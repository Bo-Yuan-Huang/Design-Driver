
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire [15:0] _26851_;
  wire [7:0] _26852_;
  wire [7:0] _26853_;
  wire [7:0] _26854_;
  wire [7:0] _26855_;
  wire [7:0] _26856_;
  wire [7:0] _26857_;
  wire [7:0] _26858_;
  wire [7:0] _26859_;
  wire [7:0] _26860_;
  wire [7:0] _26861_;
  wire [7:0] _26862_;
  wire [7:0] _26863_;
  wire [7:0] _26864_;
  wire [7:0] _26865_;
  wire [7:0] _26866_;
  wire [7:0] _26867_;
  wire _26868_;
  wire [7:0] _26869_;
  wire [2:0] _26870_;
  wire [2:0] _26871_;
  wire [1:0] _26872_;
  wire [7:0] _26873_;
  wire _26874_;
  wire [1:0] _26875_;
  wire [1:0] _26876_;
  wire [2:0] _26877_;
  wire [2:0] _26878_;
  wire [1:0] _26879_;
  wire [3:0] _26880_;
  wire [1:0] _26881_;
  wire _26882_;
  wire [7:0] _26883_;
  wire [7:0] _26884_;
  wire [7:0] _26885_;
  wire [7:0] _26886_;
  wire [7:0] _26887_;
  wire [7:0] _26888_;
  wire [7:0] _26889_;
  wire [7:0] _26890_;
  wire [15:0] _26891_;
  wire [15:0] _26892_;
  wire _26893_;
  wire [4:0] _26894_;
  wire [7:0] _26895_;
  wire [7:0] _26896_;
  wire _26897_;
  wire _26898_;
  wire [15:0] _26899_;
  wire [15:0] _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire [7:0] _26904_;
  wire [2:0] _26905_;
  wire [7:0] _26906_;
  wire _26907_;
  wire [7:0] _26908_;
  wire _26909_;
  wire _26910_;
  wire [3:0] _26911_;
  wire [31:0] _26912_;
  wire [31:0] _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire [15:0] _26917_;
  wire _26918_;
  wire _26919_;
  wire [7:0] _26920_;
  wire _26921_;
  wire [2:0] _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire [7:0] _27317_;
  wire _27318_;
  wire [3:0] _27319_;
  wire _27320_;
  wire _27321_;
  wire [7:0] _27322_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_22761_, rst);
  not (_22762_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_22763_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_22764_, _22763_, _22762_);
  not (_22765_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22767_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_22768_, _22767_, _22765_);
  and (_22769_, _22768_, _22764_);
  and (_22770_, _22769_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_22771_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_22772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_22773_, _22770_, _22772_);
  or (_22774_, _22773_, _22771_);
  and (_26891_[11], _22774_, _22761_);
  and (_22775_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_22776_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_22777_, _22770_, _22776_);
  or (_22778_, _22777_, _22775_);
  and (_26891_[12], _22778_, _22761_);
  and (_22779_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_22780_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_22781_, _22770_, _22780_);
  or (_22782_, _22781_, _22779_);
  and (_26891_[13], _22782_, _22761_);
  and (_22783_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_22784_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_22785_, _22770_, _22784_);
  or (_22787_, _22785_, _22783_);
  and (_26891_[14], _22787_, _22761_);
  and (_22788_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_22789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22790_, _22770_, _22789_);
  or (_22791_, _22790_, _22788_);
  and (_26892_[0], _22791_, _22761_);
  and (_22792_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_22794_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_22795_, _22770_, _22794_);
  or (_22796_, _22795_, _22792_);
  and (_26892_[1], _22796_, _22761_);
  and (_22797_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_22798_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_22799_, _22770_, _22798_);
  or (_22800_, _22799_, _22797_);
  and (_26892_[2], _22800_, _22761_);
  and (_22801_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_22802_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22803_, _22770_, _22802_);
  or (_22804_, _22803_, _22801_);
  and (_26892_[3], _22804_, _22761_);
  or (_22805_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not (_22807_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_22808_, _22770_, _22807_);
  and (_22809_, _22808_, _22761_);
  and (_26892_[4], _22809_, _22805_);
  and (_22810_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_22811_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_22812_, _22770_, _22811_);
  or (_22813_, _22812_, _22810_);
  and (_26892_[5], _22813_, _22761_);
  and (_22814_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_22815_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_22816_, _22770_, _22815_);
  or (_22817_, _22816_, _22814_);
  and (_26892_[6], _22817_, _22761_);
  and (_22818_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_22820_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22821_, _22770_, _22820_);
  or (_22822_, _22821_, _22818_);
  and (_26892_[7], _22822_, _22761_);
  or (_22823_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not (_22824_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_22825_, _22770_, _22824_);
  and (_22826_, _22825_, _22761_);
  and (_26892_[8], _22826_, _22823_);
  and (_22827_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not (_22828_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_22829_, _22770_, _22828_);
  or (_22830_, _22829_, _22827_);
  and (_26892_[9], _22830_, _22761_);
  and (_22832_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not (_22833_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_22834_, _22770_, _22833_);
  or (_22835_, _22834_, _22832_);
  and (_26892_[10], _22835_, _22761_);
  and (_22836_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_22837_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_22838_, _22770_, _22837_);
  or (_22839_, _22838_, _22836_);
  and (_26892_[11], _22839_, _22761_);
  or (_22840_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nand (_22841_, _22770_, _22776_);
  and (_22842_, _22841_, _22761_);
  and (_26892_[12], _22842_, _22840_);
  and (_22843_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_22844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_22846_, _22770_, _22844_);
  or (_22847_, _22846_, _22843_);
  and (_26892_[13], _22847_, _22761_);
  or (_22848_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand (_22849_, _22770_, _22784_);
  and (_22850_, _22849_, _22761_);
  and (_26892_[14], _22850_, _22848_);
  and (_22852_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_22853_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_22854_, _22770_, _22853_);
  or (_22855_, _22854_, _22852_);
  and (_26891_[10], _22855_, _22761_);
  not (_22856_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not (_22857_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22858_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _22765_);
  and (_22860_, _22858_, _22857_);
  and (_22861_, _22860_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_22862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_22863_, _22862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_22864_, _22863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_22865_, _22864_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_22866_, _22865_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_22867_, _22866_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_22868_, _22867_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_22869_, _22867_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_22870_, _22869_, _22868_);
  and (_22871_, _22870_, _22861_);
  not (_22872_, _22871_);
  and (_22873_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22874_, _22873_, _22858_);
  nor (_22875_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_22876_, _22875_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_22877_, _22876_, _22857_);
  and (_22878_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_22880_, _22878_, _22874_);
  nor (_22881_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22883_, _22881_, _22858_);
  and (_22884_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_22885_, _22876_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22886_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_22887_, _22886_, _22884_);
  and (_22889_, _22887_, _22880_);
  nand (_22890_, _22889_, _22872_);
  nor (_22891_, _22890_, _22856_);
  not (_22892_, _22864_);
  not (_22893_, _22861_);
  nor (_22895_, _22863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_22896_, _22895_, _22893_);
  and (_22897_, _22896_, _22892_);
  not (_22899_, _22897_);
  nor (_22900_, _22881_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_22902_, _22900_, _22858_);
  not (_22903_, _22902_);
  and (_22905_, _22903_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_22906_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_22908_, _22906_, _22905_);
  and (_22909_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_22910_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_22911_, _22910_, _22909_);
  and (_22912_, _22911_, _22908_);
  and (_22913_, _22912_, _22899_);
  not (_22914_, _22913_);
  and (_22915_, _22914_, _22891_);
  and (_22916_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_22917_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_22918_, _22917_, _22916_);
  and (_22919_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_22920_, _22919_);
  not (_22921_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_22922_, _22861_, _22921_);
  and (_22923_, _22903_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_22924_, _22923_, _22922_);
  and (_22925_, _22924_, _22920_);
  and (_22926_, _22925_, _22918_);
  nor (_22927_, _22926_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22928_, _22927_, _22915_);
  and (_22929_, \oc8051_top_1.oc8051_decoder1.wr , _22765_);
  not (_22930_, _22929_);
  not (_22931_, _22890_);
  nor (_22932_, _22931_, _22860_);
  nor (_22933_, _22932_, _22930_);
  not (_22934_, _22933_);
  nor (_22936_, _22934_, _22928_);
  nor (_22937_, _22864_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_22938_, _22937_);
  nor (_22939_, _22893_, _22865_);
  and (_22940_, _22939_, _22938_);
  not (_22941_, _22940_);
  and (_22942_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_22943_, _22942_, _22874_);
  and (_22944_, _22903_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_22945_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_22946_, _22945_, _22944_);
  and (_22947_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_22948_, _22947_);
  and (_22949_, _22948_, _22946_);
  and (_22950_, _22949_, _22943_);
  and (_22951_, _22950_, _22941_);
  not (_22952_, _22951_);
  and (_22953_, _22952_, _22891_);
  nor (_22954_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_22955_, _22954_, _22862_);
  and (_22956_, _22955_, _22861_);
  and (_22957_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_22958_, _22957_, _22956_);
  and (_22959_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_22960_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_22962_, _22903_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_22963_, _22962_, _22960_);
  nor (_22964_, _22963_, _22959_);
  and (_22965_, _22964_, _22958_);
  nor (_22966_, _22965_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22967_, _22966_, _22953_);
  nor (_22968_, _22967_, _22934_);
  and (_22969_, _22968_, _22936_);
  nor (_22970_, _22866_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_22971_, _22970_);
  nor (_22972_, _22893_, _22867_);
  and (_22973_, _22972_, _22971_);
  not (_22974_, _22973_);
  and (_22975_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_22976_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_22977_, _22976_, _22975_);
  and (_22978_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  nor (_22979_, _22978_, _22874_);
  and (_22980_, _22979_, _22977_);
  and (_22981_, _22980_, _22974_);
  not (_22982_, _22981_);
  and (_22983_, _22982_, _22891_);
  nor (_22984_, _22913_, _22891_);
  nor (_22985_, _22984_, _22983_);
  nor (_22986_, _22985_, _22934_);
  nor (_22987_, _22865_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_22988_, _22987_);
  nor (_22989_, _22893_, _22866_);
  and (_22990_, _22989_, _22988_);
  not (_22991_, _22990_);
  and (_22992_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_22993_, _22992_, _22874_);
  and (_22994_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_22995_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor (_22996_, _22995_, _22994_);
  and (_22997_, _22996_, _22993_);
  and (_22998_, _22997_, _22991_);
  not (_22999_, _22998_);
  and (_23000_, _22999_, _22891_);
  nor (_23001_, _22862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_23002_, _23001_, _22863_);
  and (_23003_, _23002_, _22861_);
  and (_23004_, _22877_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_23005_, _23004_, _23003_);
  and (_23006_, _22903_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  not (_23007_, _23006_);
  and (_23008_, _22885_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_23009_, _22883_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_23010_, _23009_, _23008_);
  and (_23011_, _23010_, _23007_);
  and (_23012_, _23011_, _23005_);
  nor (_23013_, _23012_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23014_, _23013_, _23000_);
  nor (_23015_, _23014_, _22934_);
  and (_23016_, _23015_, _22986_);
  and (_23017_, _23016_, _22969_);
  nor (_23018_, _22951_, _22891_);
  and (_23019_, _23018_, _22933_);
  nor (_23020_, _22999_, _22891_);
  not (_23021_, _23020_);
  and (_23022_, _23021_, _22933_);
  nor (_23023_, _23022_, _23019_);
  nor (_23024_, _22981_, _22891_);
  and (_23025_, _23024_, _22933_);
  and (_23027_, _23025_, _22931_);
  and (_23028_, _23027_, _23023_);
  and (_23029_, _23028_, _23017_);
  not (_23030_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_23031_, _22765_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23032_, _23031_, _23030_);
  and (_23033_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _22765_);
  and (_23034_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _22765_);
  nor (_23035_, _23034_, _23033_);
  and (_23037_, _23035_, _23032_);
  not (_23038_, _23037_);
  not (_23039_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_23040_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_23041_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_23042_, _23041_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_23043_, _23042_, _23040_);
  or (_23044_, _23043_, _23039_);
  nor (_23045_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_23046_, _23045_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_23047_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_23049_, _23047_, _23044_);
  not (_23050_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or (_23051_, _23042_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23052_, _23051_, _23050_);
  nor (_23054_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_23055_, _23054_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_23056_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_23057_, _23056_, _23052_);
  and (_23058_, _23057_, _23049_);
  nand (_23059_, _23054_, _23041_);
  or (_23060_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_23061_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23062_, _23061_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_23063_, _23062_, _23060_);
  not (_23064_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_23065_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23064_);
  or (_23066_, _23065_, _23063_);
  nand (_23067_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23064_);
  or (_23068_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_23069_, _23068_, _23066_);
  or (_23070_, _23069_, _23059_);
  and (_23071_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_23072_, _23071_, _23040_);
  nand (_23073_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_23074_, _23071_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_23075_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_23076_, _23075_, _23073_);
  and (_23077_, _23076_, _23070_);
  and (_23078_, _23077_, _23058_);
  or (_23080_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_23081_, _23080_, _23069_);
  and (_23082_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_23083_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_23084_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_23086_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_23087_, _23086_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor (_23088_, _23087_, _23084_);
  nor (_23089_, _23088_, _23083_);
  and (_23090_, _23089_, _23081_);
  nor (_23091_, _23090_, _23078_);
  not (_23092_, _23091_);
  not (_23093_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_23095_, _23043_, _23093_);
  nand (_23096_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_23098_, _23096_, _23095_);
  not (_23099_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_23100_, _23051_, _23099_);
  nand (_23101_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_23102_, _23101_, _23100_);
  and (_23103_, _23102_, _23098_);
  or (_23104_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_23105_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23061_);
  and (_23106_, _23105_, _23104_);
  or (_23107_, _23106_, _23065_);
  or (_23108_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_23109_, _23108_, _23107_);
  or (_23110_, _23109_, _23059_);
  nand (_23111_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nand (_23112_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_23113_, _23112_, _23111_);
  and (_23114_, _23113_, _23110_);
  nand (_23115_, _23114_, _23103_);
  or (_23116_, _23109_, _23080_);
  nand (_23117_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not (_23118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_23119_, _23087_, _23118_);
  and (_23120_, _23119_, _23117_);
  nand (_23121_, _23120_, _23116_);
  and (_23122_, _23121_, _23115_);
  nor (_23123_, _23121_, _23115_);
  nor (_23124_, _23123_, _23122_);
  not (_23125_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_23126_, _23043_, _23125_);
  nand (_23127_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_23128_, _23127_, _23126_);
  nand (_23129_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  not (_23130_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_23131_, _23051_, _23130_);
  and (_23132_, _23131_, _23129_);
  and (_23133_, _23132_, _23128_);
  or (_23134_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_23135_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23061_);
  and (_23136_, _23135_, _23134_);
  or (_23137_, _23136_, _23065_);
  or (_23138_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_23139_, _23138_, _23137_);
  or (_23140_, _23139_, _23059_);
  nand (_23141_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_23142_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_23143_, _23142_, _23141_);
  and (_23145_, _23143_, _23140_);
  and (_23146_, _23145_, _23133_);
  or (_23147_, _23139_, _23080_);
  nand (_23148_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_23149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_23150_, _23087_, _23149_);
  and (_23151_, _23150_, _23148_);
  and (_23152_, _23151_, _23147_);
  nor (_23153_, _23152_, _23146_);
  and (_23154_, _23152_, _23146_);
  nor (_23155_, _23154_, _23153_);
  not (_23156_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_23158_, _23043_, _23156_);
  nand (_23159_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_23160_, _23159_, _23158_);
  not (_23161_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_23162_, _23051_, _23161_);
  nand (_23163_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_23164_, _23163_, _23162_);
  and (_23165_, _23164_, _23160_);
  or (_23166_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_23167_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23061_);
  and (_23168_, _23167_, _23166_);
  or (_23169_, _23168_, _23065_);
  or (_23170_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_23171_, _23170_, _23169_);
  or (_23172_, _23171_, _23059_);
  nand (_23174_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nand (_23175_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_23176_, _23175_, _23174_);
  and (_23177_, _23176_, _23172_);
  and (_23178_, _23177_, _23165_);
  or (_23179_, _23171_, _23080_);
  nand (_23180_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not (_23181_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_23182_, _23087_, _23181_);
  and (_23183_, _23182_, _23180_);
  and (_23184_, _23183_, _23179_);
  nor (_23185_, _23184_, _23178_);
  and (_23187_, _23184_, _23178_);
  nor (_23188_, _23187_, _23185_);
  nand (_23189_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand (_23190_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_23191_, _23190_, _23189_);
  not (_23192_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_23193_, _23043_, _23192_);
  nand (_23194_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_23195_, _23194_, _23193_);
  and (_23196_, _23195_, _23191_);
  or (_23197_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_23198_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23061_);
  and (_23199_, _23198_, _23197_);
  or (_23200_, _23199_, _23065_);
  or (_23202_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_23203_, _23202_, _23200_);
  or (_23205_, _23203_, _23059_);
  not (_23206_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_23207_, _23051_, _23206_);
  nand (_23208_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_23209_, _23208_, _23207_);
  and (_23210_, _23209_, _23205_);
  nand (_23211_, _23210_, _23196_);
  or (_23212_, _23203_, _23080_);
  nand (_23213_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_23214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_23215_, _23087_, _23214_);
  and (_23216_, _23215_, _23213_);
  nand (_23217_, _23216_, _23212_);
  and (_23218_, _23217_, _23211_);
  nor (_23219_, _23217_, _23211_);
  nor (_23220_, _23219_, _23218_);
  not (_23221_, _23220_);
  not (_23222_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_23223_, _23043_, _23222_);
  nand (_23224_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_23225_, _23224_, _23223_);
  nand (_23226_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  not (_23227_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_23228_, _23051_, _23227_);
  and (_23229_, _23228_, _23226_);
  and (_23230_, _23229_, _23225_);
  or (_23231_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_23232_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23061_);
  and (_23233_, _23232_, _23231_);
  or (_23234_, _23233_, _23065_);
  or (_23235_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_23236_, _23235_, _23234_);
  or (_23237_, _23236_, _23059_);
  nand (_23238_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand (_23239_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_23240_, _23239_, _23238_);
  and (_23241_, _23240_, _23237_);
  nand (_23242_, _23241_, _23230_);
  or (_23243_, _23236_, _23080_);
  nand (_23244_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not (_23245_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_23246_, _23087_, _23245_);
  and (_23247_, _23246_, _23244_);
  nand (_23248_, _23247_, _23243_);
  and (_23249_, _23248_, _23242_);
  and (_23251_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_23252_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_23253_, _23043_, _23252_);
  nor (_23254_, _23253_, _23251_);
  and (_23255_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_23256_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_23257_, _23256_, _23255_);
  and (_23258_, _23257_, _23254_);
  or (_23259_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_23260_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23061_);
  and (_23261_, _23260_, _23259_);
  or (_23262_, _23261_, _23065_);
  or (_23263_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_23264_, _23263_, _23262_);
  or (_23265_, _23264_, _23059_);
  not (_23266_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_23267_, _23051_, _23266_);
  and (_23268_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_23269_, _23268_, _23267_);
  and (_23270_, _23269_, _23265_);
  and (_23271_, _23270_, _23258_);
  or (_23273_, _23264_, _23080_);
  nand (_23274_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not (_23275_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_23276_, _23087_, _23275_);
  and (_23277_, _23276_, _23274_);
  and (_23278_, _23277_, _23273_);
  nor (_23279_, _23278_, _23271_);
  nor (_23280_, _23248_, _23242_);
  nor (_23281_, _23280_, _23249_);
  and (_23282_, _23281_, _23279_);
  nor (_23283_, _23282_, _23249_);
  nor (_23284_, _23283_, _23221_);
  nor (_23285_, _23284_, _23218_);
  nor (_23286_, _23285_, _23188_);
  and (_23287_, _23285_, _23188_);
  nor (_23288_, _23287_, _23286_);
  not (_23289_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_23290_, _23289_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  or (_23291_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_23292_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23061_);
  and (_23293_, _23292_, _23291_);
  nand (_23295_, _23293_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_23296_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23297_, _23199_, _23296_);
  nand (_23298_, _23297_, _23295_);
  nand (_23299_, _23298_, _23290_);
  not (_23300_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23301_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _23300_);
  nand (_23302_, _23233_, _23296_);
  nand (_23303_, _23106_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23304_, _23303_, _23302_);
  nand (_23305_, _23304_, _23301_);
  and (_23306_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23307_, _23306_, _23296_);
  nand (_23308_, _23307_, _23168_);
  and (_23309_, _23306_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23310_, _23309_, _23063_);
  and (_23311_, _23310_, _23308_);
  nor (_23312_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23313_, _23312_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23314_, _23313_, _23136_);
  and (_23315_, _23312_, _23296_);
  nand (_23316_, _23315_, _23261_);
  and (_23317_, _23316_, _23314_);
  and (_23318_, _23317_, _23311_);
  and (_23319_, _23318_, _23305_);
  nand (_23320_, _23319_, _23299_);
  nand (_23321_, _23320_, _23067_);
  and (_23322_, _23065_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_23323_, _23322_);
  nand (_23324_, _23323_, _23321_);
  and (_23325_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_23326_, _23325_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_23327_, _23326_);
  and (_23328_, _23327_, _23324_);
  and (_23329_, _23327_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_23330_, _23329_, _23328_);
  and (_23332_, _23278_, _23271_);
  nor (_23333_, _23332_, _23279_);
  and (_23334_, _23333_, _23330_);
  and (_23335_, _23334_, _23281_);
  and (_23337_, _23283_, _23221_);
  nor (_23338_, _23337_, _23284_);
  and (_23339_, _23338_, _23335_);
  not (_23340_, _23339_);
  nor (_23341_, _23340_, _23288_);
  nor (_23342_, _23285_, _23187_);
  or (_23344_, _23342_, _23185_);
  or (_23345_, _23344_, _23341_);
  and (_23346_, _23345_, _23155_);
  and (_23347_, _23346_, _23124_);
  not (_23348_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_23349_, _23043_, _23348_);
  nand (_23350_, _23046_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_23351_, _23350_, _23349_);
  not (_23352_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_23353_, _23051_, _23352_);
  nand (_23354_, _23055_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_23355_, _23354_, _23353_);
  and (_23356_, _23355_, _23351_);
  or (_23358_, _23293_, _23065_);
  or (_23359_, _23067_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_23360_, _23359_, _23358_);
  or (_23361_, _23360_, _23059_);
  nand (_23362_, _23072_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_23363_, _23074_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_23364_, _23363_, _23362_);
  and (_23365_, _23364_, _23361_);
  and (_23366_, _23365_, _23356_);
  or (_23367_, _23360_, _23080_);
  nand (_23368_, _23082_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_23369_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_23370_, _23087_, _23369_);
  and (_23371_, _23370_, _23368_);
  nand (_23372_, _23371_, _23367_);
  not (_23373_, _23372_);
  nor (_23374_, _23373_, _23366_);
  and (_23375_, _23373_, _23366_);
  nor (_23376_, _23375_, _23374_);
  not (_23377_, _23376_);
  and (_23378_, _23153_, _23124_);
  nor (_23379_, _23378_, _23122_);
  nor (_23380_, _23379_, _23377_);
  and (_23381_, _23379_, _23377_);
  nor (_23382_, _23381_, _23380_);
  and (_23383_, _23382_, _23347_);
  not (_23384_, _23383_);
  nor (_23385_, _23380_, _23374_);
  and (_23386_, _23385_, _23384_);
  and (_23387_, _23090_, _23078_);
  nor (_23388_, _23387_, _23091_);
  not (_23389_, _23388_);
  or (_23390_, _23389_, _23386_);
  and (_23391_, _23390_, _23092_);
  nor (_23392_, _23391_, _23038_);
  not (_23393_, _23392_);
  not (_23394_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23395_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22765_);
  and (_23397_, _23395_, _23394_);
  and (_23398_, _23397_, _23035_);
  not (_23399_, _23398_);
  not (_23401_, _23090_);
  and (_23402_, _23401_, _23078_);
  nor (_23403_, _23372_, _23366_);
  and (_23404_, _23120_, _23116_);
  and (_23405_, _23404_, _23115_);
  nand (_23406_, _23151_, _23147_);
  and (_23407_, _23406_, _23146_);
  nor (_23408_, _23407_, _23124_);
  nor (_23409_, _23408_, _23405_);
  nor (_23410_, _23409_, _23376_);
  nor (_23411_, _23410_, _23403_);
  and (_23412_, _23409_, _23376_);
  nor (_23413_, _23412_, _23410_);
  not (_23414_, _23413_);
  and (_23415_, _23407_, _23124_);
  nor (_23416_, _23415_, _23408_);
  not (_23417_, _23416_);
  not (_23418_, _23155_);
  nand (_23419_, _23277_, _23273_);
  and (_23420_, _23419_, _23271_);
  nor (_23422_, _23420_, _23281_);
  and (_23423_, _23247_, _23243_);
  and (_23424_, _23423_, _23242_);
  nor (_23425_, _23424_, _23422_);
  nor (_23426_, _23425_, _23220_);
  and (_23427_, _23216_, _23212_);
  and (_23428_, _23427_, _23211_);
  nor (_23429_, _23428_, _23426_);
  nor (_23430_, _23429_, _23188_);
  and (_23431_, _23429_, _23188_);
  nor (_23432_, _23431_, _23430_);
  and (_23433_, _23425_, _23220_);
  nor (_23434_, _23433_, _23426_);
  not (_23435_, _23434_);
  and (_23436_, _23420_, _23281_);
  nor (_23437_, _23436_, _23422_);
  not (_23438_, _23437_);
  not (_23439_, _23333_);
  and (_23440_, _23439_, _23330_);
  and (_23441_, _23440_, _23438_);
  and (_23442_, _23441_, _23435_);
  not (_23443_, _23442_);
  nor (_23444_, _23443_, _23432_);
  nand (_23445_, _23183_, _23179_);
  or (_23446_, _23445_, _23178_);
  and (_23447_, _23445_, _23178_);
  or (_23448_, _23429_, _23447_);
  and (_23449_, _23448_, _23446_);
  or (_23451_, _23449_, _23444_);
  and (_23452_, _23451_, _23418_);
  and (_23453_, _23452_, _23417_);
  and (_23454_, _23453_, _23414_);
  nor (_23455_, _23454_, _23411_);
  nor (_23456_, _23455_, _23388_);
  nor (_23457_, _23456_, _23402_);
  nor (_23458_, _23457_, _23399_);
  not (_23459_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_23460_, _23033_, _23459_);
  and (_23461_, _23460_, _23032_);
  not (_23462_, _23461_);
  nor (_23463_, _23242_, _23211_);
  nor (_23464_, _23463_, _23178_);
  and (_23465_, _23323_, _23321_);
  or (_23466_, _23326_, _23465_);
  not (_23467_, _23329_);
  and (_23468_, _23467_, _23466_);
  not (_23469_, _23115_);
  and (_23470_, _23366_, _23469_);
  nor (_23471_, _23470_, _23078_);
  and (_23472_, _23471_, _23468_);
  nor (_23473_, _23472_, _23464_);
  nor (_23474_, _23473_, _23462_);
  not (_23475_, _23474_);
  and (_23476_, _23467_, _23465_);
  not (_23477_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23478_, _23034_, _23477_);
  and (_23479_, _23478_, _23032_);
  nor (_23480_, _23395_, _23031_);
  and (_23481_, _23480_, _23478_);
  and (_23482_, _23481_, _23466_);
  nor (_23483_, _23482_, _23479_);
  nor (_23484_, _23483_, _23476_);
  not (_23485_, _23484_);
  and (_23486_, _23326_, _23324_);
  and (_23487_, _23478_, _23397_);
  and (_23488_, _23395_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23489_, _23488_, _23460_);
  and (_23490_, _23489_, _23324_);
  nor (_23491_, _23490_, _23487_);
  nor (_23492_, _23491_, _23486_);
  not (_23493_, _23492_);
  and (_23494_, _23480_, _23035_);
  nor (_23495_, _23471_, _23462_);
  nor (_23496_, _23495_, _23494_);
  nor (_23497_, _23496_, _23468_);
  and (_23498_, _23460_, _23397_);
  and (_23499_, _23498_, _23467_);
  and (_23500_, _23034_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23501_, _23500_, _23480_);
  and (_23502_, _23501_, _23329_);
  nor (_23503_, _23502_, _23499_);
  nor (_23504_, _23503_, _23328_);
  not (_23505_, _23271_);
  and (_23506_, _23500_, _23032_);
  and (_23507_, _23506_, _23505_);
  not (_23508_, _23078_);
  and (_23509_, _23488_, _23478_);
  and (_23510_, _23509_, _23508_);
  nor (_23511_, _23510_, _23507_);
  not (_23512_, _23511_);
  nor (_23513_, _23512_, _23504_);
  not (_23514_, _23513_);
  nor (_23515_, _23514_, _23497_);
  and (_23517_, _23515_, _23493_);
  and (_23518_, _23517_, _23485_);
  and (_23519_, _23518_, _23475_);
  not (_23520_, _23519_);
  nor (_23521_, _23520_, _23458_);
  and (_23522_, _23521_, _23393_);
  and (_23523_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23524_, _23523_, _23306_);
  nor (_23525_, _23524_, _23522_);
  nor (_23526_, _23309_, _22856_);
  and (_23527_, _23526_, _23063_);
  and (_23528_, _23480_, _23460_);
  not (_23529_, _23528_);
  and (_23530_, _23032_, _23459_);
  and (_23531_, _23488_, _23035_);
  nor (_23532_, _23531_, _23530_);
  and (_23533_, _23532_, _23529_);
  and (_23534_, _23500_, _23030_);
  not (_23535_, _23534_);
  and (_23536_, _23478_, _23395_);
  nor (_23537_, _23536_, _23494_);
  and (_23538_, _23537_, _23535_);
  and (_23540_, _23538_, _23533_);
  nor (_23541_, _23540_, _23078_);
  not (_23542_, _23541_);
  and (_23543_, _23500_, _23397_);
  not (_23544_, _23543_);
  and (_23545_, _23463_, _23271_);
  and (_23546_, _23545_, _23178_);
  and (_23547_, _23546_, _23146_);
  and (_23548_, _23547_, _23470_);
  nor (_23549_, _23548_, _23468_);
  not (_23550_, _23366_);
  not (_23551_, _23146_);
  not (_23552_, _23178_);
  and (_23553_, _23505_, _23242_);
  and (_23554_, _23553_, _23211_);
  and (_23555_, _23554_, _23552_);
  and (_23556_, _23555_, _23551_);
  and (_23557_, _23556_, _23115_);
  and (_23558_, _23557_, _23550_);
  nor (_23560_, _23558_, _23330_);
  or (_23561_, _23560_, _23549_);
  nor (_23562_, _23561_, _23508_);
  and (_23563_, _23561_, _23508_);
  nor (_23564_, _23563_, _23562_);
  nor (_23565_, _23564_, _23544_);
  and (_23566_, _23330_, _23090_);
  not (_23567_, _23566_);
  and (_23568_, _23500_, _23488_);
  not (_23569_, _23568_);
  and (_23570_, _23468_, _23078_);
  nor (_23571_, _23570_, _23569_);
  and (_23572_, _23571_, _23567_);
  and (_23573_, _23481_, _23388_);
  and (_23574_, _23489_, _23091_);
  not (_23575_, _23479_);
  nor (_23576_, _23575_, _23387_);
  and (_23577_, _23498_, _23078_);
  or (_23578_, _23577_, _23576_);
  or (_23579_, _23578_, _23574_);
  nor (_23580_, _23579_, _23573_);
  not (_23581_, _23580_);
  nor (_23582_, _23581_, _23572_);
  not (_23583_, _23582_);
  nor (_23584_, _23583_, _23565_);
  and (_23585_, _23584_, _23542_);
  nor (_23586_, _23585_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or (_23587_, _23586_, _23527_);
  or (_23588_, _23587_, _23525_);
  and (_23589_, _23588_, _22933_);
  and (_23590_, _23589_, _23029_);
  not (_23591_, _23029_);
  and (_23592_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or (_24563_, _23592_, _23590_);
  nor (_23593_, _23015_, _22986_);
  and (_23594_, _23593_, _22969_);
  and (_23595_, _23019_, _22999_);
  nor (_23596_, _22982_, _22890_);
  nor (_23597_, _23596_, _22891_);
  not (_23598_, _23597_);
  and (_23599_, _23598_, _23595_);
  and (_23601_, _23599_, _23594_);
  nand (_23602_, _23523_, _23301_);
  nor (_23603_, _23602_, _23522_);
  and (_23604_, _23468_, _23469_);
  not (_23605_, _23604_);
  and (_23606_, _23330_, _23404_);
  nor (_23607_, _23606_, _23569_);
  and (_23608_, _23607_, _23605_);
  nor (_23609_, _23556_, _23330_);
  nor (_23610_, _23547_, _23468_);
  nor (_23611_, _23610_, _23609_);
  and (_23612_, _23611_, _23115_);
  nor (_23613_, _23611_, _23115_);
  or (_23614_, _23613_, _23544_);
  nor (_23615_, _23614_, _23612_);
  nor (_23616_, _23615_, _23608_);
  and (_23617_, _23481_, _23124_);
  and (_23618_, _23489_, _23122_);
  nor (_23619_, _23575_, _23123_);
  and (_23620_, _23498_, _23469_);
  or (_23621_, _23620_, _23619_);
  or (_23622_, _23621_, _23618_);
  nor (_23623_, _23622_, _23617_);
  not (_23624_, _23540_);
  and (_23625_, _23624_, _23115_);
  not (_23626_, _23625_);
  and (_23627_, _23626_, _23623_);
  and (_23628_, _23627_, _23616_);
  nor (_23629_, _23628_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23630_, _23301_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_23631_, _23106_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23632_, _23631_, _23630_);
  or (_23633_, _23632_, _23629_);
  or (_23634_, _23633_, _23603_);
  and (_23635_, _23634_, _22933_);
  and (_23636_, _23635_, _23601_);
  not (_23637_, _23601_);
  and (_23638_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or (_27242_, _23638_, _23636_);
  and (_23639_, _22968_, _22928_);
  and (_23640_, _23015_, _22985_);
  and (_23641_, _23640_, _23639_);
  and (_23642_, _22981_, _22890_);
  and (_23643_, _23642_, _23595_);
  and (_23644_, _23643_, _23641_);
  and (_23645_, _23644_, _23589_);
  not (_23646_, _23644_);
  and (_23647_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_27084_, _23647_, _23645_);
  nor (_23648_, _22968_, _22936_);
  and (_23649_, _23648_, _23593_);
  and (_23650_, _23019_, _22998_);
  and (_23651_, _23650_, _23027_);
  and (_23652_, _23651_, _23649_);
  and (_23653_, _23296_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23654_, _23653_, _23312_);
  not (_23655_, _23654_);
  nor (_23656_, _23655_, _23522_);
  and (_23657_, _23568_, _23419_);
  and (_23658_, _23543_, _23271_);
  nor (_23659_, _23658_, _23657_);
  and (_23660_, _23489_, _23279_);
  and (_23661_, _23498_, _23271_);
  nor (_23662_, _23661_, _23660_);
  and (_23663_, _23662_, _23659_);
  nor (_23664_, _23540_, _23271_);
  and (_23665_, _23481_, _23333_);
  nor (_23666_, _23575_, _23332_);
  or (_23667_, _23666_, _23665_);
  nor (_23668_, _23667_, _23664_);
  and (_23669_, _23668_, _23663_);
  nand (_23670_, _23669_, _22856_);
  or (_23671_, _23261_, _22856_);
  and (_23672_, _23671_, _23655_);
  and (_23673_, _23672_, _23670_);
  or (_23674_, _23673_, _23656_);
  and (_23676_, _23674_, _22933_);
  and (_23677_, _23676_, _23652_);
  not (_23678_, _23652_);
  and (_23680_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or (_11638_, _23680_, _23677_);
  nand (_23681_, _23653_, _23290_);
  nor (_23682_, _23681_, _23522_);
  and (_23683_, _23568_, _23217_);
  not (_23684_, _23211_);
  or (_23685_, _23271_, _23242_);
  or (_23687_, _23468_, _23242_);
  or (_23688_, _23330_, _23271_);
  nand (_23690_, _23688_, _23687_);
  nand (_23691_, _23690_, _23685_);
  nand (_23692_, _23691_, _23684_);
  or (_23693_, _23691_, _23684_);
  and (_23694_, _23693_, _23543_);
  and (_23695_, _23694_, _23692_);
  nor (_23696_, _23695_, _23683_);
  and (_23697_, _23624_, _23211_);
  not (_23698_, _23697_);
  and (_23699_, _23481_, _23220_);
  nor (_23700_, _23575_, _23219_);
  not (_23701_, _23700_);
  and (_23702_, _23489_, _23218_);
  and (_23703_, _23498_, _23684_);
  nor (_23704_, _23703_, _23702_);
  nand (_23705_, _23704_, _23701_);
  nor (_23706_, _23705_, _23699_);
  and (_23707_, _23706_, _23698_);
  nand (_23709_, _23707_, _23696_);
  and (_23710_, _23709_, _22856_);
  and (_23711_, _23653_, _23300_);
  and (_23712_, _23653_, _23306_);
  or (_23713_, _23712_, _23523_);
  or (_23714_, _23713_, _23711_);
  and (_23715_, _23714_, _23199_);
  or (_23716_, _23715_, _23710_);
  or (_23717_, _23716_, _23682_);
  and (_23718_, _23717_, _22933_);
  and (_23719_, _23718_, _23652_);
  and (_23720_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or (_14343_, _23720_, _23719_);
  nand (_23721_, _23523_, _23290_);
  nor (_23722_, _23721_, _23522_);
  and (_23723_, _23372_, _23330_);
  and (_23724_, _23550_, _23468_);
  nor (_23725_, _23724_, _23723_);
  nor (_23726_, _23725_, _23569_);
  nor (_23728_, _23557_, _23550_);
  not (_23729_, _23728_);
  and (_23730_, _23729_, _23560_);
  and (_23731_, _23547_, _23469_);
  nor (_23732_, _23731_, _23366_);
  nor (_23733_, _23732_, _23548_);
  nor (_23734_, _23733_, _23468_);
  nor (_23735_, _23734_, _23730_);
  nor (_23736_, _23735_, _23544_);
  nor (_23737_, _23736_, _23726_);
  and (_23738_, _23481_, _23376_);
  and (_23739_, _23489_, _23374_);
  nor (_23740_, _23575_, _23375_);
  and (_23741_, _23498_, _23366_);
  or (_23742_, _23741_, _23740_);
  or (_23743_, _23742_, _23739_);
  nor (_23744_, _23743_, _23738_);
  nor (_23745_, _23540_, _23366_);
  not (_23746_, _23745_);
  and (_23747_, _23746_, _23744_);
  and (_23748_, _23747_, _23737_);
  nor (_23749_, _23748_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23750_, _23290_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_23751_, _23293_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23752_, _23751_, _23750_);
  or (_23753_, _23752_, _23749_);
  or (_23754_, _23753_, _23722_);
  and (_23755_, _23754_, _22933_);
  and (_23756_, _23755_, _23644_);
  and (_23757_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_18789_, _23757_, _23756_);
  nand (_23758_, _23653_, _23301_);
  nor (_23759_, _23758_, _23522_);
  and (_23760_, _23624_, _23242_);
  not (_23762_, _23760_);
  nand (_23763_, _23271_, _23242_);
  and (_23765_, _23763_, _23685_);
  or (_23766_, _23765_, _23468_);
  nand (_23767_, _23765_, _23468_);
  and (_23768_, _23767_, _23543_);
  nand (_23769_, _23768_, _23766_);
  and (_23770_, _23481_, _23281_);
  not (_23771_, _23770_);
  and (_23772_, _23489_, _23249_);
  not (_23773_, _23772_);
  nor (_23774_, _23575_, _23280_);
  not (_23775_, _23774_);
  and (_23776_, _23568_, _23248_);
  not (_23777_, _23242_);
  and (_23778_, _23498_, _23777_);
  nor (_23779_, _23778_, _23776_);
  and (_23780_, _23779_, _23775_);
  and (_23781_, _23780_, _23773_);
  and (_23782_, _23781_, _23771_);
  and (_23783_, _23782_, _23769_);
  and (_23784_, _23783_, _23762_);
  nor (_23785_, _23784_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23786_, _23653_, _23289_);
  or (_23787_, _23786_, _23713_);
  and (_23788_, _23787_, _23233_);
  or (_23789_, _23788_, _23785_);
  or (_23790_, _23789_, _23759_);
  and (_23791_, _23790_, _22933_);
  and (_23792_, _23791_, _23652_);
  and (_23793_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or (_20210_, _23793_, _23792_);
  and (_23794_, _23676_, _23644_);
  and (_23795_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_22709_, _23795_, _23794_);
  and (_23796_, _23014_, _22986_);
  and (_23797_, _23796_, _23639_);
  and (_23798_, _23797_, _23599_);
  and (_23799_, _23798_, _23676_);
  not (_23800_, _23798_);
  and (_23801_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or (_22729_, _23801_, _23799_);
  and (_23802_, _22967_, _22936_);
  and (_23803_, _23802_, _23016_);
  not (_23804_, _23018_);
  and (_23805_, _23022_, _23804_);
  and (_23806_, _23805_, _23027_);
  and (_23807_, _23806_, _23803_);
  and (_23808_, _23807_, _23791_);
  not (_23809_, _23807_);
  and (_23810_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_22744_, _23810_, _23808_);
  and (_23811_, _23651_, _23594_);
  not (_23812_, _23522_);
  and (_23813_, _23712_, _23812_);
  nand (_23814_, _23554_, _23468_);
  nand (_23815_, _23545_, _23330_);
  and (_23816_, _23815_, _23814_);
  nand (_23817_, _23816_, _23178_);
  or (_23818_, _23816_, _23178_);
  and (_23819_, _23818_, _23543_);
  and (_23820_, _23819_, _23817_);
  and (_23821_, _23568_, _23445_);
  nor (_23822_, _23821_, _23820_);
  and (_23823_, _23489_, _23185_);
  and (_23824_, _23498_, _23178_);
  nor (_23825_, _23824_, _23823_);
  nor (_23826_, _23540_, _23178_);
  and (_23827_, _23481_, _23188_);
  nor (_23828_, _23575_, _23187_);
  or (_23829_, _23828_, _23827_);
  nor (_23830_, _23829_, _23826_);
  and (_23831_, _23830_, _23825_);
  and (_23832_, _23831_, _23822_);
  nor (_23833_, _23832_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23834_, _23307_, _22856_);
  and (_23835_, _23834_, _23168_);
  or (_23836_, _23835_, _23833_);
  or (_23837_, _23836_, _23813_);
  and (_23838_, _23837_, _22933_);
  and (_23839_, _23838_, _23811_);
  not (_23840_, _23811_);
  and (_23841_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or (_23727_, _23841_, _23839_);
  and (_23842_, _23648_, _23016_);
  and (_23843_, _23842_, _23806_);
  and (_23844_, _23843_, _23755_);
  not (_23845_, _23843_);
  and (_23846_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or (_26943_, _23846_, _23844_);
  and (_23847_, _23843_, _23589_);
  and (_23848_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_26944_, _23848_, _23847_);
  and (_23849_, _23639_, _23016_);
  and (_23850_, _23849_, _23651_);
  and (_23851_, _23850_, _23755_);
  not (_23852_, _23850_);
  and (_23853_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or (_27310_, _23853_, _23851_);
  and (_23854_, _23796_, _22969_);
  and (_23855_, _23854_, _23806_);
  and (_23857_, _23855_, _23791_);
  not (_23858_, _23855_);
  and (_23859_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or (_24159_, _23859_, _23857_);
  and (_23861_, _23807_, _23589_);
  and (_23862_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_24183_, _23862_, _23861_);
  and (_23863_, _23802_, _23640_);
  and (_23864_, _23863_, _23643_);
  and (_23865_, _23864_, _23589_);
  not (_23866_, _23864_);
  and (_23867_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_24231_, _23867_, _23865_);
  and (_23868_, _23838_, _23807_);
  and (_23869_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_24419_, _23869_, _23868_);
  and (_23870_, _23807_, _23635_);
  and (_23871_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_24454_, _23871_, _23870_);
  and (_23872_, _23807_, _23718_);
  and (_23873_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_24727_, _23873_, _23872_);
  and (_23874_, _22998_, _22951_);
  and (_23875_, _23874_, _23642_);
  not (_23876_, _22926_);
  and (_23877_, _22965_, _23876_);
  and (_23878_, _23877_, _23012_);
  nor (_23879_, _22930_, _22860_);
  and (_23880_, _23879_, _22856_);
  not (_23881_, _23880_);
  nor (_23882_, _23881_, _22913_);
  and (_23883_, _23882_, _23878_);
  and (_23884_, _23883_, _23875_);
  or (_23885_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_23886_, _23885_, _22761_);
  and (_23887_, _23878_, _22914_);
  and (_23888_, _23875_, _23880_);
  and (_23889_, _23888_, _23887_);
  nor (_23890_, _23540_, _23146_);
  nand (_23891_, _23555_, _23468_);
  nand (_23892_, _23546_, _23330_);
  and (_23893_, _23892_, _23891_);
  or (_23894_, _23893_, _23146_);
  nand (_23895_, _23893_, _23146_);
  and (_23896_, _23895_, _23894_);
  and (_23897_, _23896_, _23543_);
  and (_23898_, _23468_, _23146_);
  and (_23899_, _23330_, _23152_);
  or (_23900_, _23899_, _23569_);
  nor (_23901_, _23900_, _23898_);
  and (_23902_, _23481_, _23155_);
  and (_23903_, _23489_, _23153_);
  nor (_23904_, _23575_, _23154_);
  and (_23906_, _23498_, _23146_);
  or (_23907_, _23906_, _23904_);
  or (_23908_, _23907_, _23903_);
  nor (_23909_, _23908_, _23902_);
  not (_23910_, _23909_);
  or (_23911_, _23910_, _23901_);
  or (_23913_, _23911_, _23897_);
  nor (_23914_, _23913_, _23890_);
  nand (_23915_, _23914_, _23889_);
  and (_24756_, _23915_, _23886_);
  and (_23916_, _23843_, _23635_);
  and (_23917_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_24790_, _23917_, _23916_);
  not (_23918_, _23012_);
  and (_23919_, _23877_, _23918_);
  and (_23920_, _23919_, _23882_);
  and (_23921_, _23920_, _23875_);
  not (_23922_, _23921_);
  or (_23923_, _23922_, _23709_);
  nor (_23924_, _22965_, _22926_);
  and (_23925_, _23924_, _23012_);
  and (_23926_, _23925_, _23882_);
  and (_23927_, _23926_, _23875_);
  not (_23928_, _23927_);
  not (_23929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  not (_23930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_23931_, _23930_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not (_23932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_23933_, _23932_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_23934_, t1_i);
  and (_23935_, _23934_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_23936_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or (_23937_, _23936_, _23933_);
  and (_23938_, _23937_, _23931_);
  and (_23939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_23940_, _23939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_23941_, _23940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_23942_, _23941_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_23943_, _23942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_23944_, _23943_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_23945_, _23944_, _23938_);
  not (_23946_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_23947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_23948_, _23947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_23949_, _23948_, _23946_);
  nor (_23950_, _23949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_23951_, _23950_, _23945_);
  nor (_23952_, _23951_, _23929_);
  and (_23953_, _23951_, _23929_);
  or (_23954_, _23953_, _23952_);
  or (_23955_, _23921_, _23954_);
  and (_23956_, _23955_, _23928_);
  and (_23958_, _23956_, _23923_);
  and (_23959_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_23961_, _23959_, _23958_);
  and (_24831_, _23961_, _22761_);
  and (_23962_, _23639_, _23593_);
  and (_23963_, _23962_, _23651_);
  and (_23964_, _23963_, _23755_);
  not (_23966_, _23963_);
  and (_23967_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_25022_, _23967_, _23964_);
  and (_23968_, _23963_, _23635_);
  and (_23969_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_25114_, _23969_, _23968_);
  and (_23971_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_23972_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_23973_, _22770_, _23972_);
  or (_23974_, _23973_, _23971_);
  and (_26891_[7], _23974_, _22761_);
  nand (_23975_, _23523_, _23312_);
  nor (_23976_, _23975_, _23522_);
  nor (_23977_, _23914_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23978_, _23313_, _22856_);
  and (_23979_, _23978_, _23136_);
  or (_23980_, _23979_, _23977_);
  or (_23981_, _23980_, _23976_);
  and (_23982_, _23981_, _22933_);
  and (_23983_, _23982_, _23963_);
  and (_23984_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_27296_, _23984_, _23983_);
  and (_23985_, _22965_, _22926_);
  and (_23986_, _23985_, _23918_);
  and (_23987_, _23986_, _23882_);
  and (_23988_, _23987_, _23875_);
  nand (_23989_, _23988_, _23585_);
  not (_23990_, _22965_);
  and (_23991_, _23990_, _22926_);
  and (_23992_, _23991_, _23012_);
  and (_23993_, _23992_, _23882_);
  and (_23994_, _23993_, _23875_);
  not (_23995_, _23994_);
  not (_23996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_23997_, _23996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_23998_, _23996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_23999_, _23998_, _23997_);
  and (_24000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_24001_, _24000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_24002_, _24001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_24003_, _24002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_24004_, _24003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_24005_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_24006_, _24005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_24007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_24009_, t0_i);
  and (_24010_, _24009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  nor (_24011_, _24010_, _24007_);
  not (_24012_, _24011_);
  not (_24013_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_24015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_24016_, _24015_, _24013_);
  and (_24017_, _24016_, _24012_);
  and (_24018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_24019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_24020_, _24019_, _24018_);
  and (_24021_, _24020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_24023_, _24021_, _24017_);
  and (_24024_, _24023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_24025_, _24024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_24026_, _24025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand (_24027_, _24026_, _24006_);
  or (_24028_, _24027_, _23997_);
  and (_24029_, _24028_, _23999_);
  and (_24030_, _24021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_24031_, _24030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_24032_, _24031_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_24033_, _24017_, _23996_);
  and (_24034_, _24033_, _24032_);
  and (_24035_, _24034_, _24005_);
  or (_24036_, _24035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_24037_, _24036_, _24029_);
  and (_24038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_24039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_24040_, _24039_, _24005_);
  not (_24041_, _24040_);
  nor (_24042_, _24041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_24043_, _24041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_24044_, _24043_, _24042_);
  and (_24045_, _24044_, _24038_);
  and (_24046_, _24017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_24047_, _24046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_24048_, _24047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_24049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_24050_, _24049_, _24048_);
  and (_24051_, _24050_, _24005_);
  or (_24052_, _24051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_24053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_24054_, _24053_);
  and (_24055_, _24023_, _24006_);
  nor (_24056_, _24055_, _24054_);
  and (_24057_, _24056_, _24052_);
  or (_24058_, _24057_, _24045_);
  or (_24059_, _24058_, _24037_);
  or (_24061_, _23988_, _24059_);
  and (_24062_, _24061_, _23995_);
  and (_24063_, _24062_, _23989_);
  and (_24064_, _23994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_24065_, _24064_, _24063_);
  and (_25345_, _24065_, _22761_);
  and (_24067_, _23718_, _23644_);
  and (_24068_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_25535_, _24068_, _24067_);
  and (_24069_, _23811_, _23791_);
  and (_24070_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or (_25648_, _24070_, _24069_);
  and (_24071_, _23811_, _23676_);
  and (_24072_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or (_25732_, _24072_, _24071_);
  and (_24073_, _23791_, _23644_);
  and (_24074_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_25768_, _24074_, _24073_);
  and (_24075_, _23963_, _23589_);
  and (_24077_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_25817_, _24077_, _24075_);
  and (_24078_, _23802_, _23593_);
  and (_24080_, _24078_, _23651_);
  and (_24081_, _24080_, _23635_);
  not (_24083_, _24080_);
  and (_24084_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_26162_, _24084_, _24081_);
  and (_24085_, _24080_, _23589_);
  and (_24086_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_26223_, _24086_, _24085_);
  and (_24087_, _24080_, _23755_);
  and (_24088_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_26374_, _24088_, _24087_);
  and (_24089_, _23962_, _23643_);
  and (_24090_, _24089_, _23676_);
  not (_24091_, _24089_);
  and (_24092_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_26425_, _24092_, _24090_);
  and (_24093_, _24078_, _23643_);
  and (_24094_, _24093_, _23589_);
  not (_24095_, _24093_);
  and (_24096_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_27079_, _24096_, _24094_);
  and (_24097_, _23963_, _23718_);
  and (_24098_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_00107_, _24098_, _24097_);
  and (_24099_, _23963_, _23791_);
  and (_24100_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_00278_, _24100_, _24099_);
  and (_24101_, _23963_, _23676_);
  and (_24102_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_00329_, _24102_, _24101_);
  and (_24103_, _23648_, _23640_);
  and (_24104_, _24103_, _23599_);
  and (_24105_, _24104_, _23676_);
  not (_24106_, _24104_);
  and (_24107_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or (_00420_, _24107_, _24105_);
  and (_24108_, _24089_, _23838_);
  and (_24109_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_00511_, _24109_, _24108_);
  and (_24110_, _24089_, _23718_);
  and (_24111_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_00592_, _24111_, _24110_);
  and (_24112_, _24089_, _23791_);
  and (_24113_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_00681_, _24113_, _24112_);
  and (_24115_, _24080_, _23838_);
  and (_24116_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_00743_, _24116_, _24115_);
  and (_24117_, _23640_, _22969_);
  and (_24118_, _23805_, _23598_);
  and (_24119_, _24118_, _24117_);
  and (_24120_, _24119_, _23755_);
  not (_24121_, _24119_);
  and (_24122_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_01076_, _24122_, _24120_);
  and (_24123_, _23849_, _23028_);
  and (_24124_, _24123_, _23791_);
  not (_24125_, _24123_);
  and (_24126_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_01170_, _24126_, _24124_);
  and (_24127_, _24093_, _23791_);
  and (_24128_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_01193_, _24128_, _24127_);
  and (_24129_, _23798_, _23791_);
  and (_24130_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or (_01215_, _24130_, _24129_);
  and (_24131_, _24123_, _23676_);
  and (_24132_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_27286_, _24132_, _24131_);
  or (_24133_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_24134_, _24133_, _22761_);
  nand (_24135_, _23889_, _23628_);
  and (_01337_, _24135_, _24134_);
  and (_24136_, _24093_, _23718_);
  and (_24137_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_01413_, _24137_, _24136_);
  and (_24138_, _24123_, _23635_);
  and (_24139_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_01582_, _24139_, _24138_);
  and (_24140_, _24123_, _23982_);
  and (_24141_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_01818_, _24141_, _24140_);
  and (_24142_, _24123_, _23838_);
  and (_24144_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_01878_, _24144_, _24142_);
  nand (_24145_, _23927_, _23585_);
  not (_24146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_24147_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_24148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _23946_);
  nor (_24149_, _24148_, _24147_);
  nor (_24150_, _24149_, _23921_);
  not (_24152_, _24150_);
  and (_24153_, _24152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_24154_, _24149_);
  and (_24155_, _23942_, _23938_);
  and (_24156_, _24155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_24158_, _24156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_24160_, _24158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_24161_, _24158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_24162_, _24161_, _24160_);
  and (_24164_, _24162_, _24154_);
  and (_24165_, _24161_, _24148_);
  and (_24166_, _24165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_24168_, _24166_, _24164_);
  nor (_24169_, _24168_, _23921_);
  or (_24170_, _24169_, _24153_);
  or (_24171_, _24170_, _23927_);
  and (_24172_, _24171_, _22761_);
  and (_01918_, _24172_, _24145_);
  and (_24174_, _24093_, _23635_);
  and (_24176_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_02051_, _24176_, _24174_);
  nand (_24178_, _23921_, _23832_);
  and (_24179_, _23945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_24180_, _24179_, _23948_);
  or (_24181_, _24180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not (_24182_, _24147_);
  and (_24184_, _24180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_24186_, _24184_, _24182_);
  and (_24187_, _24186_, _24181_);
  and (_24189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_24190_, _24179_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_24191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not (_24192_, _24191_);
  and (_24193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_24194_, _24193_, _23945_);
  nor (_24195_, _24194_, _24192_);
  and (_24196_, _24195_, _24190_);
  or (_24197_, _24196_, _24189_);
  or (_24198_, _24197_, _24187_);
  or (_24199_, _24198_, _23921_);
  and (_24200_, _24199_, _23928_);
  and (_24201_, _24200_, _24178_);
  and (_24203_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_24204_, _24203_, _24201_);
  and (_02094_, _24204_, _22761_);
  and (_24206_, _24093_, _23982_);
  and (_24207_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_27078_, _24207_, _24206_);
  and (_24209_, _23803_, _23028_);
  and (_24210_, _24209_, _23838_);
  not (_24211_, _24209_);
  and (_24213_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_27282_, _24213_, _24210_);
  and (_24214_, _23649_, _23643_);
  and (_24215_, _24214_, _23635_);
  not (_24216_, _24214_);
  and (_24217_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or (_27075_, _24217_, _24215_);
  and (_24218_, _24209_, _23755_);
  and (_24219_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_27284_, _24219_, _24218_);
  and (_24220_, _24209_, _23635_);
  and (_24221_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_27283_, _24221_, _24220_);
  and (_24222_, _24214_, _23982_);
  and (_24223_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or (_27074_, _24223_, _24222_);
  and (_24224_, _23676_, _23029_);
  and (_24225_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_27288_, _24225_, _24224_);
  and (_24226_, _24123_, _23589_);
  and (_24227_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_27287_, _24227_, _24226_);
  and (_24228_, _24214_, _23589_);
  and (_24229_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or (_27077_, _24229_, _24228_);
  not (_24232_, _22769_);
  not (_24233_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_24234_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_24235_, _24234_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_24236_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  not (_24237_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_24238_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_24239_, _24238_, _24237_);
  and (_24240_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_24241_, _24240_, _24236_);
  nor (_24242_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_24243_, _24242_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_24244_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not (_24245_, _24244_);
  and (_24246_, _24245_, _24241_);
  not (_24247_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_24248_, _24247_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_24250_, _24248_, _24237_);
  and (_24251_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_24252_, _24251_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_24253_, _24234_, _24237_);
  and (_24254_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_24255_, _24234_, _24237_);
  and (_24256_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_24257_, _24256_, _24254_);
  and (_24258_, _24257_, _24252_);
  and (_24259_, _24258_, _24246_);
  and (_24260_, _24259_, _24233_);
  nor (_24261_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _24233_);
  nor (_24262_, _24261_, _24260_);
  nor (_24263_, _24262_, _24232_);
  not (_24264_, _24263_);
  not (_24265_, _22764_);
  nor (_24266_, _22768_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_24267_, _24266_, _24265_);
  and (_24268_, _24267_, _24264_);
  not (_24269_, _24268_);
  not (_24270_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24271_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_24272_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_24273_, _24272_, _24271_);
  nand (_24274_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_24275_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_24276_, _24275_, _24274_);
  nand (_24277_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_24278_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_24279_, _24278_, _24277_);
  and (_24280_, _24279_, _24276_);
  nand (_24281_, _24280_, _24273_);
  nand (_24282_, _24281_, _24270_);
  nand (_24283_, _24282_, _24233_);
  nor (_24285_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _24233_);
  not (_24286_, _24285_);
  and (_24288_, _24286_, _24283_);
  or (_24289_, _24288_, _24232_);
  nor (_24291_, _22768_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_24292_, _24291_, _24265_);
  and (_24294_, _24292_, _24289_);
  or (_24295_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24296_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_24297_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_24299_, _24297_, _24296_);
  nand (_24300_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_24301_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_24302_, _24301_, _24300_);
  nand (_24303_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_24304_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_24305_, _24304_, _24303_);
  and (_24306_, _24305_, _24302_);
  and (_24307_, _24306_, _24299_);
  or (_24308_, _24307_, _24295_);
  and (_24309_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24310_, _24309_);
  and (_24311_, _24310_, _24308_);
  nand (_24313_, _24311_, _22769_);
  nor (_24314_, _22768_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_24316_, _24314_, _24265_);
  and (_24317_, _24316_, _24313_);
  not (_24318_, _24317_);
  and (_24319_, _24318_, _24294_);
  and (_24321_, _24319_, _24269_);
  and (_24322_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_24324_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_24325_, _24324_, _24322_);
  nand (_24327_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand (_24328_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_24329_, _24328_, _24327_);
  nand (_24330_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_24331_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_24332_, _24331_, _24330_);
  and (_24334_, _24332_, _24329_);
  and (_24335_, _24334_, _24325_);
  or (_24336_, _24335_, _24295_);
  and (_24337_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24338_, _24337_);
  and (_24340_, _24338_, _24336_);
  nand (_24341_, _24340_, _22769_);
  nor (_24343_, _22768_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_24344_, _24343_, _24265_);
  and (_24346_, _24344_, _24341_);
  not (_24347_, _24346_);
  and (_24348_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_24349_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_24350_, _24349_, _24348_);
  nand (_24351_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nand (_24352_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_24353_, _24352_, _24351_);
  nand (_24354_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_24356_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_24357_, _24356_, _24354_);
  and (_24358_, _24357_, _24353_);
  and (_24359_, _24358_, _24350_);
  or (_24360_, _24359_, _24295_);
  and (_24361_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24362_, _24361_);
  and (_24363_, _24362_, _24360_);
  nand (_24364_, _24363_, _22769_);
  nor (_24365_, _22768_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_24366_, _24365_, _24265_);
  and (_24367_, _24366_, _24364_);
  not (_24368_, _24367_);
  nor (_24369_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_24371_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_24372_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_24373_, _24372_, _24371_);
  nand (_24374_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand (_24375_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_24376_, _24375_, _24374_);
  and (_24377_, _24376_, _24373_);
  and (_24378_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_24379_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_24380_, _24379_, _24378_);
  nand (_24381_, _24380_, _24377_);
  nand (_24382_, _24381_, _24369_);
  and (_24383_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_24384_, _24383_);
  and (_24385_, _24384_, _24382_);
  nand (_24386_, _24385_, _22769_);
  nor (_24387_, _22768_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_24388_, _24387_, _24265_);
  and (_24389_, _24388_, _24386_);
  and (_24390_, _24389_, _24368_);
  and (_24391_, _24390_, _24347_);
  and (_24392_, _24391_, _24321_);
  nor (_24393_, _24367_, _24346_);
  and (_24394_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_24395_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_24396_, _24395_, _24394_);
  and (_24397_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_24398_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_24399_, _24398_, _24397_);
  and (_24400_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_24401_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_24402_, _24401_, _24400_);
  and (_24403_, _24402_, _24399_);
  nand (_24404_, _24403_, _24396_);
  nand (_24405_, _24404_, _24270_);
  nand (_24406_, _24405_, _24233_);
  nor (_24407_, _24233_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  not (_24408_, _24407_);
  and (_24409_, _24408_, _24406_);
  or (_24410_, _24409_, _24232_);
  nor (_24411_, _22768_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_24412_, _24411_, _24265_);
  and (_24413_, _24412_, _24410_);
  not (_24414_, _24294_);
  and (_24415_, _24318_, _24268_);
  and (_24416_, _24415_, _24414_);
  nand (_24417_, _24416_, _24413_);
  not (_24418_, _24417_);
  and (_24420_, _24418_, _24393_);
  and (_24421_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_24422_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_24423_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_24424_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_24425_, _24424_, _24423_);
  and (_24426_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_24427_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_24428_, _24427_, _24426_);
  nand (_24429_, _24428_, _24425_);
  or (_24430_, _24429_, _24422_);
  nor (_24431_, _24430_, _24421_);
  and (_24432_, _24431_, _24270_);
  and (_24433_, _24432_, _24233_);
  nor (_24435_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _24233_);
  nor (_24436_, _24435_, _24433_);
  nor (_24438_, _24436_, _24232_);
  not (_24439_, _24438_);
  nor (_24440_, _22768_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_24441_, _24440_, _24265_);
  and (_24443_, _24441_, _24439_);
  not (_24445_, _24443_);
  and (_24446_, _24368_, _24346_);
  and (_24447_, _24446_, _24389_);
  and (_24448_, _24447_, _24445_);
  and (_24449_, _24448_, _24418_);
  or (_24450_, _24449_, _24420_);
  and (_24451_, _24367_, _24347_);
  and (_24452_, _24451_, _24389_);
  and (_24453_, _24452_, _24445_);
  and (_24456_, _24453_, _24321_);
  and (_24457_, _24391_, _24317_);
  and (_24458_, _24443_, _24317_);
  not (_24459_, _24389_);
  and (_24460_, _24451_, _24459_);
  and (_24461_, _24460_, _24458_);
  or (_24463_, _24461_, _24457_);
  or (_24464_, _24463_, _24456_);
  or (_24465_, _24464_, _24450_);
  and (_24466_, _24319_, _24268_);
  and (_24468_, _24466_, _24445_);
  and (_24469_, _24468_, _24460_);
  and (_24470_, _24446_, _24459_);
  and (_24471_, _24470_, _24443_);
  and (_24472_, _24471_, _24466_);
  or (_24473_, _24472_, _24469_);
  nor (_24474_, _24443_, _24318_);
  and (_24475_, _24389_, _24367_);
  or (_24476_, _24475_, _24451_);
  and (_24478_, _24476_, _24474_);
  and (_24479_, _24460_, _24443_);
  and (_24480_, _24479_, _24466_);
  or (_24481_, _24480_, _24478_);
  or (_24482_, _24481_, _24473_);
  or (_24483_, _24482_, _24465_);
  or (_24484_, _24483_, _24392_);
  nor (_24485_, _24413_, _24268_);
  and (_24486_, _24485_, _24319_);
  and (_24487_, _24452_, _24443_);
  and (_24488_, _24487_, _24486_);
  and (_24489_, _24413_, _24321_);
  nand (_24490_, _24367_, _24346_);
  nor (_24491_, _24490_, _24459_);
  and (_24492_, _24491_, _24445_);
  and (_24493_, _24492_, _24489_);
  or (_24494_, _24493_, _24488_);
  nor (_24495_, _24317_, _24294_);
  and (_24496_, _24495_, _24485_);
  and (_24497_, _24496_, _24471_);
  and (_24499_, _24460_, _24445_);
  and (_24500_, _24499_, _24321_);
  or (_24501_, _24500_, _24497_);
  and (_24502_, _24491_, _24486_);
  or (_24503_, _24502_, _24501_);
  or (_24505_, _24503_, _24494_);
  and (_24506_, _24468_, _24475_);
  and (_24507_, _24471_, _24321_);
  and (_24508_, _24479_, _24321_);
  or (_24509_, _24508_, _24507_);
  or (_24510_, _24509_, _24506_);
  and (_24511_, _24466_, _24391_);
  and (_24513_, _24471_, _24317_);
  or (_24514_, _24513_, _24511_);
  and (_24515_, _24393_, _24459_);
  nor (_24516_, _24490_, _24389_);
  and (_24517_, _24516_, _24443_);
  or (_24518_, _24517_, _24515_);
  and (_24519_, _24518_, _24486_);
  or (_24520_, _24519_, _24514_);
  or (_24521_, _24520_, _24510_);
  or (_24522_, _24521_, _24505_);
  or (_24523_, _24522_, _24484_);
  and (_24524_, _24523_, _22768_);
  and (_24525_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_24526_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_24527_, \oc8051_top_1.oc8051_decoder1.state [0], _22765_);
  and (_24528_, _24527_, _24526_);
  not (_24529_, _24528_);
  nor (_24531_, _24496_, _24416_);
  not (_24533_, _24531_);
  and (_24534_, _24533_, _24492_);
  and (_24536_, _24470_, _24418_);
  nor (_24537_, _24536_, _24534_);
  nor (_24538_, _24537_, _24529_);
  or (_24539_, _24538_, _24525_);
  or (_24540_, _24539_, _24524_);
  and (_26875_[0], _24540_, _22761_);
  and (_24541_, _23796_, _23648_);
  and (_24542_, _24541_, _23028_);
  and (_24544_, _24542_, _23791_);
  not (_24545_, _24542_);
  and (_24546_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_27274_, _24546_, _24544_);
  and (_24547_, _23651_, _23017_);
  and (_24549_, _24547_, _23791_);
  not (_24550_, _24547_);
  and (_24552_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_27311_, _24552_, _24549_);
  and (_24554_, _23838_, _23029_);
  and (_24555_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_27290_, _24555_, _24554_);
  and (_24556_, _23718_, _23029_);
  and (_24557_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_27289_, _24557_, _24556_);
  and (_24558_, _23805_, _23642_);
  and (_24559_, _24558_, _23017_);
  not (_24560_, _24559_);
  and (_24561_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_24562_, _24559_, _23589_);
  or (_27071_, _24562_, _24561_);
  or (_24564_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_24565_, _24564_, _22761_);
  nand (_24566_, _23889_, _23748_);
  and (_04534_, _24566_, _24565_);
  and (_24567_, _24117_, _23643_);
  and (_24568_, _24567_, _23755_);
  not (_24569_, _24567_);
  and (_24570_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or (_27087_, _24570_, _24568_);
  and (_24571_, _22982_, _22890_);
  and (_24572_, _24571_, _23805_);
  and (_24573_, _24572_, _23842_);
  and (_24574_, _24573_, _23676_);
  not (_24575_, _24573_);
  and (_24576_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or (_27162_, _24576_, _24574_);
  and (_24577_, _24118_, _23842_);
  and (_24578_, _24577_, _23838_);
  not (_24579_, _24577_);
  and (_24580_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or (_27232_, _24580_, _24578_);
  and (_24581_, _23635_, _23029_);
  and (_24582_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or (_27291_, _24582_, _24581_);
  and (_24583_, _23650_, _23598_);
  and (_24584_, _24583_, _24103_);
  and (_24585_, _24584_, _23676_);
  not (_24586_, _24584_);
  and (_24587_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or (_27125_, _24587_, _24585_);
  and (_24588_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_24590_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_24591_, _22770_, _24590_);
  or (_24592_, _24591_, _24588_);
  and (_26891_[9], _24592_, _22761_);
  and (_24593_, _24583_, _23594_);
  and (_24594_, _24593_, _23589_);
  not (_24595_, _24593_);
  and (_24596_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or (_27111_, _24596_, _24594_);
  and (_24597_, _23797_, _23643_);
  and (_24598_, _24597_, _23755_);
  not (_24599_, _24597_);
  and (_24600_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or (_27090_, _24600_, _24598_);
  and (_24601_, _24214_, _23791_);
  and (_24602_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or (_27072_, _24602_, _24601_);
  and (_24603_, _24214_, _23718_);
  and (_24604_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or (_27073_, _24604_, _24603_);
  and (_24605_, _24583_, _23017_);
  and (_24606_, _24605_, _23589_);
  not (_24607_, _24605_);
  and (_24608_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_27211_, _24608_, _24606_);
  and (_24610_, _24118_, _23649_);
  and (_24611_, _24610_, _23676_);
  not (_24612_, _24610_);
  and (_24613_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_27212_, _24613_, _24611_);
  and (_24614_, _24571_, _22933_);
  and (_24615_, _24614_, _23023_);
  and (_24616_, _24615_, _23641_);
  not (_24617_, _24616_);
  and (_24618_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and (_24619_, _24616_, _23635_);
  or (_27109_, _24619_, _24618_);
  and (_24620_, _24610_, _23791_);
  and (_24621_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_27213_, _24621_, _24620_);
  and (_24622_, _24583_, _23842_);
  and (_24623_, _24622_, _23982_);
  not (_24624_, _24622_);
  and (_24625_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_27201_, _24625_, _24623_);
  and (_24626_, _24622_, _23755_);
  and (_24627_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_27202_, _24627_, _24626_);
  and (_24628_, _22999_, _22981_);
  and (_24629_, _23879_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not (_24630_, _24629_);
  nor (_24631_, _24630_, _22913_);
  and (_24632_, _24631_, _22952_);
  and (_24633_, _24632_, _22890_);
  and (_24634_, _24633_, _24628_);
  and (_24635_, _23925_, _23812_);
  nor (_24636_, _23924_, _23918_);
  and (_24637_, _24636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_24638_, _24637_, _24635_);
  and (_24639_, _24638_, _24634_);
  not (_24640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_24641_, _24634_, _23012_);
  nor (_24642_, _24641_, _24640_);
  nor (_24643_, _22998_, _22951_);
  and (_24644_, _24643_, _23642_);
  and (_24645_, _23918_, _22913_);
  and (_24646_, _23924_, _23880_);
  and (_24647_, _24646_, _24645_);
  and (_24648_, _24647_, _24644_);
  or (_24649_, _24648_, _24642_);
  or (_24650_, _24649_, _24639_);
  nand (_24651_, _24648_, _23832_);
  and (_24652_, _24651_, _22761_);
  and (_06483_, _24652_, _24650_);
  not (_24653_, _24648_);
  and (_24654_, _24634_, _23992_);
  or (_24655_, _24654_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24656_, _24655_, _24653_);
  nand (_24657_, _24654_, _23522_);
  and (_24658_, _24657_, _24656_);
  and (_24659_, _24648_, _23709_);
  or (_24660_, _24659_, _24658_);
  and (_06503_, _24660_, _22761_);
  and (_24661_, _24634_, _23878_);
  or (_24662_, _24661_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24663_, _24662_, _24653_);
  nand (_24664_, _24661_, _23522_);
  and (_24665_, _24664_, _24663_);
  nor (_24666_, _24653_, _23784_);
  or (_24667_, _24666_, _24665_);
  and (_06526_, _24667_, _22761_);
  nand (_24668_, _24641_, _23985_);
  nor (_24669_, _24668_, _23522_);
  and (_24670_, _23880_, _22913_);
  and (_24671_, _23924_, _23918_);
  and (_24672_, _24671_, _24670_);
  and (_24673_, _24672_, _23642_);
  and (_24674_, _24673_, _24643_);
  and (_24675_, _24668_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_24676_, _24675_, _24674_);
  or (_24677_, _24676_, _24669_);
  nand (_24678_, _24648_, _23669_);
  and (_24679_, _24678_, _22761_);
  and (_06545_, _24679_, _24677_);
  and (_24680_, _24583_, _23803_);
  and (_24681_, _24680_, _23791_);
  not (_24682_, _24680_);
  and (_24683_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or (_27203_, _24683_, _24681_);
  and (_24684_, _24680_, _23838_);
  and (_24685_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or (_27204_, _24685_, _24684_);
  and (_24686_, _24680_, _23635_);
  and (_24687_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or (_27206_, _24687_, _24686_);
  and (_24688_, _23991_, _23918_);
  and (_24689_, _24688_, _24634_);
  nand (_24690_, _24689_, _23522_);
  or (_24691_, _24689_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_24692_, _24691_, _24653_);
  and (_24693_, _24692_, _24690_);
  nor (_24694_, _24653_, _23748_);
  or (_24695_, _24694_, _24693_);
  and (_06717_, _24695_, _22761_);
  and (_24696_, _24634_, _23919_);
  nand (_24697_, _24696_, _23522_);
  or (_24698_, _24696_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24699_, _24698_, _24653_);
  and (_24700_, _24699_, _24697_);
  nor (_24701_, _24653_, _23628_);
  or (_24702_, _24701_, _24700_);
  and (_06761_, _24702_, _22761_);
  and (_24703_, _24680_, _23755_);
  and (_24704_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or (_06852_, _24704_, _24703_);
  and (_24705_, _22951_, _22914_);
  and (_24706_, _24629_, _22890_);
  and (_24707_, _24706_, _24628_);
  and (_24708_, _24707_, _24705_);
  and (_24709_, _24708_, _23878_);
  or (_24710_, _24709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24711_, _22999_, _22951_);
  and (_24712_, _24711_, _23642_);
  and (_24713_, _23985_, _23012_);
  and (_24714_, _24713_, _23882_);
  and (_24715_, _24714_, _24712_);
  not (_24716_, _24715_);
  and (_24717_, _24716_, _24710_);
  nand (_24718_, _24709_, _23522_);
  and (_24719_, _24718_, _24717_);
  nor (_24720_, _24716_, _23784_);
  or (_24721_, _24720_, _24719_);
  and (_06907_, _24721_, _22761_);
  and (_24722_, _24583_, _23849_);
  and (_24723_, _24722_, _23718_);
  not (_24724_, _24722_);
  and (_24725_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or (_06935_, _24725_, _24723_);
  not (_24726_, _24708_);
  nor (_24728_, _23985_, _23012_);
  or (_24729_, _24728_, _24726_);
  and (_24730_, _24729_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  not (_24731_, _23986_);
  nor (_24732_, _24731_, _23522_);
  and (_24733_, _24732_, _24708_);
  or (_24734_, _24733_, _24730_);
  and (_24735_, _24708_, _23012_);
  and (_24736_, _24735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_24737_, _24736_, _24715_);
  or (_24738_, _24737_, _24734_);
  nand (_24739_, _24715_, _23914_);
  and (_24740_, _24739_, _22761_);
  and (_06955_, _24740_, _24738_);
  not (_24741_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor (_24742_, _24735_, _24741_);
  or (_24743_, _24742_, _24715_);
  and (_24744_, _24636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_24745_, _24744_, _24635_);
  and (_24746_, _24745_, _24708_);
  or (_24747_, _24746_, _24743_);
  nand (_24748_, _24715_, _23832_);
  and (_24749_, _24748_, _22761_);
  and (_07003_, _24749_, _24747_);
  and (_24750_, _24708_, _23992_);
  or (_24751_, _24750_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24752_, _24751_, _24716_);
  nand (_24753_, _24750_, _23522_);
  and (_24754_, _24753_, _24752_);
  and (_24755_, _24715_, _23709_);
  or (_24757_, _24755_, _24754_);
  and (_07039_, _24757_, _22761_);
  and (_24758_, _24708_, _24713_);
  or (_24759_, _24758_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24760_, _24759_, _24716_);
  nand (_24761_, _24758_, _23522_);
  and (_24762_, _24761_, _24760_);
  not (_24763_, _23669_);
  and (_24764_, _24715_, _24763_);
  or (_24765_, _24764_, _24762_);
  and (_07060_, _24765_, _22761_);
  and (_24766_, _24722_, _23838_);
  and (_24767_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or (_07105_, _24767_, _24766_);
  and (_24768_, _23802_, _23796_);
  and (_24769_, _24768_, _23643_);
  and (_24770_, _24769_, _23982_);
  not (_24771_, _24769_);
  and (_24772_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or (_07159_, _24772_, _24770_);
  and (_24773_, _24722_, _23635_);
  and (_24774_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or (_07183_, _24774_, _24773_);
  and (_24775_, _24722_, _23589_);
  and (_24776_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or (_07210_, _24776_, _24775_);
  and (_24777_, _24118_, _23017_);
  and (_24778_, _24777_, _23676_);
  not (_24779_, _24777_);
  and (_24780_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or (_27236_, _24780_, _24778_);
  and (_24782_, _24708_, _24688_);
  or (_24783_, _24782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_24784_, _24783_, _24716_);
  nand (_24785_, _24782_, _23522_);
  and (_24786_, _24785_, _24784_);
  nor (_24787_, _24716_, _23748_);
  or (_24788_, _24787_, _24786_);
  and (_07403_, _24788_, _22761_);
  and (_24789_, _24605_, _23791_);
  and (_24791_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_27210_, _24791_, _24789_);
  and (_24792_, _24605_, _23718_);
  and (_24793_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_07484_, _24793_, _24792_);
  and (_24794_, _24605_, _23982_);
  and (_24795_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_07516_, _24795_, _24794_);
  and (_24796_, _22998_, _22981_);
  and (_24797_, _24705_, _24706_);
  and (_24798_, _24797_, _24796_);
  and (_24799_, _24798_, _23986_);
  or (_24800_, _24799_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_24801_, _24714_, _23875_);
  not (_24802_, _24801_);
  and (_24803_, _24802_, _24800_);
  nand (_24804_, _24799_, _23522_);
  and (_24805_, _24804_, _24803_);
  nor (_24806_, _24802_, _23914_);
  or (_24807_, _24806_, _24805_);
  and (_07585_, _24807_, _22761_);
  and (_24808_, _24798_, _23992_);
  or (_24809_, _24808_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_24810_, _24809_, _24802_);
  nand (_24811_, _24808_, _23522_);
  and (_24812_, _24811_, _24810_);
  and (_24813_, _24801_, _23709_);
  or (_24814_, _24813_, _24812_);
  and (_07604_, _24814_, _22761_);
  and (_24815_, _24798_, _24713_);
  or (_24816_, _24815_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_24817_, _24816_, _24802_);
  nand (_24818_, _24815_, _23522_);
  and (_24819_, _24818_, _24817_);
  and (_24820_, _24801_, _24763_);
  or (_24821_, _24820_, _24819_);
  and (_07624_, _24821_, _22761_);
  and (_24822_, _24605_, _23635_);
  and (_24823_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_07690_, _24823_, _24822_);
  and (_24824_, _24610_, _23982_);
  and (_24825_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_07709_, _24825_, _24824_);
  and (_24826_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_24827_, _24559_, _23791_);
  or (_07729_, _24827_, _24826_);
  and (_24828_, _24610_, _23635_);
  and (_24829_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_27214_, _24829_, _24828_);
  and (_24830_, _24610_, _23589_);
  and (_24832_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_07831_, _24832_, _24830_);
  and (_24833_, _24118_, _24078_);
  and (_24834_, _24833_, _23676_);
  not (_24835_, _24833_);
  and (_24836_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or (_07877_, _24836_, _24834_);
  and (_24837_, _24833_, _23838_);
  and (_24838_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or (_27216_, _24838_, _24837_);
  and (_24839_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_24840_, _24559_, _23676_);
  or (_07957_, _24840_, _24839_);
  and (_24841_, _24833_, _23982_);
  and (_24842_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or (_07976_, _24842_, _24841_);
  and (_24843_, _23676_, _23601_);
  and (_24844_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or (_08021_, _24844_, _24843_);
  and (_24845_, _24833_, _23755_);
  and (_24846_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or (_08063_, _24846_, _24845_);
  and (_24847_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_24848_, _24847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_24849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_24850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_24851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _24850_);
  and (_24852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24853_, _24852_, _24851_);
  and (_24854_, _24853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_24855_, _24854_, _24849_);
  not (_24856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_24857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_24858_, _24857_, _24856_);
  nand (_24859_, _24858_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_24860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_24861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_24862_, _24861_, _24860_);
  and (_24863_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_24864_, _24863_);
  and (_24865_, _24864_, _24859_);
  and (_24866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24867_, _24866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_24868_, _24867_);
  and (_24869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24870_, _24869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24872_, _24871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_24873_, _24872_, _24870_);
  and (_24874_, _24873_, _24868_);
  and (_24875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_24876_, _24875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_24877_, _24876_);
  and (_24879_, _24877_, _24874_);
  and (_24880_, _24879_, _24865_);
  nor (_24881_, _24880_, _24855_);
  and (_24882_, _24849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not (_24883_, _24882_);
  not (_24884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_24885_, _24858_, _24884_);
  not (_24886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24887_, _24862_, _24886_);
  nor (_24888_, _24887_, _24885_);
  and (_24889_, _24875_, _24640_);
  not (_24890_, _24889_);
  and (_24891_, _24890_, _24888_);
  nor (_24892_, _24891_, _24883_);
  not (_24893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_24894_, _24866_, _24893_);
  not (_24895_, _24894_);
  not (_24896_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24897_, _24869_, _24896_);
  not (_24898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24899_, _24871_, _24898_);
  nor (_24900_, _24899_, _24897_);
  and (_24901_, _24900_, _24895_);
  nor (_24902_, _24901_, _24883_);
  nor (_24903_, _24902_, _24892_);
  nor (_24904_, _24903_, _24881_);
  nand (_24905_, _24904_, _24848_);
  and (_24906_, _24881_, _24848_);
  or (_24907_, _24906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_24908_, _24907_, _22761_);
  and (_08082_, _24908_, _24905_);
  and (_24909_, _24118_, _23962_);
  and (_24910_, _24909_, _23718_);
  not (_24911_, _24909_);
  and (_24912_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or (_08181_, _24912_, _24910_);
  and (_24913_, _24909_, _23982_);
  and (_24914_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or (_08224_, _24914_, _24913_);
  and (_24915_, _24909_, _23755_);
  and (_24916_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or (_27218_, _24916_, _24915_);
  and (_24917_, _24909_, _23589_);
  and (_24918_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or (_27219_, _24918_, _24917_);
  nor (_24919_, _24847_, _24850_);
  and (_24920_, _24919_, _24881_);
  not (_24921_, _24919_);
  or (_24922_, _24921_, _24903_);
  and (_24923_, _24922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_24924_, _24923_, _24920_);
  and (_08337_, _24924_, _22761_);
  and (_24925_, _24118_, _23594_);
  and (_24926_, _24925_, _23791_);
  not (_24927_, _24925_);
  and (_24928_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_08374_, _24928_, _24926_);
  and (_24929_, _24925_, _23838_);
  and (_24930_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_08392_, _24930_, _24929_);
  and (_24931_, _23718_, _23601_);
  and (_24932_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or (_08411_, _24932_, _24931_);
  not (_24933_, _24881_);
  and (_24934_, _24903_, _24933_);
  nor (_24935_, _24934_, _24847_);
  not (_24936_, _24935_);
  and (_24937_, _24936_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_24938_, _24847_);
  nor (_24939_, _24859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24940_, _24939_, _24876_);
  not (_24941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_24942_, _24863_, _24850_);
  or (_24943_, _24942_, _24941_);
  nand (_24944_, _24943_, _24940_);
  and (_24945_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24946_, _24945_, _24877_);
  and (_24947_, _24946_, _24944_);
  or (_24948_, _24947_, _24872_);
  not (_24949_, _24870_);
  not (_24950_, _24872_);
  or (_24951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _24850_);
  or (_24952_, _24951_, _24950_);
  and (_24953_, _24952_, _24949_);
  and (_24954_, _24953_, _24948_);
  and (_24955_, _24945_, _24870_);
  or (_24956_, _24955_, _24867_);
  or (_24957_, _24956_, _24954_);
  or (_24958_, _24951_, _24868_);
  and (_24959_, _24958_, _24881_);
  and (_24960_, _24959_, _24957_);
  or (_24961_, _24951_, _24895_);
  and (_24962_, _24885_, _24850_);
  nor (_24963_, _24962_, _24889_);
  and (_24964_, _24887_, _24850_);
  or (_24965_, _24964_, _24941_);
  nand (_24966_, _24965_, _24963_);
  or (_24967_, _24945_, _24890_);
  and (_24968_, _24967_, _24966_);
  or (_24969_, _24968_, _24899_);
  not (_24970_, _24897_);
  not (_24971_, _24899_);
  or (_24972_, _24951_, _24971_);
  and (_24973_, _24972_, _24970_);
  and (_24974_, _24973_, _24969_);
  and (_24975_, _24945_, _24897_);
  or (_24976_, _24975_, _24894_);
  or (_24977_, _24976_, _24974_);
  and (_24978_, _24977_, _24904_);
  and (_24979_, _24978_, _24961_);
  or (_24980_, _24979_, _24960_);
  and (_24981_, _24980_, _24938_);
  or (_24982_, _24981_, _24937_);
  and (_08453_, _24982_, _22761_);
  and (_24983_, _24925_, _23635_);
  and (_24984_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_08475_, _24984_, _24983_);
  nand (_24985_, _24934_, _24848_);
  nor (_24986_, _24881_, _24847_);
  or (_24987_, _24986_, _24850_);
  and (_24988_, _24987_, _22761_);
  and (_08562_, _24988_, _24985_);
  and (_24989_, _24925_, _23755_);
  and (_24990_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_08595_, _24990_, _24989_);
  and (_24991_, _24118_, _24103_);
  and (_24992_, _24991_, _23791_);
  not (_24993_, _24991_);
  and (_24994_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_27221_, _24994_, _24992_);
  and (_24995_, _24991_, _23838_);
  and (_24996_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_08658_, _24996_, _24995_);
  not (_24997_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_24998_, _24935_, _24997_);
  or (_24999_, _24877_, _24872_);
  and (_25000_, _24999_, _24949_);
  and (_25001_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _24850_);
  or (_25002_, _25001_, _25000_);
  and (_25003_, _24863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25004_, _25003_, _24997_);
  nor (_25005_, _24859_, _24850_);
  nor (_25006_, _25005_, _24876_);
  nand (_25008_, _25006_, _24873_);
  or (_25009_, _25008_, _25004_);
  and (_25010_, _25009_, _25002_);
  or (_25011_, _25010_, _24867_);
  or (_25012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25013_, _24950_, _24870_);
  and (_25014_, _25013_, _24868_);
  or (_25015_, _25014_, _25012_);
  and (_25016_, _25015_, _24881_);
  and (_25017_, _25016_, _25011_);
  and (_25018_, _24885_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25019_, _25018_, _24889_);
  and (_25020_, _24887_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25021_, _25020_, _24997_);
  nand (_25023_, _25021_, _25019_);
  or (_25024_, _25001_, _24890_);
  and (_25025_, _25024_, _25023_);
  or (_25026_, _25025_, _24899_);
  or (_25027_, _25012_, _24971_);
  and (_25028_, _25027_, _24970_);
  and (_25029_, _25028_, _25026_);
  and (_25030_, _25001_, _24897_);
  or (_25031_, _25030_, _24894_);
  or (_25032_, _25031_, _25029_);
  and (_25033_, _24904_, _24895_);
  and (_25034_, _25012_, _24904_);
  or (_25035_, _25034_, _25033_);
  and (_25036_, _25035_, _25032_);
  or (_25037_, _25036_, _25017_);
  and (_25038_, _25037_, _24938_);
  or (_25039_, _25038_, _24998_);
  and (_08759_, _25039_, _22761_);
  and (_25040_, _24991_, _23635_);
  and (_25041_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_08780_, _25041_, _25040_);
  and (_25042_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_25043_, _24559_, _23838_);
  or (_08829_, _25043_, _25042_);
  and (_25044_, _24991_, _23755_);
  and (_25045_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_08852_, _25045_, _25044_);
  and (_25046_, _24118_, _23863_);
  and (_25047_, _25046_, _23676_);
  not (_25048_, _25046_);
  and (_25049_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or (_08972_, _25049_, _25047_);
  and (_25050_, _25046_, _23718_);
  and (_25051_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or (_08996_, _25051_, _25050_);
  and (_25052_, _25046_, _23982_);
  and (_25053_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or (_09029_, _25053_, _25052_);
  and (_25054_, _25046_, _23635_);
  and (_25055_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or (_09049_, _25055_, _25054_);
  and (_25056_, _24847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_25058_, _25056_, _24935_);
  and (_09078_, _25058_, _22761_);
  or (_25059_, _24899_, _24889_);
  nor (_25060_, _24897_, _24894_);
  nand (_25061_, _25060_, _24882_);
  or (_25063_, _25061_, _25059_);
  or (_25064_, _25063_, _24888_);
  nor (_25066_, _25064_, _24881_);
  and (_25067_, _24847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_25068_, _24855_, _24847_);
  not (_25069_, _24865_);
  and (_25070_, _24879_, _25069_);
  and (_25071_, _25070_, _25068_);
  or (_25072_, _25071_, _25067_);
  or (_25073_, _25072_, _25066_);
  and (_09104_, _25073_, _22761_);
  and (_25074_, _24888_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_25075_, _25074_, _25059_);
  and (_25076_, _25075_, _25060_);
  and (_25077_, _25076_, _24904_);
  nor (_25078_, _24870_, _24867_);
  or (_25079_, _24876_, _24872_);
  and (_25080_, _24865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_25081_, _25080_, _25079_);
  and (_25082_, _25081_, _25078_);
  and (_25083_, _25082_, _24881_);
  or (_25084_, _25083_, _25077_);
  or (_25085_, _25084_, _24847_);
  or (_25086_, _24938_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_25087_, _25086_, _22761_);
  and (_09132_, _25087_, _25085_);
  and (_25088_, _24118_, _23641_);
  and (_25089_, _25088_, _23676_);
  not (_25090_, _25088_);
  and (_25091_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or (_27223_, _25091_, _25089_);
  nor (_25092_, _24887_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_25093_, _25092_, _24885_);
  or (_25094_, _25093_, _24889_);
  and (_25095_, _25094_, _24971_);
  or (_25097_, _25095_, _24897_);
  and (_25098_, _25097_, _25033_);
  or (_25099_, _24863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25100_, _25099_, _24859_);
  or (_25101_, _25100_, _24876_);
  and (_25102_, _25101_, _24950_);
  or (_25103_, _25102_, _24870_);
  and (_25104_, _24881_, _24868_);
  and (_25105_, _25104_, _25103_);
  or (_25106_, _25105_, _24847_);
  or (_25107_, _25106_, _25098_);
  not (_25108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nand (_25109_, _24847_, _25108_);
  and (_25110_, _25109_, _22761_);
  and (_09188_, _25110_, _25107_);
  and (_25111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _22761_);
  and (_09242_, _25111_, _24847_);
  and (_25113_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_25115_, _24559_, _23982_);
  or (_09285_, _25115_, _25113_);
  nor (_25116_, _22951_, _22914_);
  and (_25117_, _25116_, _22890_);
  and (_25118_, _25117_, _24628_);
  and (_25119_, _25118_, _23925_);
  nand (_25120_, _25119_, _23522_);
  or (_25121_, _25119_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_25122_, _25121_, _24629_);
  and (_25123_, _25122_, _25120_);
  and (_25124_, _25118_, _24713_);
  nand (_25125_, _25124_, _23832_);
  or (_25126_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_25127_, _25126_, _23880_);
  and (_25128_, _25127_, _25125_);
  not (_25129_, _23879_);
  and (_25130_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_25131_, _25130_, rst);
  or (_25132_, _25131_, _25128_);
  or (_09305_, _25132_, _25123_);
  and (_25133_, _25088_, _23791_);
  and (_25134_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or (_09325_, _25134_, _25133_);
  and (_25135_, _25118_, _23992_);
  nand (_25136_, _25135_, _23522_);
  or (_25137_, _25135_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_25138_, _25137_, _24629_);
  and (_25139_, _25138_, _25136_);
  not (_25140_, _25124_);
  or (_25141_, _25140_, _23709_);
  or (_25142_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_25143_, _25142_, _23880_);
  and (_25144_, _25143_, _25141_);
  and (_25145_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_25146_, _25145_, rst);
  or (_25147_, _25146_, _25144_);
  or (_09347_, _25147_, _25139_);
  and (_25148_, _25118_, _23878_);
  nand (_25149_, _25148_, _23522_);
  or (_25150_, _25148_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_25151_, _25150_, _24629_);
  and (_25152_, _25151_, _25149_);
  nand (_25153_, _25124_, _23784_);
  or (_25154_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_25155_, _25154_, _23880_);
  and (_25156_, _25155_, _25153_);
  and (_25157_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_25158_, _25157_, rst);
  or (_25159_, _25158_, _25156_);
  or (_09369_, _25159_, _25152_);
  nand (_25160_, _25124_, _23522_);
  or (_25161_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_25162_, _25161_, _24629_);
  and (_25163_, _25162_, _25160_);
  nand (_25164_, _25124_, _23669_);
  and (_25165_, _25164_, _23880_);
  and (_25166_, _25165_, _25161_);
  not (_25167_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_25168_, _23879_, _25167_);
  or (_25169_, _25168_, rst);
  or (_25170_, _25169_, _25166_);
  or (_09390_, _25170_, _25163_);
  and (_25171_, _25088_, _23838_);
  and (_25172_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or (_27225_, _25172_, _25171_);
  and (_25173_, _25088_, _23635_);
  and (_25174_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or (_09452_, _25174_, _25173_);
  and (_25175_, _25088_, _23589_);
  and (_25176_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or (_09490_, _25176_, _25175_);
  and (_25177_, _25118_, _24688_);
  nand (_25178_, _25177_, _23522_);
  or (_25179_, _25177_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_25180_, _25179_, _24629_);
  and (_25181_, _25180_, _25178_);
  nand (_25182_, _25124_, _23748_);
  or (_25183_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_25184_, _25183_, _23880_);
  and (_25185_, _25184_, _25182_);
  and (_25186_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_25187_, _25186_, rst);
  or (_25188_, _25187_, _25185_);
  or (_09507_, _25188_, _25181_);
  and (_25189_, _24119_, _23676_);
  and (_25190_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_09607_, _25190_, _25189_);
  and (_25191_, _25118_, _23919_);
  nand (_25192_, _25191_, _23522_);
  or (_25193_, _25191_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_25194_, _25193_, _24629_);
  and (_25195_, _25194_, _25192_);
  nand (_25196_, _25124_, _23628_);
  or (_25197_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_25198_, _25197_, _23880_);
  and (_25199_, _25198_, _25196_);
  and (_25200_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_25201_, _25200_, rst);
  or (_25202_, _25201_, _25199_);
  or (_09650_, _25202_, _25195_);
  and (_25203_, _24119_, _23718_);
  and (_25204_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_09750_, _25204_, _25203_);
  and (_25205_, _24119_, _23982_);
  and (_25206_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_09775_, _25206_, _25205_);
  and (_25207_, _22951_, _22913_);
  and (_25208_, _25207_, _22890_);
  and (_25209_, _25208_, _24628_);
  and (_25210_, _25209_, _23878_);
  nand (_25211_, _25210_, _23522_);
  or (_25212_, _25210_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_25213_, _25212_, _24629_);
  and (_25214_, _25213_, _25211_);
  and (_25215_, _24713_, _22913_);
  and (_25216_, _25215_, _24712_);
  nand (_25217_, _25216_, _23784_);
  or (_25218_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_25219_, _25218_, _23880_);
  and (_25220_, _25219_, _25217_);
  and (_25221_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_25222_, _25221_, rst);
  or (_25223_, _25222_, _25220_);
  or (_09827_, _25223_, _25214_);
  and (_25224_, _25209_, _23919_);
  nand (_25226_, _25224_, _23522_);
  or (_25227_, _25224_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_25228_, _25227_, _24629_);
  and (_25230_, _25228_, _25226_);
  nand (_25231_, _25216_, _23628_);
  or (_25233_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_25234_, _25233_, _23880_);
  and (_25235_, _25234_, _25231_);
  and (_25236_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_25237_, _25236_, rst);
  or (_25238_, _25237_, _25235_);
  or (_09875_, _25238_, _25230_);
  and (_25239_, _25209_, _23986_);
  nand (_25240_, _25239_, _23522_);
  or (_25241_, _25239_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_25242_, _25241_, _24629_);
  and (_25243_, _25242_, _25240_);
  nand (_25244_, _25216_, _23914_);
  or (_25245_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_25246_, _25245_, _23880_);
  and (_25247_, _25246_, _25244_);
  and (_25248_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_25249_, _25248_, rst);
  or (_25250_, _25249_, _25247_);
  or (_09902_, _25250_, _25243_);
  and (_25251_, _25209_, _23925_);
  nand (_25252_, _25251_, _23522_);
  or (_25253_, _25251_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_25254_, _25253_, _24629_);
  and (_25255_, _25254_, _25252_);
  nand (_25256_, _25216_, _23832_);
  or (_25257_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_25258_, _25257_, _23880_);
  and (_25259_, _25258_, _25256_);
  and (_25260_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_25261_, _25260_, rst);
  or (_25262_, _25261_, _25259_);
  or (_09928_, _25262_, _25255_);
  and (_25263_, _25209_, _23992_);
  nand (_25264_, _25263_, _23522_);
  or (_25265_, _25263_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_25266_, _25265_, _24629_);
  and (_25267_, _25266_, _25264_);
  not (_25268_, _23709_);
  nand (_25269_, _25216_, _25268_);
  or (_25270_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_25271_, _25270_, _23880_);
  and (_25272_, _25271_, _25269_);
  and (_25273_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_25274_, _25273_, rst);
  or (_25275_, _25274_, _25272_);
  or (_09956_, _25275_, _25267_);
  and (_25276_, _25209_, _24713_);
  nand (_25277_, _25276_, _23522_);
  or (_25278_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_25279_, _25278_, _24629_);
  and (_25280_, _25279_, _25277_);
  nand (_25281_, _25216_, _23669_);
  and (_25282_, _25281_, _23880_);
  and (_25283_, _25282_, _25278_);
  not (_25284_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_25285_, _23879_, _25284_);
  or (_25286_, _25285_, rst);
  or (_25288_, _25286_, _25283_);
  or (_09994_, _25288_, _25280_);
  and (_25289_, _24584_, _23718_);
  and (_25290_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or (_27126_, _25290_, _25289_);
  and (_25291_, _24584_, _23791_);
  and (_25292_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or (_10167_, _25292_, _25291_);
  and (_25294_, _24558_, _23849_);
  not (_25295_, _25294_);
  and (_25296_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and (_25297_, _25294_, _23982_);
  or (_10243_, _25297_, _25296_);
  and (_25298_, _24573_, _23718_);
  and (_25299_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or (_10254_, _25299_, _25298_);
  and (_25301_, _23854_, _23643_);
  and (_25302_, _25301_, _23791_);
  not (_25303_, _25301_);
  and (_25304_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_10287_, _25304_, _25302_);
  and (_25305_, _24593_, _23718_);
  and (_25306_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or (_10331_, _25306_, _25305_);
  and (_25307_, _24593_, _23791_);
  and (_25308_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or (_10354_, _25308_, _25307_);
  and (_25309_, _25117_, _24796_);
  and (_25310_, _25309_, _23925_);
  nand (_25311_, _25310_, _23522_);
  or (_25312_, _25310_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_25313_, _25312_, _24629_);
  and (_25314_, _25313_, _25311_);
  and (_25315_, _22998_, _22952_);
  and (_25316_, _25315_, _23642_);
  and (_25317_, _25316_, _25215_);
  nand (_25319_, _25317_, _23832_);
  or (_25320_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_25321_, _25320_, _23880_);
  and (_25322_, _25321_, _25319_);
  and (_25323_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_25324_, _25323_, rst);
  or (_25325_, _25324_, _25322_);
  or (_10378_, _25325_, _25314_);
  and (_25327_, _25309_, _23992_);
  nand (_25328_, _25327_, _23522_);
  or (_25329_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_25331_, _25329_, _24629_);
  and (_25332_, _25331_, _25328_);
  not (_25333_, _25317_);
  or (_25334_, _25333_, _23709_);
  or (_25335_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_25336_, _25335_, _23880_);
  and (_25337_, _25336_, _25334_);
  and (_25338_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_25339_, _25338_, rst);
  or (_25340_, _25339_, _25337_);
  or (_10401_, _25340_, _25332_);
  and (_25341_, _25309_, _23878_);
  nand (_25342_, _25341_, _23522_);
  or (_25343_, _25341_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_25344_, _25343_, _24629_);
  and (_25346_, _25344_, _25342_);
  nand (_25348_, _25317_, _23784_);
  or (_25349_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_25351_, _25349_, _23880_);
  and (_25352_, _25351_, _25348_);
  and (_25353_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_25354_, _25353_, rst);
  or (_25355_, _25354_, _25352_);
  or (_10424_, _25355_, _25346_);
  and (_25356_, _25309_, _24713_);
  nand (_25357_, _25356_, _23522_);
  or (_25358_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_25359_, _25358_, _24629_);
  and (_25360_, _25359_, _25357_);
  nand (_25361_, _25317_, _23669_);
  and (_25362_, _25361_, _23880_);
  and (_25363_, _25362_, _25358_);
  not (_25364_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_25365_, _23879_, _25364_);
  or (_25366_, _25365_, rst);
  or (_25367_, _25366_, _25363_);
  or (_10447_, _25367_, _25360_);
  and (_25368_, _24593_, _23676_);
  and (_25369_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or (_10469_, _25369_, _25368_);
  and (_25370_, _25309_, _24688_);
  nand (_25371_, _25370_, _23522_);
  or (_25372_, _25370_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_25373_, _25372_, _24629_);
  and (_25374_, _25373_, _25371_);
  nand (_25375_, _25317_, _23748_);
  or (_25376_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_25377_, _25376_, _23880_);
  and (_25378_, _25377_, _25375_);
  and (_25379_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_25380_, _25379_, rst);
  or (_25381_, _25380_, _25378_);
  or (_10777_, _25381_, _25374_);
  and (_25382_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and (_25383_, _25294_, _23755_);
  or (_10904_, _25383_, _25382_);
  and (_25384_, _25309_, _23919_);
  nand (_25385_, _25384_, _23522_);
  or (_25386_, _25384_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_25387_, _25386_, _24629_);
  and (_25388_, _25387_, _25385_);
  nand (_25389_, _25317_, _23628_);
  or (_25390_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_25391_, _25390_, _23880_);
  and (_25392_, _25391_, _25389_);
  and (_25394_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_25395_, _25394_, rst);
  or (_25397_, _25395_, _25392_);
  or (_10980_, _25397_, _25388_);
  and (_25398_, _24593_, _23635_);
  and (_25399_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or (_11031_, _25399_, _25398_);
  and (_25400_, _24078_, _23599_);
  and (_25401_, _25400_, _23755_);
  not (_25402_, _25400_);
  and (_25403_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_11111_, _25403_, _25401_);
  and (_25405_, _24593_, _23982_);
  and (_25406_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or (_11143_, _25406_, _25405_);
  and (_25407_, _25208_, _24796_);
  and (_25408_, _25407_, _23992_);
  nand (_25409_, _25408_, _23522_);
  or (_25410_, _25408_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25411_, _25410_, _24629_);
  and (_25412_, _25411_, _25409_);
  and (_25413_, _25215_, _23875_);
  not (_25414_, _25413_);
  or (_25415_, _25414_, _23709_);
  or (_25416_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25417_, _25416_, _23880_);
  and (_25418_, _25417_, _25415_);
  and (_25419_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_25420_, _25419_, rst);
  or (_25422_, _25420_, _25418_);
  or (_11331_, _25422_, _25412_);
  and (_25423_, _25407_, _23878_);
  nand (_25424_, _25423_, _23522_);
  or (_25425_, _25423_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_25426_, _25425_, _24629_);
  and (_25428_, _25426_, _25424_);
  nand (_25429_, _25413_, _23784_);
  or (_25430_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_25431_, _25430_, _23880_);
  and (_25432_, _25431_, _25429_);
  and (_25433_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_25434_, _25433_, rst);
  or (_25435_, _25434_, _25432_);
  or (_11355_, _25435_, _25428_);
  and (_25436_, _25407_, _24713_);
  nand (_25437_, _25436_, _23522_);
  or (_25438_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_25440_, _25438_, _24629_);
  and (_25441_, _25440_, _25437_);
  nand (_25442_, _25413_, _23669_);
  and (_25443_, _25438_, _23880_);
  and (_25444_, _25443_, _25442_);
  not (_25445_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_25446_, _23879_, _25445_);
  or (_25447_, _25446_, rst);
  or (_25448_, _25447_, _25444_);
  or (_11382_, _25448_, _25441_);
  and (_25449_, _25400_, _23589_);
  and (_25450_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_11495_, _25450_, _25449_);
  and (_25451_, _25407_, _23919_);
  nand (_25452_, _25451_, _23522_);
  or (_25453_, _25451_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25454_, _25453_, _24629_);
  and (_25455_, _25454_, _25452_);
  nand (_25456_, _25413_, _23628_);
  or (_25457_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25458_, _25457_, _23880_);
  and (_25459_, _25458_, _25456_);
  and (_25461_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_25462_, _25461_, rst);
  or (_25463_, _25462_, _25459_);
  or (_11654_, _25463_, _25455_);
  and (_25464_, _24558_, _23803_);
  not (_25465_, _25464_);
  and (_25466_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  and (_25467_, _25464_, _23589_);
  or (_11687_, _25467_, _25466_);
  and (_25468_, _24583_, _23962_);
  and (_25469_, _25468_, _23982_);
  not (_25470_, _25468_);
  and (_25471_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_11746_, _25471_, _25469_);
  and (_25472_, _25407_, _24688_);
  nand (_25473_, _25472_, _23522_);
  or (_25474_, _25472_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25476_, _25474_, _24629_);
  and (_25477_, _25476_, _25473_);
  nand (_25478_, _25413_, _23748_);
  or (_25479_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25481_, _25479_, _23880_);
  and (_25482_, _25481_, _25478_);
  and (_25483_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_25484_, _25483_, rst);
  or (_25485_, _25484_, _25482_);
  or (_11786_, _25485_, _25477_);
  not (_25486_, _25407_);
  or (_25487_, _25486_, _24728_);
  and (_25488_, _25487_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25489_, _23012_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_25491_, _25489_, _24732_);
  and (_25492_, _25491_, _25407_);
  or (_25493_, _25492_, _25488_);
  and (_25494_, _25493_, _24629_);
  nand (_25495_, _25413_, _23914_);
  or (_25496_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25497_, _25496_, _23880_);
  and (_25498_, _25497_, _25495_);
  and (_25499_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_25501_, _25499_, rst);
  or (_25502_, _25501_, _25498_);
  or (_11811_, _25502_, _25494_);
  and (_25503_, _25400_, _23718_);
  and (_25504_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_11935_, _25504_, _25503_);
  and (_25505_, _25468_, _23838_);
  and (_25506_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_12030_, _25506_, _25505_);
  and (_25507_, _25468_, _23589_);
  and (_25508_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_27096_, _25508_, _25507_);
  and (_25509_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and (_25510_, _25294_, _23791_);
  or (_12238_, _25510_, _25509_);
  and (_25512_, _25468_, _23755_);
  and (_25513_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_27095_, _25513_, _25512_);
  and (_25515_, _25468_, _23635_);
  and (_25516_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_12299_, _25516_, _25515_);
  and (_25517_, _24103_, _23028_);
  and (_25518_, _25517_, _23589_);
  not (_25519_, _25517_);
  and (_25520_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_13746_, _25520_, _25518_);
  and (_25521_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and (_25522_, _25464_, _23838_);
  or (_13781_, _25522_, _25521_);
  and (_25523_, _22929_, _22856_);
  and (_25525_, _23878_, _22913_);
  and (_25526_, _25315_, _23596_);
  and (_25528_, _25526_, _25525_);
  and (_25529_, _25528_, _25523_);
  and (_25530_, _25529_, _23589_);
  not (_25531_, _25529_);
  and (_25532_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_13902_, _25532_, _25530_);
  and (_25533_, _25529_, _23755_);
  and (_25534_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_14374_, _25534_, _25533_);
  and (_25536_, _23962_, _23599_);
  and (_25537_, _25536_, _23982_);
  not (_25538_, _25536_);
  and (_25539_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_14495_, _25539_, _25537_);
  and (_25540_, _25529_, _23635_);
  and (_25541_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_14596_, _25541_, _25540_);
  and (_25542_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and (_25543_, _25464_, _23982_);
  or (_14645_, _25543_, _25542_);
  and (_25544_, _23798_, _23755_);
  and (_25546_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or (_14741_, _25546_, _25544_);
  nor (_25547_, _22768_, _23206_);
  and (_25548_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_25549_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_25550_, _25549_, _25548_);
  and (_25551_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_25552_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_25553_, _25552_, _25551_);
  and (_25554_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_25555_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_25556_, _25555_, _25554_);
  and (_25558_, _25556_, _25553_);
  and (_25559_, _25558_, _25550_);
  and (_25561_, _22768_, _24270_);
  not (_25562_, _25561_);
  nor (_25564_, _25562_, _25559_);
  nor (_25565_, _25564_, _25547_);
  nor (_26896_[2], _25565_, rst);
  not (_25566_, _22768_);
  and (_25568_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_25569_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_25570_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_25571_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_25572_, _25571_, _25570_);
  and (_25573_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_25574_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_25575_, _25574_, _25573_);
  or (_25576_, _25575_, _25572_);
  and (_25577_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_25578_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_25579_, _25578_, _25577_);
  or (_25580_, _25579_, _25576_);
  and (_25581_, _25580_, _24270_);
  or (_25582_, _25581_, _25569_);
  and (_25583_, _25582_, _22768_);
  nor (_25584_, _25583_, _25568_);
  nor (_26906_[4], _25584_, rst);
  and (_25585_, _25468_, _23791_);
  and (_25586_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_16909_, _25586_, _25585_);
  and (_25587_, _25468_, _23676_);
  and (_25588_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_17026_, _25588_, _25587_);
  and (_25589_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_25590_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_25591_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_25592_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_25593_, _25592_, _25591_);
  and (_25594_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_25595_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_25596_, _25595_, _25594_);
  and (_25597_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_25598_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_25599_, _25598_, _25597_);
  and (_25600_, _25599_, _25596_);
  and (_25601_, _25600_, _25593_);
  nor (_25602_, _25601_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_25603_, _25602_, _25590_);
  nor (_25604_, _25603_, _25566_);
  nor (_25605_, _25604_, _25589_);
  nor (_26906_[7], _25605_, rst);
  and (_25606_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and (_25607_, _25464_, _23635_);
  or (_17209_, _25607_, _25606_);
  and (_25608_, _25526_, _25215_);
  and (_25609_, _25608_, _25523_);
  and (_25610_, _25609_, _23589_);
  not (_25611_, _25609_);
  and (_25612_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or (_17708_, _25612_, _25610_);
  and (_25613_, _24496_, _24491_);
  nor (_25614_, _25613_, _24536_);
  and (_25615_, _22768_, _22761_);
  not (_25616_, _25615_);
  or (_26871_[1], _25616_, _25614_);
  nor (_25617_, _25611_, _23748_);
  and (_25618_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or (_18030_, _25618_, _25617_);
  and (_25619_, _24558_, _23842_);
  not (_25620_, _25619_);
  and (_25621_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_25622_, _25619_, _23589_);
  or (_27067_, _25622_, _25621_);
  and (_25625_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_25627_, _25619_, _23755_);
  or (_27066_, _25627_, _25625_);
  nor (_25628_, _22768_, _23227_);
  and (_25629_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_25630_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_25631_, _25630_, _25629_);
  and (_25632_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_25633_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_25634_, _25633_, _25632_);
  and (_25635_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_25636_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_25637_, _25636_, _25635_);
  and (_25638_, _25637_, _25634_);
  and (_25639_, _25638_, _25631_);
  nor (_25640_, _25639_, _25562_);
  nor (_25641_, _25640_, _25628_);
  nor (_26896_[1], _25641_, rst);
  and (_25642_, _25529_, _23791_);
  and (_25643_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_18475_, _25643_, _25642_);
  and (_25644_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_25646_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_25647_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_25650_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_25651_, _25650_, _25647_);
  and (_25652_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_25653_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_25654_, _25653_, _25652_);
  and (_25655_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_25656_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_25657_, _25656_, _25655_);
  and (_25658_, _25657_, _25654_);
  and (_25659_, _25658_, _25651_);
  nor (_25660_, _25659_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_25661_, _25660_, _25646_);
  nor (_25662_, _25661_, _25566_);
  nor (_25663_, _25662_, _25644_);
  nor (_26906_[3], _25663_, rst);
  and (_25664_, _23798_, _23635_);
  and (_25665_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or (_18556_, _25665_, _25664_);
  and (_25666_, _24571_, _23874_);
  and (_25667_, _25666_, _23987_);
  and (_25668_, _25667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_25669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_25670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_25671_, _25670_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_25672_, _25671_, _25669_);
  not (_25673_, _25672_);
  and (_25674_, _25673_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_25675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_25676_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_25677_, _25676_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_25678_, _25677_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_25679_, _25678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_25680_, _25679_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_25681_, _25680_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_25682_, _25681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_25683_, _25682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_25685_, _25683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_25687_, _25685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_25688_, _25687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_25689_, _25688_, _25675_);
  and (_25690_, _25689_, _25674_);
  nand (_25691_, _25690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_25692_, _25690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_25693_, _25692_, _25691_);
  not (_25694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor (_25695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_25696_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_25697_, _25696_, _25695_);
  and (_25699_, _25697_, _25694_);
  and (_25700_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_25701_, _25700_, _25689_);
  and (_25702_, _25695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_25703_, _25702_);
  and (_25704_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_25705_, _25704_, _25674_);
  and (_25706_, _25705_, _25701_);
  or (_25707_, _25706_, _25699_);
  or (_25708_, _25707_, _25693_);
  not (_25709_, _25699_);
  or (_25710_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_25711_, _25666_, _23920_);
  nor (_25712_, _25711_, _25667_);
  and (_25713_, _25712_, _25710_);
  and (_25715_, _25713_, _25708_);
  not (_25716_, _25711_);
  nor (_25717_, _25716_, _23748_);
  or (_25718_, _25717_, _25715_);
  or (_25720_, _25718_, _25668_);
  and (_18587_, _25720_, _22761_);
  and (_25721_, _25529_, _23718_);
  and (_25722_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_18678_, _25722_, _25721_);
  nor (_25723_, _22768_, _23050_);
  and (_25724_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_25725_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_25727_, _25725_, _25724_);
  and (_25728_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_25729_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_25730_, _25729_, _25728_);
  and (_25731_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_25733_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_25734_, _25733_, _25731_);
  and (_25735_, _25734_, _25730_);
  and (_25736_, _25735_, _25727_);
  nor (_25738_, _25736_, _25562_);
  nor (_25739_, _25738_, _25723_);
  nor (_26896_[7], _25739_, rst);
  and (_25740_, _23982_, _23798_);
  and (_25741_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or (_19697_, _25741_, _25740_);
  and (_25742_, _23863_, _23028_);
  and (_25743_, _25742_, _23676_);
  not (_25744_, _25742_);
  and (_25745_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_19788_, _25745_, _25743_);
  and (_25746_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and (_25748_, _25464_, _23676_);
  or (_27068_, _25748_, _25746_);
  nor (_25749_, _25611_, _23784_);
  and (_25750_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or (_19939_, _25750_, _25749_);
  and (_25751_, _25609_, _24763_);
  and (_25752_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or (_20400_, _25752_, _25751_);
  nor (_25753_, _22768_, _23266_);
  and (_25754_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_25755_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_25756_, _25755_, _25754_);
  and (_25758_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_25759_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_25760_, _25759_, _25758_);
  and (_25761_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_25762_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_25763_, _25762_, _25761_);
  and (_25764_, _25763_, _25760_);
  and (_25765_, _25764_, _25756_);
  nor (_25766_, _25765_, _25562_);
  nor (_25767_, _25766_, _25753_);
  nor (_26896_[0], _25767_, rst);
  nor (_26869_[7], _24340_, rst);
  and (_26894_[0], _24413_, _22761_);
  and (_26894_[1], _24268_, _22761_);
  and (_26894_[2], _24294_, _22761_);
  and (_25769_, _24670_, _24713_);
  and (_25770_, _25769_, _25315_);
  and (_25771_, _25770_, _24571_);
  not (_25772_, _25771_);
  and (_25773_, _25772_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_25774_, _25315_, _24571_);
  and (_25775_, _25774_, _25769_);
  not (_25776_, _25775_);
  nor (_25777_, _25776_, _23832_);
  nor (_25778_, _25777_, _25773_);
  nor (_26894_[3], _25778_, rst);
  nor (_25779_, _24238_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_25780_, _25779_, _25566_);
  nor (_25781_, _25780_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_25782_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  not (_25783_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand (_25784_, _25781_, _25783_);
  and (_25785_, _25784_, _22761_);
  and (_26912_[0], _25785_, _25782_);
  or (_25786_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  not (_25787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_25788_, _25781_, _25787_);
  and (_25789_, _25788_, _22761_);
  and (_26912_[1], _25789_, _25786_);
  or (_25790_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  not (_25791_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_25792_, _25781_, _25791_);
  and (_25793_, _25792_, _22761_);
  and (_26912_[2], _25793_, _25790_);
  or (_25794_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not (_25795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand (_25796_, _25781_, _25795_);
  and (_25797_, _25796_, _22761_);
  and (_26912_[3], _25797_, _25794_);
  or (_25798_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not (_25799_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand (_25800_, _25781_, _25799_);
  and (_25801_, _25800_, _22761_);
  and (_26912_[4], _25801_, _25798_);
  or (_25802_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not (_25803_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_25804_, _25781_, _25803_);
  and (_25805_, _25804_, _22761_);
  and (_26912_[5], _25805_, _25802_);
  or (_25806_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  not (_25807_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_25808_, _25781_, _25807_);
  and (_25809_, _25808_, _22761_);
  and (_26912_[6], _25809_, _25806_);
  or (_25810_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  not (_25811_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand (_25812_, _25781_, _25811_);
  and (_25813_, _25812_, _22761_);
  and (_26912_[7], _25813_, _25810_);
  or (_25814_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not (_25815_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_25816_, _25781_, _25815_);
  and (_25818_, _25816_, _22761_);
  and (_26912_[8], _25818_, _25814_);
  or (_25819_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  not (_25820_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_25821_, _25781_, _25820_);
  and (_25822_, _25821_, _22761_);
  and (_26912_[9], _25822_, _25819_);
  or (_25823_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  not (_25824_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_25825_, _25781_, _25824_);
  and (_25826_, _25825_, _22761_);
  and (_26912_[10], _25826_, _25823_);
  or (_25827_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  not (_25828_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_25829_, _25781_, _25828_);
  and (_25830_, _25829_, _22761_);
  and (_26912_[11], _25830_, _25827_);
  or (_25832_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  not (_25833_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand (_25834_, _25781_, _25833_);
  and (_25835_, _25834_, _22761_);
  and (_26912_[12], _25835_, _25832_);
  or (_25836_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not (_25837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_25838_, _25781_, _25837_);
  and (_25839_, _25838_, _22761_);
  and (_26912_[13], _25839_, _25836_);
  or (_25840_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  not (_25841_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_25842_, _25781_, _25841_);
  and (_25843_, _25842_, _22761_);
  and (_26912_[14], _25843_, _25840_);
  and (_25844_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not (_25845_, _25781_);
  and (_25846_, _25845_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  or (_25847_, _25846_, _25844_);
  and (_26912_[15], _25847_, _22761_);
  or (_25848_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  not (_25849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_25850_, _25781_, _25849_);
  and (_25852_, _25850_, _22761_);
  and (_26912_[16], _25852_, _25848_);
  or (_25853_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not (_25855_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_25856_, _25781_, _25855_);
  and (_25857_, _25856_, _22761_);
  and (_26912_[17], _25857_, _25853_);
  or (_25858_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not (_25859_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_25860_, _25781_, _25859_);
  and (_25861_, _25860_, _22761_);
  and (_26912_[18], _25861_, _25858_);
  or (_25862_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not (_25863_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_25864_, _25781_, _25863_);
  and (_25865_, _25864_, _22761_);
  and (_26912_[19], _25865_, _25862_);
  or (_25866_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  not (_25867_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_25868_, _25781_, _25867_);
  and (_25869_, _25868_, _22761_);
  and (_26912_[20], _25869_, _25866_);
  or (_25870_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  not (_25871_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_25872_, _25781_, _25871_);
  and (_25873_, _25872_, _22761_);
  and (_26912_[21], _25873_, _25870_);
  or (_25874_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not (_25875_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_25876_, _25781_, _25875_);
  and (_25877_, _25876_, _22761_);
  and (_26912_[22], _25877_, _25874_);
  and (_25878_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_25879_, _25845_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or (_25880_, _25879_, _25878_);
  and (_26912_[23], _25880_, _22761_);
  or (_25881_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  not (_25882_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_25883_, _25781_, _25882_);
  and (_25885_, _25883_, _22761_);
  and (_26912_[24], _25885_, _25881_);
  or (_25887_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  not (_25888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_25889_, _25781_, _25888_);
  and (_25890_, _25889_, _22761_);
  and (_26912_[25], _25890_, _25887_);
  or (_25891_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not (_25892_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_25893_, _25781_, _25892_);
  and (_25895_, _25893_, _22761_);
  and (_26912_[26], _25895_, _25891_);
  and (_25896_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_25897_, _25845_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or (_25898_, _25897_, _25896_);
  and (_26912_[27], _25898_, _22761_);
  and (_25899_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_25900_, _25845_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or (_25901_, _25900_, _25899_);
  and (_26912_[28], _25901_, _22761_);
  or (_25902_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not (_25903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_25904_, _25781_, _25903_);
  and (_25905_, _25904_, _22761_);
  and (_26912_[29], _25905_, _25902_);
  or (_25906_, _25781_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not (_25907_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_25908_, _25781_, _25907_);
  and (_25909_, _25908_, _22761_);
  and (_26912_[30], _25909_, _25906_);
  nor (_25910_, _25611_, _23914_);
  and (_25911_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or (_21584_, _25911_, _25910_);
  and (_25913_, _25772_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_25914_, _25776_, _23914_);
  nor (_25915_, _25914_, _25913_);
  not (_25916_, _25915_);
  and (_25917_, _25778_, _24413_);
  and (_25918_, _25917_, _25916_);
  and (_25920_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_25921_, _25917_, _25915_);
  and (_25922_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_25923_, _25922_, _25920_);
  not (_25924_, _24413_);
  nor (_25925_, _25778_, _25924_);
  and (_25926_, _25925_, _25916_);
  and (_25927_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_25928_, _25778_, _25924_);
  and (_25929_, _25928_, _25916_);
  and (_25930_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_25932_, _25930_, _25927_);
  and (_25933_, _25932_, _25923_);
  nor (_25934_, _25915_, _22951_);
  and (_25935_, _25915_, _22951_);
  nor (_25936_, _25935_, _25934_);
  not (_25937_, _25936_);
  or (_25938_, _25778_, _22913_);
  nand (_25940_, _25778_, _22913_);
  nand (_25941_, _25940_, _25938_);
  and (_25942_, _24413_, _22926_);
  not (_25943_, _25942_);
  nor (_25945_, _24413_, _22926_);
  not (_25946_, _25523_);
  and (_25948_, _23874_, _23596_);
  and (_25949_, _25948_, _25215_);
  and (_25950_, _25948_, _25525_);
  nor (_25952_, _25950_, _25949_);
  and (_25953_, _24713_, _22914_);
  and (_25955_, _25948_, _25953_);
  not (_25956_, _25955_);
  and (_25958_, _25948_, _23887_);
  nor (_25959_, _25958_, _25608_);
  and (_25960_, _25959_, _25956_);
  and (_25961_, _25960_, _25952_);
  and (_25963_, _25526_, _23887_);
  and (_25964_, _25526_, _25953_);
  nor (_25965_, _25964_, _25528_);
  not (_25966_, _25965_);
  nor (_25967_, _25966_, _25963_);
  and (_25968_, _25967_, _25961_);
  or (_25970_, _25968_, _25946_);
  nor (_25971_, _25970_, _25945_);
  and (_25972_, _25971_, _25943_);
  and (_25974_, _25972_, _25941_);
  and (_25975_, _25974_, _25937_);
  not (_25976_, _25975_);
  and (_25977_, _25925_, _25915_);
  nand (_25978_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_25979_, _25778_, _24413_);
  and (_25980_, _25979_, _25915_);
  nand (_25981_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_25983_, _25981_, _25978_);
  and (_25984_, _25979_, _25916_);
  nand (_25985_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_25986_, _25928_, _25915_);
  nand (_25987_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_25988_, _25987_, _25985_);
  and (_25989_, _25988_, _25983_);
  and (_25990_, _25989_, _25976_);
  and (_25991_, _25990_, _25933_);
  and (_25993_, _25975_, _23669_);
  nor (_25994_, _25993_, _25991_);
  and (_26895_[0], _25994_, _22761_);
  and (_25995_, _25975_, _23784_);
  and (_25996_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_25997_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_25999_, _25997_, _25996_);
  and (_26000_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_26001_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_26002_, _26001_, _26000_);
  and (_26003_, _26002_, _25999_);
  and (_26004_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_26005_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_26006_, _26005_, _26004_);
  and (_26008_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_26010_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_26011_, _26010_, _26008_);
  and (_26013_, _26011_, _26006_);
  and (_26014_, _26013_, _25976_);
  and (_26015_, _26014_, _26003_);
  nor (_26016_, _26015_, _25995_);
  and (_26895_[1], _26016_, _22761_);
  and (_26017_, _25975_, _25268_);
  and (_26018_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_26019_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_26020_, _26019_, _26018_);
  and (_26021_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_26022_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_26023_, _26022_, _26021_);
  and (_26024_, _26023_, _26020_);
  and (_26025_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_26026_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_26027_, _26026_, _26025_);
  and (_26028_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_26029_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_26030_, _26029_, _26028_);
  and (_26032_, _26030_, _26027_);
  and (_26033_, _26032_, _25976_);
  and (_26034_, _26033_, _26024_);
  nor (_26035_, _26034_, _26017_);
  and (_26895_[2], _26035_, _22761_);
  and (_26036_, _25975_, _23832_);
  and (_26037_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_26038_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_26039_, _26038_, _26037_);
  and (_26040_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_26041_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_26042_, _26041_, _26040_);
  and (_26044_, _26042_, _26039_);
  nand (_26045_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nand (_26046_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_26047_, _26046_, _26045_);
  nand (_26048_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nand (_26049_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_26050_, _26049_, _26048_);
  and (_26051_, _26050_, _26047_);
  and (_26052_, _26051_, _25976_);
  and (_26053_, _26052_, _26044_);
  nor (_26054_, _26053_, _26036_);
  and (_26895_[3], _26054_, _22761_);
  and (_26055_, _25975_, _23914_);
  and (_26056_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_26057_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_26058_, _26057_, _26056_);
  and (_26059_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_26060_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_26061_, _26060_, _26059_);
  and (_26062_, _26061_, _26058_);
  and (_26063_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_26064_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_26065_, _26064_, _26063_);
  and (_26066_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_26067_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_26068_, _26067_, _26066_);
  and (_26069_, _26068_, _26065_);
  and (_26070_, _26069_, _25976_);
  and (_26071_, _26070_, _26062_);
  nor (_26072_, _26071_, _26055_);
  and (_26895_[4], _26072_, _22761_);
  and (_26073_, _25975_, _23628_);
  and (_26074_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_26075_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_26076_, _26075_, _26074_);
  and (_26077_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_26078_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_26079_, _26078_, _26077_);
  and (_26080_, _26079_, _26076_);
  and (_26081_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_26082_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor (_26083_, _26082_, _26081_);
  and (_26084_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_26085_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_26086_, _26085_, _26084_);
  and (_26087_, _26086_, _26083_);
  and (_26088_, _26087_, _25976_);
  and (_26089_, _26088_, _26080_);
  nor (_26090_, _26089_, _26073_);
  and (_26895_[5], _26090_, _22761_);
  and (_26091_, _25975_, _23748_);
  and (_26092_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_26093_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_26094_, _26093_, _26092_);
  and (_26095_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_26096_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_26097_, _26096_, _26095_);
  and (_26098_, _26097_, _26094_);
  and (_26099_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_26100_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_26101_, _26100_, _26099_);
  and (_26102_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_26103_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_26104_, _26103_, _26102_);
  and (_26105_, _26104_, _26101_);
  and (_26106_, _26105_, _25976_);
  and (_26107_, _26106_, _26098_);
  nor (_26108_, _26107_, _26091_);
  and (_26895_[6], _26108_, _22761_);
  nor (_26109_, _25611_, _23832_);
  and (_26110_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or (_21895_, _26110_, _26109_);
  and (_26111_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_26112_, _25619_, _23838_);
  or (_21926_, _26112_, _26111_);
  and (_26113_, _25400_, _23982_);
  and (_26114_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_21947_, _26114_, _26113_);
  and (_26115_, _25609_, _23718_);
  and (_26116_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or (_21968_, _26116_, _26115_);
  and (_26117_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_26118_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_26119_, _22770_, _26118_);
  or (_26120_, _26119_, _26117_);
  and (_26891_[6], _26120_, _22761_);
  and (_26121_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_26122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_26123_, _22770_, _26122_);
  or (_26124_, _26123_, _26121_);
  and (_26891_[5], _26124_, _22761_);
  and (_26125_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_26126_, _22770_, _22807_);
  or (_26127_, _26126_, _26125_);
  and (_26891_[4], _26127_, _22761_);
  and (_26128_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_26129_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26130_, _22770_, _26129_);
  or (_26131_, _26130_, _26128_);
  and (_26891_[3], _26131_, _22761_);
  and (_26132_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_26133_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_26134_, _22770_, _26133_);
  or (_26135_, _26134_, _26132_);
  and (_26891_[2], _26135_, _22761_);
  and (_26136_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_26137_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_26138_, _22770_, _26137_);
  or (_26139_, _26138_, _26136_);
  and (_26891_[1], _26139_, _22761_);
  and (_26140_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_26141_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26142_, _22770_, _26141_);
  or (_26143_, _26142_, _26140_);
  and (_26891_[0], _26143_, _22761_);
  nor (_26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_26145_, _26144_, _23271_);
  nor (_26146_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_26147_, _26146_, _26145_);
  and (_26148_, _23419_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_26149_, _26148_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_26150_, _26149_);
  and (_26151_, _23373_, _23090_);
  nor (_26152_, _26151_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26153_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_26154_, _23445_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26155_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26156_, _23121_, _26155_);
  nand (_26157_, _26156_, _26154_);
  or (_26158_, _23406_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26159_, _23372_, _26155_);
  nand (_26160_, _26159_, _26158_);
  and (_26161_, _26160_, _26157_);
  or (_26163_, _23217_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26164_, _23406_, _26155_);
  nand (_26165_, _26164_, _26163_);
  or (_26166_, _23121_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26167_, _23090_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26168_, _26167_, _26166_);
  and (_26169_, _26168_, _26165_);
  nand (_26170_, _26169_, _26161_);
  and (_26171_, _26170_, _26153_);
  nor (_26172_, _26171_, _26152_);
  or (_26173_, _23248_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26174_, _23445_, _26155_);
  nand (_26175_, _26174_, _26173_);
  and (_26176_, _26175_, _26153_);
  and (_26177_, _26168_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_26178_, _26177_, _26176_);
  not (_26179_, _26178_);
  nand (_26180_, _26144_, _23078_);
  nor (_26181_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_26182_, _26181_);
  and (_26183_, _26182_, _26180_);
  not (_26184_, _26183_);
  or (_26185_, _23419_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26186_, _23217_, _26155_);
  and (_26187_, _26186_, _26185_);
  or (_26188_, _26187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26189_, _26160_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26190_, _26189_, _26188_);
  or (_26191_, _26190_, _26184_);
  and (_26192_, _23248_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26193_, _26192_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26194_, _26157_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26195_, _26194_, _26193_);
  nand (_26196_, _26144_, _23366_);
  nor (_26197_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_26198_, _26197_);
  and (_26199_, _26198_, _26196_);
  not (_26200_, _26199_);
  or (_26201_, _26200_, _26195_);
  nand (_26202_, _26189_, _26188_);
  or (_26203_, _26202_, _26183_);
  and (_26204_, _26203_, _26191_);
  not (_26205_, _26204_);
  or (_26206_, _26205_, _26201_);
  and (_26207_, _26206_, _26191_);
  nand (_26208_, _26194_, _26193_);
  or (_26209_, _26199_, _26208_);
  and (_26210_, _26209_, _26201_);
  and (_26211_, _26210_, _26204_);
  not (_26212_, _26144_);
  or (_26213_, _26212_, _23115_);
  nor (_26214_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_26215_, _26214_);
  nand (_26216_, _26215_, _26213_);
  or (_26217_, _26148_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26218_, _26165_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26219_, _26218_, _26217_);
  or (_26220_, _26219_, _26216_);
  nor (_26221_, _26175_, _26153_);
  nor (_26222_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_26224_, _26222_);
  nand (_26225_, _26144_, _23146_);
  and (_26226_, _26225_, _26224_);
  not (_26227_, _26226_);
  or (_26228_, _26227_, _26221_);
  and (_26229_, _26215_, _26213_);
  nand (_26230_, _26218_, _26217_);
  or (_26231_, _26230_, _26229_);
  nand (_26232_, _26231_, _26220_);
  or (_26233_, _26232_, _26228_);
  nand (_26234_, _26233_, _26220_);
  nand (_26235_, _26234_, _26211_);
  and (_26236_, _26235_, _26207_);
  and (_26237_, _26187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_26238_, _26237_);
  nand (_26239_, _26144_, _23178_);
  nor (_26240_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_26241_, _26240_);
  and (_26242_, _26241_, _26239_);
  nand (_26243_, _26242_, _26238_);
  or (_26244_, _26242_, _26238_);
  nand (_26245_, _26244_, _26243_);
  nand (_26246_, _26192_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_26247_, _26212_, _23211_);
  nor (_26248_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_26249_, _26248_);
  and (_26250_, _26249_, _26247_);
  nand (_26251_, _26250_, _26246_);
  or (_26252_, _26212_, _23242_);
  nor (_26253_, _26144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_26254_, _26253_);
  nand (_26255_, _26254_, _26252_);
  and (_26256_, _26255_, _26149_);
  or (_26257_, _26250_, _26246_);
  nand (_26258_, _26257_, _26251_);
  or (_26259_, _26258_, _26256_);
  and (_26260_, _26259_, _26251_);
  or (_26261_, _26260_, _26245_);
  nand (_26262_, _26261_, _26243_);
  not (_26263_, _26221_);
  or (_26264_, _26226_, _26263_);
  and (_26265_, _26264_, _26228_);
  and (_26266_, _26231_, _26220_);
  and (_26267_, _26266_, _26265_);
  and (_26268_, _26267_, _26211_);
  nand (_26269_, _26268_, _26262_);
  nand (_26270_, _26269_, _26236_);
  and (_26271_, _26179_, _26172_);
  and (_26272_, _26271_, _26270_);
  nor (_26273_, _26272_, _26183_);
  not (_26274_, _26273_);
  and (_26275_, _26219_, _26216_);
  and (_26276_, _26265_, _26262_);
  not (_26277_, _26276_);
  and (_26278_, _26277_, _26228_);
  or (_26279_, _26278_, _26275_);
  and (_26280_, _26279_, _26220_);
  not (_26281_, _26280_);
  nand (_26282_, _26281_, _26210_);
  nand (_26283_, _26282_, _26201_);
  nand (_26284_, _26283_, _26205_);
  nand (_26285_, _26284_, _26272_);
  and (_26286_, _26285_, _26274_);
  and (_26287_, _26286_, _26179_);
  not (_26288_, _26287_);
  nor (_26289_, _26286_, _26179_);
  or (_26290_, _26281_, _26210_);
  nand (_26291_, _26290_, _26282_);
  nand (_26292_, _26291_, _26272_);
  nor (_26293_, _26272_, _26199_);
  not (_26294_, _26293_);
  nand (_26295_, _26294_, _26292_);
  or (_26296_, _26295_, _26190_);
  or (_26297_, _26296_, _26289_);
  nand (_26298_, _26297_, _26288_);
  or (_26299_, _26289_, _26287_);
  nand (_26300_, _26295_, _26190_);
  nand (_26301_, _26300_, _26296_);
  nor (_26302_, _26301_, _26299_);
  nand (_26303_, _26232_, _26278_);
  or (_26304_, _26232_, _26278_);
  nand (_26305_, _26304_, _26303_);
  nand (_26306_, _26305_, _26272_);
  nor (_26307_, _26272_, _26229_);
  not (_26308_, _26307_);
  and (_26309_, _26308_, _26306_);
  and (_26310_, _26309_, _26208_);
  not (_26311_, _26310_);
  nor (_26312_, _26272_, _26227_);
  nor (_26313_, _26265_, _26262_);
  nor (_26314_, _26313_, _26276_);
  and (_26315_, _26314_, _26272_);
  or (_26316_, _26315_, _26312_);
  and (_26317_, _26316_, _26230_);
  not (_26318_, _26317_);
  nor (_26319_, _26309_, _26208_);
  or (_26320_, _26319_, _26310_);
  or (_26321_, _26320_, _26318_);
  nand (_26322_, _26321_, _26311_);
  not (_26323_, _26272_);
  and (_26324_, _26260_, _26245_);
  not (_26325_, _26324_);
  and (_26326_, _26325_, _26261_);
  or (_26327_, _26326_, _26323_);
  or (_26328_, _26272_, _26242_);
  and (_26329_, _26328_, _26327_);
  nor (_26330_, _26329_, _26263_);
  not (_26331_, _26330_);
  or (_26332_, _26272_, _26255_);
  and (_26333_, _26255_, _26150_);
  nor (_26334_, _26255_, _26150_);
  nor (_26335_, _26334_, _26333_);
  nand (_26336_, _26272_, _26335_);
  nand (_26337_, _26336_, _26332_);
  nand (_26338_, _26337_, _26246_);
  or (_26339_, _26337_, _26246_);
  nand (_26340_, _26339_, _26338_);
  nor (_26341_, _26150_, _26147_);
  or (_26342_, _26341_, _26340_);
  and (_26343_, _26342_, _26338_);
  and (_26344_, _26258_, _26256_);
  not (_26345_, _26344_);
  and (_26346_, _26345_, _26259_);
  or (_26347_, _26346_, _26323_);
  or (_26348_, _26272_, _26250_);
  and (_26349_, _26348_, _26347_);
  nand (_26350_, _26349_, _26238_);
  or (_26351_, _26349_, _26238_);
  nand (_26352_, _26351_, _26350_);
  or (_26353_, _26352_, _26343_);
  and (_26354_, _26329_, _26263_);
  not (_26355_, _26354_);
  and (_26356_, _26355_, _26350_);
  nand (_26357_, _26356_, _26353_);
  nand (_26358_, _26357_, _26331_);
  not (_26359_, _26358_);
  nor (_26360_, _26316_, _26230_);
  nor (_26361_, _26360_, _26317_);
  not (_26362_, _26361_);
  nor (_26363_, _26320_, _26362_);
  and (_26364_, _26363_, _26359_);
  or (_26365_, _26364_, _26322_);
  and (_26366_, _26365_, _26302_);
  or (_26367_, _26366_, _26298_);
  nand (_26368_, _26367_, _26172_);
  or (_26369_, _26368_, _26150_);
  and (_26370_, _26369_, _26147_);
  nor (_26371_, _26369_, _26147_);
  or (_26372_, _26371_, _26370_);
  nand (_26373_, _26372_, _23528_);
  nor (_26375_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_26376_, _26375_);
  and (_26377_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  not (_26378_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_26379_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _26378_);
  not (_26380_, _26379_);
  or (_26381_, _26380_, _23184_);
  not (_26382_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_26383_, _26382_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_26384_, _26383_);
  or (_26385_, _26384_, _23404_);
  and (_26386_, _26385_, _26381_);
  or (_26387_, _26383_, _26379_);
  or (_26388_, _26387_, _23423_);
  and (_26389_, _26388_, _26376_);
  nand (_26390_, _26389_, _26386_);
  nand (_26391_, _26375_, _23090_);
  and (_26392_, _26391_, _26390_);
  and (_26393_, _26392_, _23242_);
  or (_26394_, _26380_, _23427_);
  or (_26395_, _26384_, _23152_);
  and (_26396_, _26395_, _26394_);
  or (_26397_, _26387_, _23278_);
  and (_26398_, _26397_, _26376_);
  nand (_26399_, _26398_, _26396_);
  or (_26400_, _26376_, _23372_);
  and (_26401_, _26400_, _26399_);
  and (_26402_, _26401_, _23211_);
  nand (_26403_, _26402_, _26393_);
  and (_26404_, _26401_, _23552_);
  nand (_26405_, _26400_, _26399_);
  or (_26406_, _26405_, _23777_);
  and (_26407_, _26392_, _23211_);
  and (_26408_, _26407_, _26406_);
  nand (_26409_, _26408_, _26404_);
  nand (_26410_, _26409_, _26403_);
  nand (_26411_, _26391_, _26390_);
  or (_26412_, _26411_, _23178_);
  or (_26413_, _26405_, _23146_);
  or (_26414_, _26413_, _26412_);
  nand (_26415_, _26413_, _26412_);
  and (_26416_, _26415_, _26414_);
  and (_26417_, _26416_, _26410_);
  and (_26418_, _26392_, _23551_);
  and (_26419_, _26418_, _26404_);
  or (_26420_, _26411_, _23469_);
  or (_26421_, _26420_, _26413_);
  and (_26422_, _26401_, _23115_);
  or (_26423_, _26422_, _26418_);
  and (_26424_, _26423_, _26421_);
  nand (_26426_, _26424_, _26419_);
  or (_26427_, _26424_, _26419_);
  and (_26428_, _26427_, _26426_);
  nand (_26429_, _26428_, _26417_);
  not (_26430_, _26420_);
  or (_26431_, _26421_, _23366_);
  and (_26432_, _26401_, _23550_);
  not (_26433_, _26432_);
  nand (_26434_, _26433_, _26421_);
  and (_26435_, _26434_, _26431_);
  nand (_26436_, _26435_, _26430_);
  or (_26437_, _26432_, _26430_);
  nand (_26438_, _26437_, _26436_);
  or (_26439_, _26438_, _26429_);
  or (_26440_, _26411_, _23271_);
  nor (_26441_, _26440_, _26406_);
  or (_26442_, _26402_, _26393_);
  and (_26443_, _26442_, _26403_);
  and (_26444_, _26443_, _26441_);
  or (_26445_, _26408_, _26404_);
  and (_26446_, _26445_, _26409_);
  and (_26447_, _26446_, _26444_);
  nand (_26448_, _26416_, _26410_);
  or (_26449_, _26416_, _26410_);
  and (_26450_, _26449_, _26448_);
  and (_26451_, _26450_, _26447_);
  or (_26452_, _26428_, _26417_);
  and (_26453_, _26452_, _26429_);
  nand (_26454_, _26453_, _26451_);
  not (_26455_, _26454_);
  and (_26456_, _26429_, _26426_);
  nand (_26457_, _26456_, _26438_);
  or (_26458_, _26456_, _26438_);
  and (_26459_, _26458_, _26457_);
  nand (_26460_, _26459_, _26455_);
  nand (_26461_, _26460_, _26439_);
  nor (_26462_, _26438_, _26426_);
  not (_26463_, _26431_);
  and (_26464_, _26435_, _26430_);
  or (_26465_, _26405_, _23078_);
  or (_26466_, _26411_, _23366_);
  or (_26467_, _26466_, _26465_);
  nand (_26468_, _26466_, _26465_);
  and (_26469_, _26468_, _26467_);
  nand (_26470_, _26469_, _26464_);
  or (_26471_, _26469_, _26464_);
  and (_26472_, _26471_, _26470_);
  nand (_26473_, _26472_, _26463_);
  or (_26474_, _26472_, _26463_);
  and (_26475_, _26474_, _26473_);
  nand (_26476_, _26475_, _26462_);
  or (_26477_, _26475_, _26462_);
  and (_26478_, _26477_, _26476_);
  nand (_26479_, _26478_, _26461_);
  or (_26480_, _26478_, _26461_);
  and (_26481_, _26480_, _26479_);
  nand (_26482_, _26481_, _26377_);
  or (_26483_, _26481_, _26377_);
  and (_26484_, _26483_, _26482_);
  and (_26485_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_26486_, _26459_, _26455_);
  and (_26487_, _26486_, _26460_);
  nand (_26488_, _26487_, _26485_);
  or (_26489_, _26487_, _26485_);
  nand (_26490_, _26489_, _26488_);
  and (_26491_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or (_26492_, _26453_, _26451_);
  and (_26493_, _26492_, _26454_);
  nand (_26494_, _26493_, _26491_);
  or (_26495_, _26493_, _26491_);
  and (_26496_, _26495_, _26494_);
  and (_26497_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nand (_26498_, _26450_, _26447_);
  or (_26499_, _26450_, _26447_);
  and (_26500_, _26499_, _26498_);
  nand (_26501_, _26500_, _26497_);
  and (_26502_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nand (_26503_, _26446_, _26444_);
  or (_26504_, _26446_, _26444_);
  and (_26505_, _26504_, _26503_);
  nand (_26506_, _26505_, _26502_);
  and (_26507_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_26508_, _26443_, _26441_);
  or (_26509_, _26443_, _26441_);
  and (_26510_, _26509_, _26508_);
  and (_26511_, _26510_, _26507_);
  not (_26512_, _26511_);
  or (_26513_, _26505_, _26502_);
  nand (_26514_, _26513_, _26506_);
  or (_26515_, _26514_, _26512_);
  nand (_26516_, _26515_, _26506_);
  or (_26517_, _26500_, _26497_);
  and (_26518_, _26517_, _26501_);
  nand (_26519_, _26518_, _26516_);
  nand (_26520_, _26519_, _26501_);
  nand (_26521_, _26520_, _26496_);
  and (_26522_, _26521_, _26494_);
  or (_26523_, _26522_, _26490_);
  nand (_26524_, _26523_, _26488_);
  nand (_26526_, _26524_, _26484_);
  nand (_26528_, _26526_, _26482_);
  and (_26529_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  nand (_26530_, _26479_, _26476_);
  and (_26531_, _26392_, _23508_);
  and (_26532_, _26531_, _26433_);
  and (_26533_, _26473_, _26470_);
  not (_26534_, _26533_);
  nand (_26535_, _26534_, _26532_);
  or (_26536_, _26534_, _26532_);
  and (_26537_, _26536_, _26535_);
  nand (_26538_, _26537_, _26530_);
  or (_26539_, _26537_, _26530_);
  and (_26540_, _26539_, _26538_);
  nand (_26541_, _26540_, _26529_);
  or (_26542_, _26540_, _26529_);
  and (_26543_, _26542_, _26541_);
  and (_26544_, _26543_, _26528_);
  nor (_26545_, _26543_, _26528_);
  nor (_26546_, _26545_, _26544_);
  and (_26547_, _26546_, _23531_);
  and (_26548_, _23509_, _23330_);
  or (_26549_, _23462_, _23271_);
  nand (_26550_, _23534_, _23242_);
  and (_26551_, _23487_, _23508_);
  not (_26552_, _23494_);
  nor (_26553_, _26552_, _23271_);
  nor (_26554_, _26553_, _26551_);
  and (_26555_, _26554_, _26550_);
  and (_26556_, _26555_, _26549_);
  nand (_26557_, _26556_, _23663_);
  nor (_26558_, _26557_, _26548_);
  and (_26559_, _23439_, _23468_);
  nor (_26560_, _26559_, _23334_);
  nor (_26561_, _23398_, _23037_);
  not (_26562_, _26561_);
  and (_26563_, _26562_, _26560_);
  nor (_26564_, _26563_, _23667_);
  and (_26565_, _26564_, _26558_);
  not (_26566_, _26565_);
  nor (_26567_, _26566_, _26547_);
  nand (_26568_, _26567_, _26373_);
  not (_26569_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_26570_, \oc8051_top_1.oc8051_decoder1.state [1], _22765_);
  and (_26571_, _26570_, _26569_);
  and (_26572_, _24487_, _24418_);
  and (_26574_, _26572_, _26571_);
  or (_26575_, _22767_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26576_, _26575_);
  and (_26577_, _24416_, _25924_);
  and (_26578_, _26577_, _24515_);
  and (_26579_, _24413_, _24269_);
  and (_26580_, _24495_, _26579_);
  nor (_26581_, _26580_, _26578_);
  nor (_26582_, _26581_, _26576_);
  nor (_26583_, _26582_, _26574_);
  and (_26584_, _24515_, _24443_);
  and (_26585_, _24496_, _26584_);
  not (_26587_, _24391_);
  nor (_26588_, _24443_, _26587_);
  and (_26589_, _24496_, _26588_);
  or (_26590_, _26589_, _26585_);
  and (_26591_, _24443_, _24391_);
  and (_26592_, _24496_, _26591_);
  nor (_26593_, _26592_, _26590_);
  and (_26594_, _24517_, _24489_);
  and (_26595_, _24447_, _24443_);
  and (_26596_, _26595_, _24321_);
  or (_26597_, _26596_, _26594_);
  and (_26598_, _26595_, _24466_);
  and (_26599_, _24458_, _24447_);
  or (_26600_, _26599_, _26598_);
  nor (_26601_, _26600_, _26597_);
  nand (_26602_, _26601_, _26593_);
  nand (_26603_, _26602_, _26571_);
  and (_26604_, _26578_, _26575_);
  not (_26605_, _26604_);
  and (_26606_, _24527_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_26607_, _26577_, _24391_);
  and (_26608_, _26607_, _26606_);
  and (_26609_, _24496_, _24391_);
  and (_26610_, _26609_, _26575_);
  nor (_26611_, _26610_, _26608_);
  and (_26612_, _26611_, _26605_);
  and (_26614_, _26612_, _26603_);
  not (_26615_, _26614_);
  not (_26616_, _26593_);
  and (_26617_, _24516_, _24458_);
  nor (_26618_, _26617_, _26597_);
  and (_26619_, _24496_, _24451_);
  not (_26620_, _26619_);
  and (_26621_, _24470_, _24445_);
  and (_26622_, _26621_, _24496_);
  nor (_26623_, _26622_, _26572_);
  nand (_26624_, _26623_, _26620_);
  nor (_26625_, _26624_, _26600_);
  nand (_26626_, _26625_, _26618_);
  or (_26627_, _26626_, _26616_);
  and (_26628_, _26627_, _26571_);
  nor (_26629_, _26628_, _26615_);
  and (_26630_, _26629_, _26583_);
  or (_26631_, _26630_, _26574_);
  and (_26632_, _26631_, _26568_);
  and (_26633_, _26619_, _26571_);
  not (_26634_, _26633_);
  nor (_26635_, _26609_, _26585_);
  and (_26636_, _26633_, _24459_);
  not (_26637_, _26636_);
  and (_26638_, _26637_, _26635_);
  nor (_26639_, _26638_, _24527_);
  and (_26640_, _26639_, _26634_);
  and (_26641_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26642_, _26641_);
  and (_26643_, _24496_, _24460_);
  and (_26644_, _26643_, _26571_);
  nor (_26645_, _26644_, _26616_);
  nor (_26646_, _26645_, _24527_);
  nor (_26647_, _26646_, _26634_);
  nor (_26648_, _24506_, _24473_);
  and (_26650_, _24468_, _24470_);
  not (_26651_, _24466_);
  nor (_26652_, _24479_, _24391_);
  nor (_26653_, _26652_, _26651_);
  nor (_26654_, _26653_, _26650_);
  and (_26655_, _26654_, _26648_);
  and (_26656_, _24466_, _24443_);
  and (_26657_, _26656_, _24447_);
  and (_26658_, _24466_, _24515_);
  nor (_26659_, _26658_, _26657_);
  not (_26660_, _24449_);
  and (_26661_, _24471_, _24418_);
  nor (_26662_, _26572_, _26661_);
  and (_26663_, _26662_, _26660_);
  and (_26664_, _24516_, _24466_);
  and (_26665_, _24517_, _24496_);
  or (_26666_, _26665_, _26607_);
  nor (_26667_, _26666_, _26664_);
  and (_26668_, _26667_, _26663_);
  and (_26670_, _26668_, _26659_);
  and (_26671_, _26670_, _26655_);
  nor (_26672_, _26671_, _26576_);
  or (_26673_, _26672_, _26608_);
  or (_26674_, _26673_, _26647_);
  nand (_26675_, _26674_, _22765_);
  and (_26676_, _26675_, _26642_);
  and (_26677_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26679_, _26677_);
  and (_26680_, _24496_, _24448_);
  and (_26681_, _26577_, _24487_);
  nor (_26682_, _26681_, _26680_);
  and (_26683_, _24499_, _24418_);
  and (_26685_, _26577_, _24499_);
  nor (_26686_, _26685_, _26683_);
  and (_26687_, _26686_, _26682_);
  and (_26688_, _24499_, _24489_);
  and (_26689_, _26584_, _24489_);
  nor (_26690_, _26689_, _26688_);
  and (_26691_, _26690_, _26687_);
  and (_26692_, _24516_, _24445_);
  and (_26693_, _26692_, _26577_);
  and (_26694_, _26595_, _24416_);
  and (_26695_, _26694_, _25924_);
  nor (_26696_, _26695_, _26693_);
  and (_26697_, _26595_, _24496_);
  nor (_26698_, _26697_, _26594_);
  and (_26699_, _26698_, _26696_);
  and (_26700_, _26699_, _26691_);
  not (_26701_, _24493_);
  and (_26702_, _26635_, _26701_);
  and (_26703_, _24453_, _24489_);
  not (_26705_, _26703_);
  nand (_26706_, _24453_, _24418_);
  nand (_26707_, _26577_, _24453_);
  and (_26708_, _26707_, _26706_);
  and (_26709_, _26708_, _26705_);
  and (_26710_, _26709_, _26702_);
  and (_26711_, _26692_, _24489_);
  not (_26712_, _26577_);
  nor (_26713_, _24517_, _24471_);
  nor (_26714_, _26713_, _26712_);
  nor (_26715_, _26714_, _26711_);
  and (_26716_, _24516_, _24496_);
  nor (_26717_, _26716_, _26607_);
  and (_26718_, _24474_, _24447_);
  nand (_26719_, _26577_, _24448_);
  not (_26720_, _26719_);
  nor (_26721_, _26720_, _26718_);
  and (_26722_, _26721_, _26717_);
  and (_26723_, _26722_, _26715_);
  and (_26724_, _26723_, _26710_);
  and (_26725_, _24471_, _24489_);
  and (_26726_, _26595_, _24489_);
  and (_26727_, _26577_, _26621_);
  and (_26728_, _24479_, _24416_);
  or (_26729_, _26728_, _26727_);
  or (_26730_, _26729_, _26726_);
  nor (_26731_, _26730_, _26725_);
  and (_26732_, _26621_, _24489_);
  not (_26733_, _24489_);
  nor (_26735_, _26652_, _26733_);
  nor (_26736_, _26735_, _26732_);
  and (_26737_, _24515_, _24445_);
  and (_26739_, _26737_, _24489_);
  and (_26740_, _24466_, _24448_);
  nor (_26741_, _26740_, _26739_);
  and (_26742_, _26741_, _26736_);
  and (_26743_, _26742_, _26731_);
  and (_26744_, _26743_, _26724_);
  nand (_26745_, _26744_, _26700_);
  nand (_26746_, _26745_, _26575_);
  nor (_26747_, _26633_, _26608_);
  nand (_26748_, _26747_, _26746_);
  nand (_26749_, _26748_, _22765_);
  and (_26750_, _26749_, _26679_);
  nor (_26751_, _26750_, _26676_);
  and (_26752_, _25525_, _23888_);
  and (_26753_, _26752_, _23585_);
  and (_26754_, _26752_, _23709_);
  not (_26755_, _26752_);
  and (_26756_, _26755_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or (_26757_, _26756_, _26754_);
  nor (_26758_, _26755_, _23784_);
  and (_26759_, _26755_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_26760_, _26759_, _26758_);
  or (_26761_, _26752_, _22921_);
  nand (_26762_, _26752_, _24763_);
  and (_26764_, _26762_, _26761_);
  and (_26765_, _26764_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_26766_, _26765_, _26760_);
  not (_26767_, _26766_);
  nor (_26768_, _26767_, _26757_);
  nor (_26769_, _26755_, _23832_);
  and (_26770_, _26755_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_26771_, _26770_, _26769_);
  nand (_26772_, _26771_, _26768_);
  nor (_26773_, _26755_, _23914_);
  and (_26774_, _26755_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_26775_, _26774_, _26773_);
  not (_26776_, _26775_);
  nor (_26777_, _26776_, _26772_);
  nor (_26778_, _26755_, _23628_);
  and (_26779_, _26755_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_26780_, _26779_, _26778_);
  and (_26781_, _26780_, _26777_);
  nor (_26782_, _26755_, _23748_);
  and (_26783_, _26755_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_26784_, _26783_, _26782_);
  and (_26785_, _26784_, _26781_);
  and (_26786_, _26755_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or (_26787_, _26786_, _26785_);
  nand (_26788_, _26786_, _26785_);
  and (_26789_, _26788_, _26787_);
  nand (_26790_, _26789_, _22893_);
  nor (_26791_, _26752_, _22871_);
  and (_26792_, _26791_, _26790_);
  nor (_26794_, _26792_, _26753_);
  nand (_26795_, _26794_, _26751_);
  not (_26796_, _26676_);
  and (_26797_, _26750_, _26796_);
  nand (_26798_, _25918_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand (_26799_, _25980_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_26800_, _26799_, _26798_);
  nand (_26801_, _25977_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand (_26802_, _25986_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_26803_, _26802_, _26801_);
  and (_26804_, _26803_, _26800_);
  nand (_26805_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand (_26806_, _25929_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_26807_, _26806_, _26805_);
  nand (_26809_, _25984_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand (_26810_, _25921_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_26811_, _26810_, _26809_);
  and (_26812_, _26811_, _26807_);
  and (_26813_, _26812_, _25976_);
  and (_26814_, _26813_, _26804_);
  and (_26815_, _25975_, _23585_);
  nor (_26816_, _26815_, _26814_);
  nand (_26817_, _26816_, _26797_);
  and (_26818_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_26819_, _24448_, _24486_);
  and (_26820_, _26819_, _22765_);
  and (_26821_, _26621_, _24486_);
  and (_26822_, _26821_, _22765_);
  nor (_26823_, _26822_, _26820_);
  nor (_26824_, _26823_, _22767_);
  not (_26825_, _26824_);
  nor (_26826_, _26821_, _26819_);
  and (_26827_, _26663_, _26826_);
  nor (_26828_, _26827_, _26576_);
  nor (_26829_, _26828_, _26633_);
  and (_26830_, _26829_, _26825_);
  nor (_26831_, _26830_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_26832_, _26831_, _26818_);
  not (_26833_, _25739_);
  nor (_26834_, _26750_, _26796_);
  nand (_26835_, _26834_, _26833_);
  and (_26836_, _26835_, _26832_);
  and (_26837_, _26836_, _26817_);
  nand (_26838_, _26837_, _26795_);
  and (_26839_, _26838_, _22890_);
  nor (_26840_, _26838_, _22890_);
  nor (_26841_, _26840_, _26839_);
  and (_26842_, _26751_, _26832_);
  not (_26843_, _26842_);
  or (_26844_, _26776_, _26772_);
  not (_26845_, _26780_);
  and (_26846_, _26845_, _26844_);
  nor (_26847_, _26846_, _26781_);
  nor (_26848_, _26847_, _22861_);
  nor (_26849_, _26848_, _22990_);
  nor (_26850_, _26849_, _26752_);
  nor (_00001_, _26850_, _26778_);
  nor (_00002_, _00001_, _26843_);
  not (_00003_, _00002_);
  and (_00004_, _26797_, _26832_);
  and (_00005_, _00004_, _26090_);
  not (_00006_, _00005_);
  and (_00007_, _26834_, _26832_);
  nor (_00008_, _22768_, _23099_);
  and (_00009_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00010_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_00011_, _00010_, _00009_);
  and (_00012_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00013_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_00014_, _00013_, _00012_);
  and (_00015_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_00016_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_00017_, _00016_, _00015_);
  and (_00018_, _00017_, _00014_);
  and (_00019_, _00018_, _00011_);
  nor (_00020_, _00019_, _25562_);
  nor (_00021_, _00020_, _00008_);
  not (_00022_, _00021_);
  and (_00023_, _00022_, _00007_);
  not (_00024_, _26797_);
  nor (_00025_, _26834_, _26832_);
  and (_00026_, _00025_, _00024_);
  nor (_00027_, _00026_, _00023_);
  and (_00028_, _00027_, _00006_);
  and (_00029_, _00028_, _00003_);
  nor (_00030_, _00029_, _22998_);
  and (_00031_, _00029_, _22998_);
  nor (_00032_, _00031_, _00030_);
  nor (_00033_, _00032_, _26841_);
  or (_00034_, _26845_, _26844_);
  not (_00035_, _26784_);
  and (_00036_, _00035_, _00034_);
  nor (_00037_, _00036_, _26785_);
  nor (_00038_, _00037_, _22861_);
  nor (_00039_, _00038_, _22973_);
  nor (_00040_, _00039_, _26752_);
  nor (_00041_, _00040_, _26782_);
  nor (_00042_, _00041_, _26843_);
  not (_00043_, _26832_);
  and (_00044_, _26797_, _00043_);
  and (_00045_, _26797_, _26108_);
  nor (_00046_, _22768_, _23352_);
  and (_00047_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00048_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_00050_, _00048_, _00047_);
  and (_00052_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00053_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_00054_, _00053_, _00052_);
  and (_00055_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_00056_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_00057_, _00056_, _00055_);
  and (_00058_, _00057_, _00054_);
  and (_00059_, _00058_, _00050_);
  nor (_00060_, _00059_, _25562_);
  nor (_00061_, _00060_, _00046_);
  not (_00062_, _00061_);
  and (_00063_, _00062_, _26834_);
  nor (_00064_, _00063_, _00045_);
  and (_00065_, _00064_, _26832_);
  nor (_00066_, _00065_, _00044_);
  nor (_00067_, _00066_, _00042_);
  nor (_00068_, _00067_, _22981_);
  and (_00069_, _00067_, _22981_);
  nor (_00070_, _00069_, _00068_);
  not (_00072_, _00070_);
  nand (_00073_, _00004_, _26054_);
  nor (_00074_, _22768_, _23161_);
  and (_00075_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00076_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_00078_, _00076_, _00075_);
  and (_00080_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00081_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_00082_, _00081_, _00080_);
  and (_00083_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00084_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_00086_, _00084_, _00083_);
  and (_00087_, _00086_, _00082_);
  and (_00088_, _00087_, _00078_);
  nor (_00089_, _00088_, _25562_);
  nor (_00090_, _00089_, _00074_);
  not (_00091_, _00090_);
  nand (_00092_, _00091_, _00007_);
  and (_00093_, _00092_, _00073_);
  or (_00094_, _26771_, _26768_);
  nand (_00095_, _00094_, _26772_);
  nand (_00096_, _00095_, _22893_);
  nand (_00097_, _00096_, _22899_);
  and (_00098_, _00097_, _26755_);
  or (_00099_, _00098_, _26769_);
  nand (_00100_, _00099_, _26842_);
  and (_00101_, _26750_, _26676_);
  and (_00102_, _00101_, _26832_);
  not (_00103_, _00102_);
  or (_00104_, _00103_, _25778_);
  and (_00105_, _00104_, _00100_);
  and (_00106_, _00105_, _00093_);
  nor (_00108_, _00106_, _22913_);
  and (_00109_, _00106_, _22913_);
  nor (_00110_, _00109_, _00108_);
  and (_00111_, _26776_, _26772_);
  nor (_00112_, _00111_, _26777_);
  nor (_00113_, _00112_, _22861_);
  nor (_00114_, _00113_, _22940_);
  nor (_00115_, _00114_, _26752_);
  nor (_00116_, _00115_, _26773_);
  nor (_00117_, _00116_, _26843_);
  not (_00118_, _00117_);
  and (_00119_, _00004_, _26072_);
  nand (_00120_, _00102_, _25916_);
  and (_00121_, _26676_, _00043_);
  nor (_00122_, _22768_, _23130_);
  and (_00123_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00124_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_00125_, _00124_, _00123_);
  and (_00126_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00127_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_00128_, _00127_, _00126_);
  and (_00129_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_00130_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_00131_, _00130_, _00129_);
  and (_00132_, _00131_, _00128_);
  and (_00133_, _00132_, _00125_);
  nor (_00135_, _00133_, _25562_);
  nor (_00136_, _00135_, _00122_);
  not (_00137_, _00136_);
  and (_00138_, _00137_, _26834_);
  nor (_00140_, _00138_, _00121_);
  nand (_00141_, _00140_, _00120_);
  nor (_00143_, _00141_, _00119_);
  and (_00144_, _00143_, _00118_);
  nor (_00145_, _00144_, _22951_);
  and (_00146_, _00144_, _22951_);
  nor (_00147_, _00146_, _00145_);
  nor (_00148_, _00147_, _00110_);
  and (_00149_, _00148_, _00072_);
  and (_00150_, _00149_, _00033_);
  nor (_00151_, _24671_, _23881_);
  and (_00152_, _00151_, _00150_);
  and (_00153_, _00152_, _26640_);
  not (_00155_, _00153_);
  and (_00156_, _00004_, _26016_);
  not (_00158_, _00156_);
  not (_00159_, _25641_);
  and (_00160_, _00007_, _00159_);
  nor (_00161_, _26765_, _26760_);
  nor (_00163_, _00161_, _26766_);
  nor (_00165_, _00163_, _22861_);
  nor (_00166_, _00165_, _22956_);
  nor (_00168_, _00166_, _26752_);
  nor (_00169_, _00168_, _26758_);
  not (_00170_, _00169_);
  nand (_00171_, _00170_, _26842_);
  and (_00172_, _00102_, _24268_);
  nor (_00173_, _00172_, _00044_);
  nand (_00174_, _00173_, _00171_);
  nor (_00175_, _00174_, _00160_);
  and (_00176_, _00175_, _00158_);
  and (_00177_, _00176_, _23990_);
  nor (_00178_, _00176_, _23990_);
  or (_00179_, _00178_, _00177_);
  nor (_00180_, _00179_, _25129_);
  nor (_00181_, _26764_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_00182_, _00181_, _26765_);
  nor (_00183_, _00182_, _22861_);
  nor (_00184_, _00183_, _22922_);
  nor (_00185_, _00184_, _26752_);
  not (_00186_, _00185_);
  and (_00187_, _00186_, _26762_);
  not (_00188_, _00187_);
  nand (_00189_, _00188_, _26842_);
  nand (_00190_, _00102_, _24413_);
  and (_00191_, _00190_, _00189_);
  nand (_00192_, _00004_, _25994_);
  not (_00193_, _25767_);
  nand (_00194_, _00007_, _00193_);
  and (_00195_, _00194_, _00192_);
  and (_00196_, _00195_, _00191_);
  nor (_00197_, _00196_, _22926_);
  and (_00198_, _00196_, _22926_);
  nor (_00199_, _00198_, _00197_);
  and (_00200_, _00102_, _24294_);
  not (_00201_, _25565_);
  and (_00202_, _00007_, _00201_);
  nor (_00203_, _00202_, _00200_);
  and (_00204_, _00004_, _26035_);
  and (_00205_, _26767_, _26757_);
  nor (_00206_, _00205_, _26768_);
  nor (_00207_, _00206_, _22861_);
  nor (_00208_, _00207_, _23003_);
  nor (_00209_, _00208_, _26752_);
  nor (_00210_, _00209_, _26754_);
  not (_00211_, _00210_);
  and (_00212_, _00211_, _26842_);
  nor (_00213_, _00212_, _00204_);
  and (_00214_, _00213_, _00203_);
  nor (_00215_, _00214_, _23012_);
  and (_00216_, _00214_, _23012_);
  nor (_00217_, _00216_, _00215_);
  nor (_00218_, _00217_, _00199_);
  and (_00219_, _00218_, _00180_);
  and (_00220_, _00219_, _00150_);
  and (_00221_, _22890_, _22856_);
  and (_00222_, _00221_, _00220_);
  not (_00223_, _00222_);
  not (_00224_, _26571_);
  not (_00225_, _24496_);
  nand (_00226_, _24451_, _24445_);
  or (_00227_, _00226_, _00225_);
  and (_00228_, _26644_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not (_00229_, _00228_);
  nor (_00230_, _23452_, _23417_);
  nor (_00231_, _00230_, _23453_);
  and (_00232_, _23455_, _23389_);
  nor (_00233_, _23455_, _23389_);
  nor (_00234_, _00233_, _00232_);
  nor (_00235_, _23453_, _23414_);
  nor (_00236_, _00235_, _23454_);
  nor (_00237_, _23451_, _23155_);
  and (_00238_, _23451_, _23155_);
  nor (_00239_, _00238_, _00237_);
  and (_00240_, _23443_, _23432_);
  nor (_00241_, _00240_, _23444_);
  nor (_00242_, _23441_, _23435_);
  nor (_00244_, _00242_, _23442_);
  and (_00245_, _00244_, _23438_);
  nand (_00246_, _00245_, _00241_);
  or (_00247_, _26633_, _26560_);
  or (_00248_, _00247_, _00246_);
  nor (_00249_, _00248_, _00239_);
  nand (_00250_, _00249_, _00236_);
  or (_00251_, _00250_, _26646_);
  nor (_00252_, _00251_, _00234_);
  and (_00253_, _00252_, _00231_);
  and (_00254_, _26646_, _26634_);
  and (_00255_, _00254_, _23324_);
  nor (_00256_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_00257_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_00258_, _00257_, _00256_);
  nor (_00259_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_00260_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00261_, _00260_, _00259_);
  and (_00262_, _00261_, _00258_);
  and (_00263_, _00262_, _26647_);
  nor (_00264_, _00263_, _00255_);
  not (_00265_, _00264_);
  nor (_00267_, _00265_, _00253_);
  and (_00268_, _00267_, _00229_);
  nor (_00269_, _00268_, _26590_);
  and (_00270_, _00269_, _00227_);
  or (_00271_, _26656_, _24458_);
  and (_00272_, _00271_, _24447_);
  and (_00273_, _26619_, _24443_);
  and (_00274_, _26609_, _24443_);
  or (_00275_, _00274_, _00273_);
  nor (_00276_, _00275_, _00272_);
  and (_00277_, _00276_, _26618_);
  and (_00279_, _00277_, _00268_);
  nor (_00280_, _00279_, _00270_);
  not (_00281_, _26607_);
  and (_00282_, _26623_, _00281_);
  not (_00283_, _00282_);
  nor (_00284_, _00283_, _00280_);
  nor (_00285_, _00284_, _00224_);
  nor (_00286_, _26608_, _26582_);
  not (_00287_, _00286_);
  nor (_00288_, _00287_, _00285_);
  nor (_00289_, _26639_, _26634_);
  not (_00290_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_00291_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _22765_);
  and (_00292_, _00291_, _00290_);
  not (_00293_, _00292_);
  not (_00294_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_00295_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _22765_);
  and (_00296_, _00295_, _00294_);
  and (_00297_, _24711_, _24571_);
  and (_00298_, _00297_, _25769_);
  nor (_00299_, _00298_, _00296_);
  and (_00300_, _00299_, _00293_);
  nor (_00301_, _22998_, _22981_);
  and (_00302_, _00301_, _24629_);
  and (_00303_, _00302_, _25208_);
  not (_00304_, _00303_);
  and (_00305_, _00304_, _00300_);
  not (_00306_, _00305_);
  and (_00307_, _00306_, _00289_);
  nor (_00308_, _22999_, _22981_);
  and (_00309_, _00308_, _24629_);
  and (_00310_, _00309_, _25117_);
  nor (_00311_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_00312_, _00311_);
  nor (_00313_, _00312_, _00310_);
  and (_00314_, _00313_, _25772_);
  nor (_00315_, _00314_, _26637_);
  nor (_00316_, _00315_, _00307_);
  not (_00317_, _00316_);
  nor (_00318_, _00317_, _00288_);
  and (_00319_, _00318_, _00223_);
  and (_00320_, _00319_, _00155_);
  or (_00321_, _26628_, _26610_);
  or (_00322_, _26615_, _26583_);
  and (_00323_, _00322_, _00321_);
  and (_00324_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_00325_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_00326_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00327_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00328_, _00327_, _00326_);
  and (_00330_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00331_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_00332_, _00331_, _00330_);
  and (_00333_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_00334_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_00335_, _00334_, _00333_);
  or (_00336_, _00335_, _00332_);
  or (_00337_, _00336_, _00328_);
  and (_00338_, _00337_, _24270_);
  or (_00339_, _00338_, _00325_);
  and (_00340_, _00339_, _22768_);
  nor (_00341_, _00340_, _00324_);
  nor (_00342_, _00341_, _26614_);
  and (_00343_, _26614_, _00193_);
  or (_00344_, _00343_, _00342_);
  nor (_00345_, _00344_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00346_, _00344_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00347_, _00346_, _00345_);
  and (_00348_, _00347_, _00323_);
  nor (_00349_, _00322_, _26628_);
  and (_00350_, _00349_, _00193_);
  nor (_00351_, _00341_, _26605_);
  and (_00352_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00353_, _00352_, _00351_);
  or (_00354_, _00353_, _00350_);
  nor (_00355_, _00354_, _00348_);
  nand (_00356_, _00355_, _00320_);
  or (_00357_, _00356_, _26632_);
  or (_00358_, _00320_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00359_, _00358_, _22761_);
  and (_26899_[0], _00359_, _00357_);
  and (_00360_, _26341_, _26340_);
  not (_00361_, _00360_);
  and (_00362_, _00361_, _26342_);
  or (_00363_, _00362_, _26368_);
  and (_00364_, _26367_, _26172_);
  or (_00365_, _00364_, _26337_);
  and (_00366_, _00365_, _00363_);
  nand (_00367_, _00366_, _23528_);
  not (_00368_, _26541_);
  nor (_00369_, _26544_, _00368_);
  and (_00370_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and (_00371_, _26535_, _26467_);
  nand (_00372_, _00371_, _26538_);
  nand (_00373_, _00372_, _00370_);
  or (_00374_, _00372_, _00370_);
  nand (_00375_, _00374_, _00373_);
  or (_00376_, _00375_, _00369_);
  nand (_00377_, _00375_, _00369_);
  and (_00378_, _00377_, _00376_);
  nand (_00379_, _00378_, _23531_);
  nor (_00380_, _23464_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_00381_, _00380_, _23242_);
  nor (_00382_, _00380_, _23242_);
  nor (_00383_, _00382_, _00381_);
  nor (_00384_, _00383_, _23462_);
  not (_00385_, _23536_);
  nor (_00386_, _00385_, _23271_);
  not (_00387_, _00386_);
  nand (_00388_, _23534_, _23211_);
  and (_00389_, _23494_, _23242_);
  not (_00390_, _00389_);
  and (_00391_, _00390_, _00388_);
  and (_00392_, _00391_, _00387_);
  not (_00393_, _00392_);
  nor (_00394_, _00393_, _00384_);
  and (_00395_, _00394_, _23783_);
  nor (_00396_, _23281_, _23279_);
  or (_00397_, _00396_, _23282_);
  and (_00398_, _00397_, _23334_);
  nor (_00399_, _00397_, _23334_);
  or (_00400_, _00399_, _00398_);
  and (_00401_, _00400_, _23037_);
  nor (_00402_, _23440_, _23438_);
  nor (_00403_, _00402_, _23441_);
  nor (_00404_, _00403_, _23399_);
  nor (_00405_, _00404_, _00401_);
  and (_00406_, _00405_, _00395_);
  and (_00407_, _00406_, _00379_);
  nand (_00408_, _00407_, _00367_);
  and (_00409_, _00408_, _26631_);
  and (_00410_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00411_, _00349_, _00159_);
  and (_00412_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_00413_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_00415_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00416_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00417_, _00416_, _00415_);
  and (_00418_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00419_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_00421_, _00419_, _00418_);
  and (_00422_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_00423_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_00424_, _00423_, _00422_);
  or (_00425_, _00424_, _00421_);
  or (_00426_, _00425_, _00417_);
  and (_00427_, _00426_, _24270_);
  or (_00428_, _00427_, _00413_);
  and (_00429_, _00428_, _22768_);
  nor (_00430_, _00429_, _00412_);
  nor (_00431_, _00430_, _26605_);
  or (_00432_, _00431_, _00411_);
  or (_00433_, _00432_, _00410_);
  or (_00434_, _00433_, _00409_);
  or (_00435_, _00430_, _26614_);
  nand (_00436_, _26614_, _00159_);
  and (_00437_, _00436_, _00435_);
  or (_00438_, _00437_, _23222_);
  nand (_00439_, _00437_, _23222_);
  and (_00440_, _00439_, _00438_);
  nor (_00441_, _00440_, _00346_);
  and (_00442_, _00440_, _00346_);
  nor (_00443_, _00442_, _00441_);
  nand (_00444_, _00443_, _00323_);
  nand (_00445_, _00444_, _00320_);
  or (_00446_, _00445_, _00434_);
  or (_00447_, _00320_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00448_, _00447_, _22761_);
  and (_26899_[1], _00448_, _00446_);
  not (_00449_, _26353_);
  and (_00450_, _26352_, _26343_);
  nor (_00451_, _00450_, _00449_);
  or (_00452_, _00451_, _26368_);
  or (_00453_, _00364_, _26349_);
  and (_00454_, _00453_, _00452_);
  nand (_00455_, _00454_, _23528_);
  and (_00456_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  nand (_00457_, _00376_, _00373_);
  nand (_00458_, _00457_, _00456_);
  or (_00459_, _00457_, _00456_);
  and (_00461_, _00459_, _00458_);
  nand (_00462_, _00461_, _23531_);
  nor (_00463_, _00244_, _23399_);
  nand (_00464_, _23536_, _23242_);
  and (_00465_, _23494_, _23211_);
  not (_00466_, _00465_);
  or (_00467_, _23535_, _23178_);
  and (_00468_, _00467_, _00466_);
  and (_00469_, _00468_, _00464_);
  and (_00470_, _00469_, _23706_);
  not (_00471_, _00470_);
  nor (_00472_, _00471_, _00463_);
  nor (_00473_, _23338_, _23335_);
  nor (_00474_, _00473_, _23038_);
  and (_00475_, _00474_, _23340_);
  and (_00476_, _23463_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00477_, _00382_, _23684_);
  nor (_00478_, _00477_, _00476_);
  nor (_00479_, _00478_, _23462_);
  nor (_00480_, _00479_, _00475_);
  and (_00481_, _00480_, _00472_);
  and (_00482_, _00481_, _23696_);
  and (_00483_, _00482_, _00462_);
  nand (_00484_, _00483_, _00455_);
  and (_00485_, _00484_, _26631_);
  not (_00486_, _00438_);
  or (_00487_, _00442_, _00486_);
  and (_00488_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_00489_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_00490_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00491_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00492_, _00491_, _00490_);
  and (_00493_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00494_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_00495_, _00494_, _00493_);
  or (_00496_, _00495_, _00492_);
  and (_00497_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00498_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00499_, _00498_, _00497_);
  or (_00500_, _00499_, _00496_);
  and (_00501_, _00500_, _24270_);
  or (_00502_, _00501_, _00489_);
  and (_00503_, _00502_, _22768_);
  nor (_00504_, _00503_, _00488_);
  nor (_00505_, _00504_, _26614_);
  and (_00506_, _26614_, _00201_);
  nor (_00507_, _00506_, _00505_);
  nor (_00508_, _00507_, _23192_);
  and (_00509_, _00507_, _23192_);
  nor (_00510_, _00509_, _00508_);
  nor (_00512_, _00510_, _00487_);
  and (_00513_, _00510_, _00487_);
  nor (_00514_, _00513_, _00512_);
  and (_00516_, _00514_, _00323_);
  and (_00517_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00518_, _00504_, _26605_);
  and (_00519_, _00349_, _00201_);
  or (_00520_, _00519_, _00518_);
  or (_00521_, _00520_, _00517_);
  nor (_00522_, _00521_, _00516_);
  nand (_00523_, _00522_, _00320_);
  or (_00524_, _00523_, _00485_);
  not (_00525_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00526_, _25781_, _00525_);
  and (_00527_, _25781_, _00525_);
  nor (_00528_, _00527_, _00526_);
  or (_00529_, _00528_, _00320_);
  and (_00530_, _00529_, _22761_);
  and (_26899_[2], _00530_, _00524_);
  or (_00531_, _26354_, _26330_);
  and (_00532_, _26353_, _26350_);
  nor (_00533_, _00532_, _00531_);
  and (_00534_, _00532_, _00531_);
  nor (_00535_, _00534_, _00533_);
  or (_00536_, _00535_, _26368_);
  or (_00537_, _00364_, _26329_);
  and (_00538_, _00537_, _00536_);
  nand (_00539_, _00538_, _23528_);
  or (_00540_, _00375_, _26541_);
  nand (_00541_, _00540_, _00373_);
  and (_00542_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_00543_, _00542_, _00456_);
  and (_00544_, _00543_, _00541_);
  and (_00545_, _00374_, _00373_);
  and (_00546_, _00545_, _26543_);
  and (_00547_, _00543_, _00546_);
  and (_00548_, _00547_, _26528_);
  or (_00549_, _00548_, _00544_);
  not (_00550_, _00549_);
  not (_00551_, _00542_);
  nand (_00552_, _00551_, _00458_);
  and (_00553_, _00552_, _00550_);
  nand (_00554_, _00553_, _23531_);
  nor (_00555_, _00241_, _23399_);
  not (_00556_, _00555_);
  and (_00557_, _23340_, _23288_);
  or (_00558_, _00557_, _23038_);
  nor (_00559_, _00558_, _23341_);
  not (_00560_, _00559_);
  not (_00561_, _23829_);
  or (_00562_, _23535_, _23146_);
  nand (_00563_, _23536_, _23211_);
  nor (_00564_, _26552_, _23178_);
  not (_00565_, _00564_);
  and (_00566_, _00565_, _00563_);
  and (_00567_, _00566_, _00562_);
  and (_00568_, _00567_, _23825_);
  not (_00569_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00570_, _23463_, _00569_);
  nor (_00571_, _00570_, _23552_);
  or (_00572_, _00571_, _23462_);
  or (_00573_, _00572_, _23464_);
  and (_00574_, _00573_, _00568_);
  and (_00575_, _00574_, _00561_);
  and (_00576_, _00575_, _23822_);
  and (_00577_, _00576_, _00560_);
  and (_00578_, _00577_, _00556_);
  and (_00579_, _00578_, _00554_);
  nand (_00580_, _00579_, _00539_);
  and (_00581_, _00580_, _26631_);
  and (_00582_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00583_, _26605_, _25663_);
  and (_00584_, _00349_, _00091_);
  or (_00585_, _00584_, _00583_);
  or (_00586_, _00585_, _00582_);
  or (_00587_, _00513_, _00508_);
  nor (_00588_, _26614_, _25663_);
  and (_00589_, _00091_, _26614_);
  nor (_00590_, _00589_, _00588_);
  nor (_00591_, _00590_, _23156_);
  and (_00593_, _00590_, _23156_);
  nor (_00594_, _00593_, _00591_);
  nand (_00595_, _00594_, _00587_);
  or (_00596_, _00594_, _00587_);
  and (_00597_, _00596_, _00595_);
  and (_00598_, _00597_, _00323_);
  or (_00599_, _00598_, _00586_);
  or (_00600_, _00599_, _00581_);
  and (_00601_, _00600_, _00320_);
  not (_00602_, _00320_);
  and (_00603_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not (_00604_, _00603_);
  nor (_00605_, _00604_, _25781_);
  nor (_00606_, _00526_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00607_, _00606_, _00605_);
  and (_00608_, _00607_, _00602_);
  or (_00609_, _00608_, _00601_);
  and (_26899_[3], _00609_, _22761_);
  and (_00610_, _00605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00611_, _00605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00612_, _00611_, _00610_);
  nor (_00613_, _00612_, _00320_);
  and (_00614_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00615_, _26362_, _26358_);
  nand (_00616_, _26362_, _26358_);
  and (_00617_, _00616_, _00615_);
  or (_00618_, _00617_, _26368_);
  or (_00619_, _00364_, _26316_);
  and (_00620_, _00619_, _00618_);
  and (_00621_, _00620_, _23528_);
  and (_00622_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_00623_, _00622_, _00549_);
  nor (_00624_, _00622_, _00549_);
  nor (_00625_, _00624_, _00623_);
  and (_00626_, _00625_, _23531_);
  and (_00627_, _00239_, _23398_);
  or (_00628_, _23345_, _23155_);
  nor (_00629_, _23346_, _23038_);
  and (_00630_, _00629_, _00628_);
  and (_00631_, _23464_, _23461_);
  and (_00632_, _00631_, _23551_);
  not (_00633_, _00632_);
  or (_00634_, _00631_, _23551_);
  and (_00635_, _00634_, _23461_);
  and (_00636_, _00635_, _00633_);
  nor (_00637_, _26552_, _23146_);
  and (_00638_, _23534_, _23115_);
  nor (_00639_, _00385_, _23178_);
  or (_00640_, _00639_, _00638_);
  or (_00641_, _00640_, _00637_);
  or (_00642_, _00641_, _00636_);
  or (_00643_, _00642_, _23913_);
  or (_00644_, _00643_, _00630_);
  or (_00645_, _00644_, _00627_);
  or (_00646_, _00645_, _00626_);
  or (_00647_, _00646_, _00621_);
  and (_00648_, _00647_, _26631_);
  and (_00649_, _00137_, _26614_);
  nor (_00650_, _26614_, _25584_);
  nor (_00651_, _00650_, _00649_);
  or (_00652_, _00651_, _23125_);
  nand (_00653_, _00651_, _23125_);
  and (_00654_, _00653_, _00652_);
  nor (_00655_, _00591_, _00587_);
  nor (_00656_, _00655_, _00593_);
  or (_00657_, _00656_, _00654_);
  nand (_00658_, _00656_, _00654_);
  and (_00659_, _00658_, _00323_);
  and (_00660_, _00659_, _00657_);
  and (_00661_, _00349_, _00137_);
  and (_00662_, _00650_, _26582_);
  or (_00663_, _00662_, _00661_);
  or (_00664_, _00663_, _00660_);
  or (_00665_, _00664_, _00648_);
  or (_00666_, _00665_, _00614_);
  and (_00667_, _00666_, _00320_);
  or (_00668_, _00667_, _00613_);
  and (_26899_[4], _00668_, _22761_);
  and (_00669_, _00615_, _26318_);
  nand (_00670_, _26320_, _00669_);
  or (_00671_, _26320_, _00669_);
  and (_00672_, _00671_, _00670_);
  or (_00673_, _00672_, _26368_);
  or (_00674_, _00364_, _26309_);
  and (_00675_, _00674_, _00673_);
  and (_00676_, _00675_, _23528_);
  and (_00677_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_00678_, _00677_, _00622_);
  nand (_00679_, _00678_, _00549_);
  or (_00680_, _00677_, _00623_);
  and (_00682_, _00680_, _00679_);
  and (_00683_, _00682_, _23531_);
  nor (_00684_, _23153_, _23124_);
  nor (_00685_, _00684_, _23378_);
  or (_00686_, _00685_, _23346_);
  nor (_00687_, _23347_, _23038_);
  and (_00688_, _00687_, _00686_);
  nor (_00689_, _00231_, _23399_);
  nor (_00690_, _00631_, _23471_);
  and (_00691_, _00690_, _23468_);
  nor (_00692_, _00691_, _00632_);
  and (_00693_, _00692_, _23469_);
  nor (_00694_, _00692_, _23469_);
  or (_00695_, _00694_, _00693_);
  and (_00696_, _00695_, _23461_);
  nor (_00697_, _23535_, _23366_);
  nand (_00698_, _23494_, _23115_);
  or (_00699_, _00385_, _23146_);
  nand (_00700_, _00699_, _00698_);
  nor (_00701_, _00700_, _00697_);
  nand (_00702_, _00701_, _23623_);
  nor (_00703_, _00702_, _00696_);
  nand (_00704_, _00703_, _23616_);
  or (_00705_, _00704_, _00689_);
  or (_00706_, _00705_, _00688_);
  or (_00707_, _00706_, _00683_);
  or (_00708_, _00707_, _00676_);
  and (_00709_, _00708_, _26631_);
  and (_00710_, _00349_, _00022_);
  and (_00711_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_00712_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_00713_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00714_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00715_, _00714_, _00713_);
  and (_00716_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00717_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or (_00718_, _00717_, _00716_);
  or (_00719_, _00718_, _00715_);
  and (_00720_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00721_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00722_, _00721_, _00720_);
  or (_00723_, _00722_, _00719_);
  and (_00724_, _00723_, _24270_);
  or (_00725_, _00724_, _00712_);
  and (_00726_, _00725_, _22768_);
  nor (_00727_, _00726_, _00711_);
  nor (_00728_, _00727_, _26605_);
  and (_00729_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00730_, _00729_, _00728_);
  or (_00731_, _00730_, _00710_);
  nand (_00732_, _00658_, _00652_);
  nor (_00733_, _00727_, _26614_);
  and (_00734_, _00022_, _26614_);
  nor (_00735_, _00734_, _00733_);
  nor (_00736_, _00735_, _23093_);
  and (_00737_, _00735_, _23093_);
  nor (_00738_, _00737_, _00736_);
  nor (_00739_, _00738_, _00732_);
  and (_00740_, _00738_, _00732_);
  nor (_00742_, _00740_, _00739_);
  and (_00744_, _00742_, _00323_);
  nor (_00745_, _00744_, _00731_);
  nand (_00746_, _00745_, _00320_);
  or (_00747_, _00746_, _00709_);
  and (_00748_, _00610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00749_, _00610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00750_, _00749_, _00748_);
  or (_00751_, _00750_, _00320_);
  and (_00752_, _00751_, _22761_);
  and (_26899_[5], _00752_, _00747_);
  not (_00753_, _26301_);
  and (_00754_, _26365_, _00753_);
  nor (_00755_, _26365_, _00753_);
  or (_00756_, _00755_, _00754_);
  and (_00757_, _00756_, _00364_);
  and (_00758_, _26368_, _26295_);
  or (_00759_, _00758_, _00757_);
  or (_00760_, _00759_, _23529_);
  not (_00761_, _23531_);
  and (_00762_, _26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not (_00763_, _00762_);
  nor (_00764_, _00763_, _00679_);
  and (_00765_, _00763_, _00679_);
  or (_00766_, _00765_, _00764_);
  or (_00767_, _00766_, _00761_);
  nor (_00768_, _00236_, _23399_);
  not (_00769_, _00768_);
  nor (_00770_, _23382_, _23347_);
  nor (_00771_, _00770_, _23038_);
  and (_00772_, _00771_, _23384_);
  nor (_00773_, _00693_, _23366_);
  and (_00774_, _00693_, _23366_);
  nor (_00775_, _00774_, _00773_);
  nor (_00776_, _00775_, _23462_);
  or (_00777_, _23535_, _23078_);
  nand (_00778_, _23536_, _23115_);
  nor (_00779_, _26552_, _23366_);
  not (_00780_, _00779_);
  and (_00781_, _00780_, _00778_);
  and (_00782_, _00781_, _00777_);
  and (_00783_, _00782_, _23744_);
  not (_00784_, _00783_);
  nor (_00785_, _00784_, _00776_);
  and (_00786_, _00785_, _23737_);
  not (_00787_, _00786_);
  nor (_00788_, _00787_, _00772_);
  and (_00789_, _00788_, _00769_);
  and (_00790_, _00789_, _00767_);
  and (_00791_, _00790_, _00760_);
  not (_00792_, _00791_);
  and (_00793_, _00792_, _26631_);
  or (_00794_, _00740_, _00736_);
  and (_00795_, _25566_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_00796_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_00797_, _24239_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00798_, _24250_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00799_, _00798_, _00797_);
  and (_00800_, _24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00801_, _24243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_00802_, _00801_, _00800_);
  or (_00803_, _00802_, _00799_);
  and (_00804_, _24253_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00805_, _24255_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00806_, _00805_, _00804_);
  or (_00807_, _00806_, _00803_);
  and (_00809_, _00807_, _24270_);
  or (_00810_, _00809_, _00796_);
  and (_00811_, _00810_, _22768_);
  nor (_00812_, _00811_, _00795_);
  not (_00813_, _00812_);
  nor (_00814_, _00813_, _26614_);
  and (_00815_, _00061_, _26614_);
  nor (_00816_, _00815_, _00814_);
  nand (_00817_, _00816_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_00818_, _00816_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00819_, _00818_, _00817_);
  nand (_00820_, _00819_, _00794_);
  or (_00821_, _00819_, _00794_);
  and (_00822_, _00821_, _00323_);
  and (_00824_, _00822_, _00820_);
  and (_00825_, _00813_, _26604_);
  and (_00826_, _00349_, _00062_);
  and (_00827_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00828_, _00827_, _00826_);
  or (_00829_, _00828_, _00825_);
  or (_00830_, _00829_, _00824_);
  or (_00831_, _00830_, _00793_);
  and (_00832_, _00831_, _00320_);
  and (_00833_, _00748_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00834_, _00748_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00835_, _00834_, _00833_);
  nor (_00836_, _00835_, _00320_);
  or (_00837_, _00836_, _00832_);
  and (_26899_[6], _00837_, _22761_);
  or (_00838_, _00364_, _26286_);
  not (_00839_, _26296_);
  or (_00840_, _00754_, _00839_);
  and (_00841_, _00840_, _26299_);
  or (_00842_, _00841_, _26368_);
  and (_00843_, _00842_, _00838_);
  and (_00844_, _00843_, _23528_);
  not (_00845_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or (_00846_, _26375_, _00845_);
  nor (_00847_, _00846_, _00764_);
  and (_00848_, _00764_, _00845_);
  or (_00849_, _00848_, _00847_);
  and (_00850_, _00849_, _23531_);
  and (_00851_, _00234_, _23398_);
  nand (_00852_, _23389_, _23386_);
  and (_00853_, _00852_, _23390_);
  and (_00855_, _00853_, _23037_);
  and (_00856_, _00633_, _23470_);
  nor (_00857_, _00691_, _00856_);
  nor (_00858_, _00857_, _23078_);
  and (_00859_, _00857_, _23078_);
  or (_00860_, _00859_, _00858_);
  and (_00861_, _00860_, _23461_);
  and (_00862_, _23506_, _23330_);
  and (_00863_, _23501_, _23505_);
  nor (_00864_, _26552_, _23078_);
  nor (_00865_, _00385_, _23366_);
  or (_00866_, _00865_, _00864_);
  or (_00867_, _00866_, _00863_);
  or (_00868_, _00867_, _00862_);
  nor (_00869_, _00868_, _00861_);
  nand (_00870_, _00869_, _23584_);
  or (_00871_, _00870_, _00855_);
  or (_00872_, _00871_, _00851_);
  or (_00873_, _00872_, _00850_);
  or (_00874_, _00873_, _00844_);
  and (_00875_, _00874_, _26631_);
  nand (_00876_, _00820_, _00817_);
  nor (_00877_, _26614_, _25605_);
  and (_00878_, _26614_, _26833_);
  nor (_00879_, _00878_, _00877_);
  nor (_00880_, _00879_, _23039_);
  and (_00881_, _00879_, _23039_);
  nor (_00882_, _00881_, _00880_);
  nand (_00883_, _00882_, _00876_);
  or (_00884_, _00882_, _00876_);
  and (_00885_, _00884_, _00323_);
  and (_00886_, _00885_, _00883_);
  and (_00887_, _00349_, _26833_);
  and (_00888_, _26608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00889_, _26605_, _25605_);
  or (_00890_, _00889_, _00888_);
  or (_00891_, _00890_, _00887_);
  nor (_00892_, _00891_, _00886_);
  nand (_00893_, _00892_, _00320_);
  or (_00894_, _00893_, _00875_);
  nor (_00895_, _00833_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00896_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_00897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00899_, _00897_, _00896_);
  and (_00900_, _00899_, _00603_);
  not (_00901_, _00900_);
  nor (_00902_, _00901_, _25781_);
  nor (_00903_, _00902_, _00895_);
  or (_00904_, _00903_, _00320_);
  and (_00905_, _00904_, _22761_);
  and (_26899_[7], _00905_, _00894_);
  and (_00906_, _26608_, _26568_);
  not (_00907_, _00879_);
  nor (_00908_, _00880_, _00876_);
  nor (_00909_, _00908_, _00881_);
  nand (_00910_, _00909_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_00911_, _00909_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00912_, _00911_, _00910_);
  or (_00914_, _00912_, _00907_);
  nand (_00915_, _00912_, _00907_);
  and (_00916_, _00915_, _00914_);
  and (_00917_, _00916_, _00323_);
  not (_00918_, _26574_);
  and (_00919_, _00364_, _23528_);
  not (_00920_, _00919_);
  nor (_00921_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_00922_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_00923_, _00922_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00924_, _00923_, _00921_);
  not (_00925_, _00924_);
  or (_00926_, _00925_, _23391_);
  and (_00927_, _00925_, _23391_);
  nor (_00928_, _00927_, _23038_);
  and (_00929_, _00928_, _00926_);
  and (_00930_, _23330_, _23508_);
  nor (_00931_, _23570_, _00930_);
  not (_00932_, _00931_);
  nor (_00933_, _00932_, _23561_);
  nor (_00934_, _00933_, _23419_);
  and (_00935_, _00933_, _23419_);
  or (_00936_, _00935_, _23544_);
  nor (_00937_, _00936_, _00934_);
  and (_00938_, _23494_, _23419_);
  and (_00939_, _26401_, _23505_);
  and (_00940_, _00939_, _23531_);
  and (_00941_, _23509_, _23551_);
  nor (_00942_, _23569_, _23271_);
  or (_00943_, _00942_, _00941_);
  or (_00944_, _00943_, _00940_);
  nor (_00945_, _00944_, _00938_);
  not (_00946_, _00945_);
  nor (_00947_, _00946_, _00937_);
  not (_00948_, _00947_);
  nor (_00949_, _00948_, _00929_);
  and (_00950_, _00949_, _00920_);
  nor (_00951_, _00950_, _00918_);
  and (_00952_, _26604_, _00193_);
  not (_00953_, _24385_);
  and (_00954_, _00349_, _00953_);
  and (_00955_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00956_, _00955_, _00954_);
  or (_00957_, _00956_, _00952_);
  or (_00958_, _00957_, _00951_);
  or (_00959_, _00958_, _00917_);
  or (_00960_, _00959_, _00906_);
  or (_00961_, _00960_, _00602_);
  and (_00962_, _00902_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00963_, _00902_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00964_, _00963_, _00962_);
  or (_00965_, _00964_, _00320_);
  and (_00966_, _00965_, _22761_);
  and (_26899_[8], _00966_, _00961_);
  not (_00967_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_00968_, _00910_, _00907_);
  nor (_00969_, _00911_, _00879_);
  nor (_00970_, _00969_, _00968_);
  nand (_00971_, _00970_, _00967_);
  or (_00972_, _00970_, _00967_);
  and (_00973_, _00972_, _00971_);
  and (_00974_, _00973_, _00323_);
  and (_00975_, _00408_, _26608_);
  nor (_00976_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00977_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _00967_);
  nor (_00978_, _00977_, _00976_);
  not (_00979_, _00978_);
  and (_00980_, _00979_, _00926_);
  not (_00981_, _00980_);
  or (_00982_, _00979_, _00926_);
  and (_00983_, _00982_, _23037_);
  and (_00984_, _00983_, _00981_);
  not (_00985_, _00984_);
  and (_00986_, _26272_, _23528_);
  not (_00987_, _00986_);
  nor (_00988_, _23278_, _23078_);
  and (_00989_, _00988_, _23558_);
  nand (_00990_, _00989_, _23468_);
  and (_00991_, _23278_, _23078_);
  and (_00992_, _00991_, _23548_);
  nand (_00993_, _00992_, _23330_);
  and (_00994_, _00993_, _00990_);
  nor (_00995_, _00994_, _23248_);
  and (_00996_, _00994_, _23248_);
  nor (_00997_, _00996_, _00995_);
  nor (_00998_, _00997_, _23544_);
  and (_00999_, _23494_, _23248_);
  and (_01000_, _26440_, _26406_);
  nor (_01001_, _01000_, _26441_);
  and (_01002_, _01001_, _23531_);
  and (_01003_, _23509_, _23115_);
  and (_01004_, _23568_, _23242_);
  or (_01005_, _01004_, _01003_);
  or (_01006_, _01005_, _01002_);
  nor (_01007_, _01006_, _00999_);
  not (_01008_, _01007_);
  nor (_01009_, _01008_, _00998_);
  and (_01010_, _01009_, _00987_);
  and (_01011_, _01010_, _00985_);
  nor (_01012_, _01011_, _00918_);
  and (_01013_, _26604_, _00159_);
  not (_01014_, _24363_);
  and (_01015_, _00349_, _01014_);
  and (_01016_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_01017_, _01016_, _01015_);
  or (_01018_, _01017_, _01013_);
  or (_01019_, _01018_, _01012_);
  nor (_01020_, _01019_, _00975_);
  nand (_01021_, _01020_, _00320_);
  or (_01022_, _01021_, _00974_);
  and (_01023_, _00962_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_01024_, _00962_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_01025_, _01024_, _01023_);
  or (_01026_, _01025_, _00320_);
  and (_01027_, _01026_, _22761_);
  and (_26899_[9], _01027_, _01022_);
  not (_01028_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01029_, _00969_, _00967_);
  and (_01030_, _00968_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_01031_, _01030_, _01029_);
  nand (_01032_, _01031_, _01028_);
  or (_01033_, _01031_, _01028_);
  and (_01034_, _01033_, _01032_);
  and (_01035_, _01034_, _00323_);
  and (_01036_, _00484_, _26608_);
  nor (_01037_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01038_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _01028_);
  nor (_01040_, _01038_, _01037_);
  not (_01041_, _01040_);
  and (_01042_, _01041_, _00982_);
  not (_01043_, _01042_);
  or (_01044_, _01041_, _00982_);
  and (_01045_, _01044_, _23037_);
  and (_01046_, _01045_, _01043_);
  not (_01047_, _01046_);
  nor (_01048_, _00993_, _23248_);
  and (_01049_, _00989_, _23248_);
  and (_01050_, _01049_, _23468_);
  nor (_01051_, _01050_, _01048_);
  and (_01052_, _01051_, _23427_);
  nor (_01053_, _01051_, _23427_);
  or (_01054_, _01053_, _23544_);
  nor (_01055_, _01054_, _01052_);
  nor (_01056_, _26510_, _26507_);
  nor (_01057_, _01056_, _26511_);
  and (_01058_, _01057_, _23531_);
  and (_01059_, _23494_, _23217_);
  and (_01060_, _23509_, _23550_);
  and (_01061_, _23568_, _23211_);
  and (_01062_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_01063_, _01062_, _01061_);
  or (_01064_, _01063_, _01060_);
  nor (_01065_, _01064_, _01059_);
  not (_01066_, _01065_);
  nor (_01067_, _01066_, _01058_);
  not (_01068_, _01067_);
  nor (_01069_, _01068_, _01055_);
  and (_01071_, _01069_, _01047_);
  nor (_01072_, _01071_, _00918_);
  and (_01073_, _26604_, _00201_);
  not (_01074_, _24340_);
  and (_01075_, _00349_, _01074_);
  and (_01077_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_01078_, _01077_, _01075_);
  or (_01079_, _01078_, _01073_);
  or (_01080_, _01079_, _01072_);
  nor (_01081_, _01080_, _01036_);
  nand (_01082_, _01081_, _00320_);
  or (_01083_, _01082_, _01035_);
  nor (_01084_, _01023_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01085_, _01023_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01086_, _01085_, _01084_);
  or (_01087_, _01086_, _00320_);
  and (_01088_, _01087_, _22761_);
  and (_26899_[10], _01088_, _01083_);
  not (_01089_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_01090_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_01091_, _01090_, _00969_);
  nand (_01093_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_01094_, _01093_, _00910_);
  nor (_01096_, _01094_, _00907_);
  nor (_01098_, _01096_, _01091_);
  nand (_01099_, _01098_, _01089_);
  or (_01100_, _01098_, _01089_);
  and (_01101_, _01100_, _01099_);
  and (_01102_, _01101_, _00323_);
  and (_01103_, _00580_, _26608_);
  nor (_01104_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01105_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _01089_);
  nor (_01106_, _01105_, _01104_);
  not (_01107_, _01106_);
  and (_01108_, _01107_, _01044_);
  nor (_01109_, _01107_, _01044_);
  nor (_01110_, _01109_, _01108_);
  and (_01111_, _01110_, _23037_);
  not (_01112_, _01111_);
  and (_01113_, _26514_, _26512_);
  not (_01114_, _01113_);
  and (_01115_, _01114_, _26515_);
  and (_01117_, _01115_, _23531_);
  not (_01118_, _01117_);
  and (_01119_, _01049_, _23217_);
  and (_01120_, _01119_, _23468_);
  and (_01121_, _23423_, _23427_);
  and (_01122_, _01121_, _00992_);
  and (_01123_, _01122_, _23330_);
  nor (_01124_, _01123_, _01120_);
  nor (_01125_, _01124_, _23184_);
  and (_01126_, _01124_, _23184_);
  or (_01127_, _01126_, _23544_);
  nor (_01128_, _01127_, _01125_);
  and (_01129_, _23494_, _23445_);
  nor (_01130_, _01129_, _23510_);
  nor (_01131_, _23569_, _23178_);
  and (_01132_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_01133_, _01132_, _01131_);
  and (_01134_, _01133_, _01130_);
  not (_01135_, _01134_);
  nor (_01136_, _01135_, _01128_);
  and (_01137_, _01136_, _01118_);
  and (_01138_, _01137_, _01112_);
  nor (_01139_, _01138_, _00918_);
  and (_01140_, _00091_, _26604_);
  not (_01141_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_01143_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01144_, _01143_, _01142_);
  nor (_01145_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_01146_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01147_, _01146_, _01145_);
  not (_01148_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_01149_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _01148_);
  nor (_01150_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_01151_, _01150_, _01149_);
  and (_01152_, _01151_, _01147_);
  and (_01153_, _01152_, _01144_);
  nor (_01154_, _01153_, _01141_);
  and (_01155_, _01153_, _01141_);
  or (_01156_, _01155_, _01154_);
  and (_01157_, _01156_, _00349_);
  and (_01158_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_01159_, _01158_, _01157_);
  or (_01160_, _01159_, _01140_);
  nor (_01161_, _01160_, _01139_);
  nand (_01162_, _01161_, _00320_);
  or (_01163_, _01162_, _01103_);
  or (_01164_, _01163_, _01102_);
  and (_01165_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01166_, _01165_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01167_, _01166_, _00900_);
  and (_01168_, _01167_, _25845_);
  nor (_01169_, _01168_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01171_, _01168_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_01172_, _01171_, _01169_);
  or (_01173_, _01172_, _00320_);
  and (_01174_, _01173_, _22761_);
  and (_26899_[11], _01174_, _01164_);
  not (_01175_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01177_, _01090_, _01089_);
  and (_01178_, _01177_, _00969_);
  or (_01179_, _01094_, _01089_);
  nor (_01180_, _01179_, _00907_);
  nor (_01181_, _01180_, _01178_);
  nand (_01182_, _01181_, _01175_);
  or (_01183_, _01181_, _01175_);
  and (_01185_, _01183_, _01182_);
  and (_01187_, _01185_, _00323_);
  not (_01188_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01189_, _01155_, _01188_);
  and (_01190_, _01155_, _01188_);
  or (_01191_, _01190_, _01189_);
  and (_01192_, _01191_, _00349_);
  and (_01194_, _00647_, _26608_);
  nor (_01195_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01196_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _01175_);
  nor (_01197_, _01196_, _01195_);
  or (_01198_, _01197_, _01109_);
  and (_01199_, _01197_, _01109_);
  nor (_01200_, _01199_, _23038_);
  and (_01201_, _01200_, _01198_);
  or (_01203_, _26518_, _26516_);
  and (_01204_, _01203_, _26519_);
  and (_01205_, _01204_, _23531_);
  and (_01206_, _01123_, _23184_);
  and (_01207_, _01120_, _23445_);
  nor (_01208_, _01207_, _01206_);
  nand (_01209_, _01208_, _23152_);
  or (_01210_, _01208_, _23152_);
  and (_01211_, _01210_, _23543_);
  and (_01212_, _01211_, _01209_);
  and (_01213_, _23330_, _23551_);
  and (_01214_, _23468_, _23406_);
  or (_01216_, _01214_, _01213_);
  and (_01218_, _01216_, _23568_);
  and (_01219_, _23509_, _23505_);
  and (_01220_, _23494_, _23406_);
  and (_01222_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_01223_, _01222_, _01220_);
  or (_01224_, _01223_, _01219_);
  or (_01225_, _01224_, _01218_);
  or (_01226_, _01225_, _01212_);
  or (_01227_, _01226_, _01205_);
  or (_01228_, _01227_, _01201_);
  and (_01229_, _01228_, _26574_);
  and (_01230_, _00137_, _26604_);
  and (_01231_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_01232_, _01231_, _01230_);
  or (_01233_, _01232_, _01229_);
  or (_01234_, _01233_, _01194_);
  nor (_01235_, _01234_, _01192_);
  nand (_01236_, _01235_, _00320_);
  or (_01237_, _01236_, _01187_);
  nor (_01238_, _01171_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01239_, _01171_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01240_, _01239_, _01238_);
  or (_01241_, _01240_, _00320_);
  and (_01243_, _01241_, _22761_);
  and (_26899_[12], _01243_, _01237_);
  or (_01244_, _01179_, _01175_);
  or (_01245_, _01244_, _00907_);
  or (_01246_, _00911_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_01247_, _01246_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_01249_, _01247_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_01250_, _01249_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_01251_, _01250_, _00879_);
  nand (_01252_, _01251_, _01245_);
  nand (_01253_, _01252_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01254_, _01252_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01255_, _01254_, _00323_);
  and (_01257_, _01255_, _01253_);
  and (_01258_, _00708_, _26608_);
  nor (_01260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_01262_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01263_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _01262_);
  nor (_01264_, _01263_, _01260_);
  or (_01266_, _01264_, _01199_);
  nand (_01267_, _01264_, _01199_);
  and (_01268_, _01267_, _23037_);
  and (_01270_, _01268_, _01266_);
  or (_01271_, _26520_, _26496_);
  and (_01272_, _01271_, _26521_);
  and (_01273_, _01272_, _23531_);
  and (_01274_, _23445_, _23406_);
  and (_01275_, _01274_, _01119_);
  nand (_01276_, _01275_, _23468_);
  and (_01278_, _23184_, _23152_);
  and (_01280_, _01278_, _01122_);
  nand (_01281_, _01280_, _23330_);
  and (_01282_, _01281_, _01276_);
  nor (_01284_, _01282_, _23121_);
  and (_01285_, _01282_, _23121_);
  or (_01286_, _01285_, _01284_);
  and (_01287_, _01286_, _23543_);
  and (_01288_, _23468_, _23121_);
  and (_01289_, _23330_, _23115_);
  or (_01290_, _01289_, _01288_);
  and (_01291_, _01290_, _23568_);
  and (_01292_, _23509_, _23242_);
  and (_01293_, _23494_, _23121_);
  and (_01294_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_01295_, _01294_, _01293_);
  or (_01296_, _01295_, _01292_);
  or (_01297_, _01296_, _01291_);
  or (_01298_, _01297_, _01287_);
  or (_01299_, _01298_, _01273_);
  or (_01300_, _01299_, _01270_);
  and (_01301_, _01300_, _26574_);
  and (_01302_, _00022_, _26604_);
  not (_01303_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01304_, _01190_, _01303_);
  and (_01305_, _01190_, _01303_);
  or (_01306_, _01305_, _01304_);
  and (_01307_, _01306_, _00349_);
  and (_01308_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_01309_, _01308_, _01307_);
  or (_01311_, _01309_, _01302_);
  nor (_01312_, _01311_, _01301_);
  nand (_01313_, _01312_, _00320_);
  or (_01314_, _01313_, _01258_);
  or (_01315_, _01314_, _01257_);
  nor (_01316_, _01239_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_01317_, _01239_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01318_, _01317_, _01316_);
  or (_01319_, _01318_, _00320_);
  and (_01320_, _01319_, _22761_);
  and (_26899_[13], _01320_, _01315_);
  not (_01321_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01322_, _01305_, _01321_);
  and (_01323_, _01305_, _01321_);
  or (_01324_, _01323_, _01322_);
  and (_01325_, _01324_, _00349_);
  not (_01326_, _26608_);
  nor (_01327_, _00791_, _01326_);
  nor (_01328_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_01329_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01330_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _01329_);
  nor (_01331_, _01330_, _01328_);
  not (_01332_, _01331_);
  and (_01333_, _01332_, _01267_);
  not (_01334_, _01333_);
  or (_01335_, _01332_, _01267_);
  and (_01336_, _01335_, _23037_);
  and (_01338_, _01336_, _01334_);
  not (_01339_, _01338_);
  and (_01340_, _26522_, _26490_);
  not (_01341_, _01340_);
  and (_01342_, _01341_, _26523_);
  and (_01343_, _01342_, _23531_);
  and (_01344_, _01280_, _23606_);
  nand (_01345_, _23558_, _23508_);
  nor (_01346_, _01345_, _23278_);
  and (_01347_, _01346_, _23248_);
  and (_01348_, _01347_, _23217_);
  and (_01349_, _01348_, _23445_);
  and (_01350_, _01349_, _23406_);
  and (_01351_, _01350_, _23121_);
  and (_01352_, _01351_, _23468_);
  nor (_01353_, _01352_, _01344_);
  nor (_01355_, _01353_, _23373_);
  and (_01356_, _01353_, _23373_);
  nor (_01357_, _01356_, _01355_);
  and (_01358_, _01357_, _23543_);
  and (_01359_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  and (_01360_, _23366_, _23330_);
  not (_01361_, _01360_);
  and (_01362_, _23373_, _23468_);
  nor (_01363_, _01362_, _23569_);
  and (_01365_, _01363_, _01361_);
  and (_01366_, _23509_, _23211_);
  and (_01368_, _23494_, _23372_);
  or (_01369_, _01368_, _01366_);
  or (_01370_, _01369_, _01365_);
  nor (_01372_, _01370_, _01359_);
  not (_01373_, _01372_);
  nor (_01374_, _01373_, _01358_);
  not (_01375_, _01374_);
  nor (_01376_, _01375_, _01343_);
  and (_01377_, _01376_, _01339_);
  nor (_01378_, _01377_, _00918_);
  and (_01379_, _00062_, _26604_);
  and (_01380_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01381_, _01380_, _01379_);
  or (_01383_, _01381_, _01378_);
  or (_01384_, _01383_, _01327_);
  or (_01385_, _01384_, _01325_);
  or (_01386_, _01250_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01387_, _01386_, _00879_);
  or (_01388_, _01244_, _01262_);
  or (_01389_, _01388_, _00907_);
  and (_01390_, _01389_, _01387_);
  nand (_01391_, _01390_, _01329_);
  or (_01392_, _01390_, _01329_);
  and (_01393_, _01392_, _01391_);
  and (_01394_, _01393_, _00323_);
  or (_01395_, _01394_, _01385_);
  or (_01396_, _01395_, _00602_);
  or (_01397_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_01398_, _01317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_01399_, _01398_, _01397_);
  or (_01400_, _01399_, _00320_);
  and (_01401_, _01400_, _22761_);
  and (_26899_[14], _01401_, _01396_);
  not (_01402_, _24409_);
  not (_01403_, _24288_);
  and (_01404_, _01403_, _24262_);
  and (_01405_, _01404_, _24311_);
  and (_01406_, _01405_, _01402_);
  and (_01408_, _24363_, _24340_);
  and (_01409_, _01408_, _24385_);
  and (_01410_, _01409_, _01406_);
  nor (_01411_, _01403_, _24262_);
  and (_01412_, _01411_, _24311_);
  and (_01414_, _01412_, _24409_);
  not (_01415_, _01414_);
  and (_01416_, _24363_, _01074_);
  nor (_01417_, _24436_, _00953_);
  and (_01418_, _01417_, _01416_);
  and (_01419_, _01014_, _24340_);
  and (_01420_, _01419_, _00953_);
  and (_01421_, _01420_, _24436_);
  nor (_01422_, _01421_, _01418_);
  nor (_01424_, _01422_, _01415_);
  nor (_01425_, _01424_, _01410_);
  not (_01426_, _01406_);
  and (_01427_, _01416_, _00953_);
  and (_01428_, _01427_, _24436_);
  nor (_01429_, _24363_, _24340_);
  and (_01430_, _01429_, _01417_);
  nor (_01432_, _01430_, _01428_);
  or (_01433_, _01432_, _01426_);
  and (_01434_, _01414_, _00953_);
  nand (_01435_, _01434_, _01408_);
  and (_01436_, _01435_, _01433_);
  and (_01437_, _01428_, _01414_);
  and (_01438_, _24436_, _24385_);
  and (_01439_, _01438_, _01419_);
  and (_01440_, _01405_, _24409_);
  and (_01441_, _01440_, _01439_);
  or (_01442_, _01441_, _01437_);
  and (_01443_, _01409_, _01414_);
  nor (_01444_, _01443_, _01442_);
  and (_01445_, _01416_, _24385_);
  and (_01446_, _01445_, _24436_);
  not (_01447_, _24436_);
  and (_01448_, _01427_, _01447_);
  nor (_01449_, _01448_, _01446_);
  or (_01450_, _01449_, _01426_);
  not (_01451_, _24311_);
  nor (_01452_, _01451_, _24262_);
  and (_01453_, _01452_, _01403_);
  and (_01454_, _01453_, _01402_);
  not (_01455_, _01454_);
  and (_01456_, _01408_, _00953_);
  and (_01457_, _01456_, _24436_);
  nor (_01458_, _01457_, _01439_);
  or (_01459_, _01458_, _01455_);
  and (_01460_, _01459_, _01450_);
  and (_01461_, _01460_, _01444_);
  and (_01462_, _01461_, _01436_);
  and (_01463_, _01462_, _01425_);
  and (_01464_, _01453_, _24409_);
  nor (_01465_, _01430_, _01446_);
  nor (_01466_, _01465_, _01415_);
  nor (_01467_, _01466_, _01464_);
  and (_01468_, _24385_, _01014_);
  and (_01469_, _01468_, _01074_);
  and (_01470_, _01469_, _24436_);
  nor (_01471_, _01421_, _01470_);
  nor (_01472_, _01471_, _01426_);
  nor (_01473_, _01412_, _01406_);
  and (_01474_, _01419_, _01417_);
  nor (_01475_, _24385_, _24363_);
  and (_01476_, _01475_, _01074_);
  and (_01477_, _01476_, _01414_);
  and (_01478_, _01477_, _24436_);
  nor (_01479_, _01478_, _01474_);
  nor (_01480_, _01479_, _01473_);
  nor (_01481_, _01480_, _01472_);
  and (_01482_, _01481_, _01467_);
  nor (_01483_, _01411_, _01404_);
  nor (_01484_, _24436_, _01451_);
  nand (_01485_, _01484_, _01420_);
  or (_01486_, _01485_, _01483_);
  and (_01487_, _01412_, _01402_);
  nand (_01488_, _01446_, _01487_);
  and (_01489_, _01440_, _01474_);
  and (_01490_, _01446_, _01454_);
  nor (_01491_, _01490_, _01489_);
  and (_01492_, _01487_, _01421_);
  and (_01493_, _01454_, _01418_);
  nor (_01495_, _01493_, _01492_);
  and (_01496_, _01495_, _01491_);
  and (_01497_, _01496_, _01488_);
  and (_01498_, _01497_, _01486_);
  and (_01499_, _01498_, _01482_);
  not (_01501_, _01427_);
  and (_01502_, _01471_, _01501_);
  nor (_01503_, _01502_, _24311_);
  and (_01504_, _01420_, _01454_);
  and (_01505_, _01418_, _01406_);
  and (_01506_, _01487_, _01456_);
  or (_01507_, _01506_, _01505_);
  or (_01508_, _01507_, _01504_);
  and (_01509_, _01428_, _01454_);
  and (_01510_, _01474_, _01454_);
  and (_01511_, _01476_, _01447_);
  and (_01512_, _01511_, _01414_);
  or (_01513_, _01512_, _01510_);
  or (_01514_, _01513_, _01509_);
  or (_01515_, _01514_, _01508_);
  nor (_01516_, _01515_, _01503_);
  and (_01517_, _01428_, _01487_);
  not (_01519_, _01517_);
  and (_01521_, _24436_, _00953_);
  nor (_01522_, _01521_, _01417_);
  and (_01524_, _01522_, _01408_);
  and (_01525_, _01524_, _01454_);
  and (_01526_, _01414_, _01470_);
  nor (_01527_, _01526_, _01525_);
  and (_01528_, _01527_, _01519_);
  nor (_01529_, _01448_, _01469_);
  nor (_01530_, _01529_, _01455_);
  not (_01531_, _01439_);
  nor (_01532_, _01473_, _01531_);
  nor (_01533_, _01532_, _01530_);
  and (_01534_, _01533_, _01528_);
  and (_01535_, _24288_, _24262_);
  and (_01536_, _01484_, _01535_);
  nand (_01537_, _01536_, _01416_);
  and (_01538_, _24436_, _24311_);
  and (_01539_, _01538_, _01535_);
  or (_01540_, _01420_, _01427_);
  and (_01541_, _01540_, _01539_);
  and (_01542_, _01418_, _01451_);
  nor (_01543_, _01542_, _01541_);
  and (_01544_, _01543_, _01537_);
  and (_01545_, _01544_, _01534_);
  and (_01546_, _01545_, _01516_);
  and (_01547_, _01546_, _01499_);
  and (_01548_, _01547_, _01463_);
  and (_01549_, _01457_, _01454_);
  and (_01550_, _01420_, _01447_);
  and (_01551_, _01440_, _01550_);
  nor (_01552_, _01551_, _01549_);
  and (_01553_, _01552_, _01491_);
  and (_01554_, _01553_, _01528_);
  nor (_01555_, _01535_, _01451_);
  not (_01556_, _01555_);
  and (_01557_, _01556_, _01428_);
  nor (_01558_, _01557_, _01442_);
  and (_01559_, _01558_, _01425_);
  and (_01560_, _01559_, _01554_);
  not (_01561_, _01560_);
  nor (_01562_, _01561_, _01548_);
  not (_01563_, _01562_);
  and (_01564_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01565_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01567_, _01565_, _01564_);
  and (_01569_, _01567_, _01563_);
  nor (_01570_, _01567_, _01563_);
  nor (_01571_, _01570_, _01569_);
  or (_01572_, _01571_, _25562_);
  not (_01573_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01574_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_01575_, _01574_, _01573_);
  and (_01576_, _01575_, _01572_);
  and (_01577_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_01578_, _01577_, _01576_);
  and (_26900_[0], _01578_, _22761_);
  and (_01579_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01580_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01581_, _01580_, _01579_);
  and (_01583_, _01581_, _01564_);
  nor (_01584_, _01581_, _01564_);
  nor (_01585_, _01584_, _01583_);
  not (_01586_, _01585_);
  nor (_01587_, _01586_, _01548_);
  and (_01588_, _01586_, _01548_);
  nor (_01589_, _01588_, _01587_);
  and (_01590_, _01589_, _01569_);
  nor (_01591_, _01589_, _01569_);
  nor (_01592_, _01591_, _01590_);
  or (_01593_, _01592_, _25562_);
  or (_01594_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01595_, _01594_, _01573_);
  and (_01596_, _01595_, _01593_);
  and (_01597_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_01598_, _01597_, _01596_);
  and (_26900_[1], _01598_, _22761_);
  nor (_01599_, _01590_, _01587_);
  not (_01600_, _01599_);
  nor (_01601_, _01583_, _01579_);
  and (_01602_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01603_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01604_, _01603_, _01602_);
  not (_01605_, _01604_);
  nor (_01606_, _01605_, _01601_);
  and (_01607_, _01605_, _01601_);
  nor (_01608_, _01607_, _01606_);
  and (_01609_, _01608_, _01600_);
  nor (_01610_, _01608_, _01600_);
  nor (_01611_, _01610_, _01609_);
  or (_01612_, _01611_, _25562_);
  or (_01613_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01614_, _01613_, _01573_);
  and (_01615_, _01614_, _01612_);
  and (_01616_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01617_, _01616_, _01615_);
  and (_26900_[2], _01617_, _22761_);
  nor (_01619_, _01606_, _01602_);
  nor (_01620_, _01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01621_, _01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_01622_, _01621_, _01620_);
  not (_01623_, _01622_);
  and (_01624_, _01623_, _01609_);
  nor (_01625_, _01623_, _01609_);
  nor (_01626_, _01625_, _01624_);
  or (_01627_, _01626_, _25562_);
  or (_01628_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01629_, _01628_, _01573_);
  and (_01630_, _01629_, _01627_);
  and (_01631_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01632_, _01631_, _01630_);
  and (_26900_[3], _01632_, _22761_);
  and (_01634_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_01635_, _01143_, _01634_);
  nand (_01636_, _01635_, _01620_);
  or (_01637_, _01635_, _01620_);
  and (_01638_, _01637_, _01636_);
  and (_01639_, _01638_, _01624_);
  nor (_01640_, _01638_, _01624_);
  nor (_01641_, _01640_, _01639_);
  or (_01642_, _01641_, _25562_);
  or (_01643_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01644_, _01643_, _01573_);
  and (_01645_, _01644_, _01642_);
  and (_01646_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01647_, _01646_, _01645_);
  and (_26900_[4], _01647_, _22761_);
  and (_01648_, _01619_, _01144_);
  and (_01649_, _01619_, _01143_);
  nor (_01650_, _01649_, _01142_);
  nor (_01651_, _01650_, _01648_);
  not (_01652_, _01651_);
  and (_01653_, _01652_, _01639_);
  nor (_01654_, _01652_, _01639_);
  nor (_01655_, _01654_, _01653_);
  or (_01656_, _01655_, _25562_);
  or (_01657_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01658_, _01657_, _01573_);
  and (_01660_, _01658_, _01656_);
  and (_01661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01662_, _01661_, _01660_);
  and (_26900_[5], _01662_, _22761_);
  not (_01663_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_01664_, _01648_, _01663_);
  and (_01665_, _01144_, _01663_);
  and (_01666_, _01665_, _01619_);
  nor (_01667_, _01666_, _01664_);
  not (_01668_, _01667_);
  and (_01669_, _01668_, _01653_);
  nor (_01670_, _01668_, _01653_);
  nor (_01671_, _01670_, _01669_);
  or (_01672_, _01671_, _25562_);
  or (_01673_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01674_, _01673_, _01573_);
  and (_01675_, _01674_, _01672_);
  and (_01676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01678_, _01676_, _01675_);
  and (_26900_[6], _01678_, _22761_);
  not (_01679_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_01680_, _01665_, _01679_);
  and (_01681_, _01680_, _01619_);
  nor (_01682_, _01666_, _01679_);
  nor (_01683_, _01682_, _01681_);
  not (_01685_, _01683_);
  and (_01686_, _01685_, _01669_);
  nor (_01687_, _01685_, _01669_);
  nor (_01688_, _01687_, _01686_);
  or (_01689_, _01688_, _25562_);
  or (_01691_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01692_, _01691_, _01573_);
  and (_01693_, _01692_, _01689_);
  and (_01694_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_01695_, _01694_, _01693_);
  and (_26900_[7], _01695_, _22761_);
  nor (_01696_, _01681_, _01148_);
  and (_01697_, _01680_, _01148_);
  and (_01698_, _01697_, _01619_);
  nor (_01699_, _01698_, _01696_);
  not (_01700_, _01699_);
  and (_01701_, _01700_, _01686_);
  nor (_01702_, _01700_, _01686_);
  nor (_01703_, _01702_, _01701_);
  or (_01704_, _01703_, _25562_);
  or (_01705_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01706_, _01705_, _01573_);
  and (_01707_, _01706_, _01704_);
  and (_01708_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01709_, _01708_, _01707_);
  and (_26900_[8], _01709_, _22761_);
  not (_01710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01712_, _01697_, _01710_);
  and (_01713_, _01712_, _01619_);
  nor (_01714_, _01698_, _01710_);
  nor (_01715_, _01714_, _01713_);
  not (_01716_, _01715_);
  and (_01717_, _01716_, _01701_);
  or (_01719_, _01716_, _01701_);
  nand (_01720_, _01719_, _25561_);
  nor (_01721_, _01720_, _01717_);
  nor (_01722_, _25561_, _00967_);
  or (_01723_, _01722_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01724_, _01723_, _01721_);
  or (_01725_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _01573_);
  and (_01726_, _01725_, _22761_);
  and (_26900_[9], _01726_, _01724_);
  not (_01727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01728_, _01713_, _01727_);
  and (_01729_, _01712_, _01727_);
  and (_01730_, _01729_, _01619_);
  nor (_01732_, _01730_, _01728_);
  not (_01733_, _01732_);
  and (_01734_, _01733_, _01717_);
  nor (_01735_, _01733_, _01717_);
  nor (_01736_, _01735_, _01734_);
  or (_01737_, _01736_, _25562_);
  or (_01738_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01739_, _01738_, _01573_);
  and (_01740_, _01739_, _01737_);
  and (_01741_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01742_, _01741_, _01740_);
  and (_26900_[10], _01742_, _22761_);
  and (_01743_, _01730_, _01141_);
  nor (_01744_, _01730_, _01141_);
  nor (_01745_, _01744_, _01743_);
  not (_01746_, _01745_);
  and (_01747_, _01746_, _01734_);
  nor (_01748_, _01746_, _01734_);
  nor (_01749_, _01748_, _01747_);
  or (_01750_, _01749_, _25562_);
  or (_01751_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01752_, _01751_, _01573_);
  and (_01753_, _01752_, _01750_);
  and (_01754_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01755_, _01754_, _01753_);
  and (_26900_[11], _01755_, _22761_);
  nor (_01756_, _01743_, _01188_);
  and (_01757_, _01729_, _01141_);
  and (_01759_, _01757_, _01188_);
  and (_01760_, _01759_, _01619_);
  nor (_01761_, _01760_, _01756_);
  not (_01762_, _01761_);
  and (_01763_, _01762_, _01747_);
  nor (_01764_, _01762_, _01747_);
  nor (_01765_, _01764_, _01763_);
  or (_01766_, _01765_, _25562_);
  or (_01767_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01768_, _01767_, _01573_);
  and (_01769_, _01768_, _01766_);
  and (_01770_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01771_, _01770_, _01769_);
  and (_26900_[12], _01771_, _22761_);
  nor (_01772_, _01760_, _01303_);
  and (_01773_, _01759_, _01303_);
  and (_01774_, _01773_, _01619_);
  nor (_01775_, _01774_, _01772_);
  not (_01776_, _01775_);
  and (_01777_, _01776_, _01763_);
  nor (_01778_, _01776_, _01763_);
  nor (_01780_, _01778_, _01777_);
  or (_01781_, _01780_, _25562_);
  or (_01782_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01783_, _01782_, _01573_);
  and (_01784_, _01783_, _01781_);
  and (_01785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01786_, _01785_, _01784_);
  and (_26900_[13], _01786_, _22761_);
  nor (_01787_, _01774_, _01321_);
  and (_01788_, _01774_, _01321_);
  nor (_01789_, _01788_, _01787_);
  not (_01790_, _01789_);
  and (_01791_, _01790_, _01777_);
  nor (_01792_, _01790_, _01777_);
  nor (_01793_, _01792_, _01791_);
  or (_01794_, _01793_, _25562_);
  or (_01795_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01796_, _01795_, _01573_);
  and (_01797_, _01796_, _01794_);
  and (_01798_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01799_, _01798_, _01797_);
  and (_26900_[14], _01799_, _22761_);
  nand (_01800_, _23597_, _22933_);
  and (_01801_, _01800_, _23023_);
  and (_01802_, _01801_, _23017_);
  and (_01803_, _01802_, _23838_);
  not (_01804_, _01802_);
  and (_01805_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_22623_, _01805_, _01803_);
  and (_01806_, _01802_, _23718_);
  and (_01807_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_22624_, _01807_, _01806_);
  nor (_01808_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_01809_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_01810_, _01809_, _01808_);
  not (_01811_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_01812_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_01813_, _01812_, _01811_);
  and (_01814_, _01813_, _01810_);
  and (_01815_, _01814_, _25108_);
  and (_01816_, _01815_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01817_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_26904_[0], _01817_, _22761_);
  and (_01819_, _01815_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01820_, _01819_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_26904_[1], _01820_, _22761_);
  and (_01821_, _01815_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_01822_, _01821_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_26904_[2], _01822_, _22761_);
  and (_01823_, _01814_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_01824_, _01823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_26904_[3], _01824_, _22761_);
  and (_01825_, _01815_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01826_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_26904_[4], _01826_, _22761_);
  and (_01827_, _01815_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_01828_, _01827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_26904_[5], _01828_, _22761_);
  and (_01829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22761_);
  and (_01830_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _22761_);
  and (_01831_, _01830_, _01815_);
  or (_26904_[6], _01831_, _01829_);
  nor (_01832_, _01562_, _25566_);
  nand (_01833_, _01832_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01834_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or (_01835_, _01832_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_01836_, _01835_, _01834_);
  and (_26905_[0], _01836_, _01833_);
  and (_01837_, _01563_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01838_, _01548_, _24247_);
  and (_01839_, _01548_, _24247_);
  nor (_01840_, _01839_, _01838_);
  and (_01841_, _01840_, _01837_);
  nor (_01842_, _01840_, _01837_);
  nor (_01843_, _01842_, _01841_);
  or (_01844_, _01843_, _25566_);
  or (_01845_, _22768_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01846_, _01845_, _01834_);
  and (_26905_[1], _01846_, _01844_);
  and (_01847_, _24567_, _23838_);
  and (_01848_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or (_22625_, _01848_, _01847_);
  nor (_26906_[5], _00727_, rst);
  and (_01849_, _01802_, _23589_);
  and (_01850_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_22626_, _01850_, _01849_);
  nor (_26906_[1], _00430_, rst);
  and (_01851_, _01802_, _23755_);
  and (_01852_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_22627_, _01852_, _01851_);
  not (_01853_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_01854_, _01853_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_01855_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_01857_, _01855_, _01854_);
  and (_26908_[0], _01857_, _22761_);
  and (_01858_, _01853_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_01859_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01860_, _01859_, _01858_);
  and (_26908_[1], _01860_, _22761_);
  and (_01861_, _01853_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_01862_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01863_, _01862_, _01861_);
  and (_26908_[2], _01863_, _22761_);
  and (_01864_, _01853_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_01865_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01866_, _01865_, _01864_);
  and (_26908_[3], _01866_, _22761_);
  and (_01867_, _01853_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_01868_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01869_, _01868_, _01867_);
  and (_26908_[4], _01869_, _22761_);
  and (_01870_, _01853_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_01871_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01872_, _01871_, _01870_);
  and (_26908_[5], _01872_, _22761_);
  and (_01873_, _01853_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_01874_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01875_, _01874_, _01873_);
  and (_26908_[6], _01875_, _22761_);
  and (_01876_, _01802_, _23635_);
  and (_01877_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_22628_, _01877_, _01876_);
  not (_01879_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01880_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor (_01881_, _01880_, _01879_);
  and (_01882_, _01880_, _01879_);
  nor (_01883_, _01882_, _01881_);
  and (_26911_[0], _01883_, _22761_);
  nor (_01884_, _01881_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01885_, _01881_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01886_, _01885_, _01884_);
  nor (_26911_[1], _01886_, rst);
  and (_01887_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01888_, _01887_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01889_, _01887_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01890_, _01889_, _01888_);
  or (_01891_, _01890_, _01880_);
  and (_26911_[2], _01891_, _22761_);
  and (_01892_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_01893_, _25781_, _25783_);
  or (_01894_, _01893_, _01892_);
  and (_26913_[0], _01894_, _22761_);
  and (_01895_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_01896_, _25781_, _25787_);
  or (_01897_, _01896_, _01895_);
  and (_26913_[1], _01897_, _22761_);
  and (_01898_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_01899_, _25781_, _25791_);
  or (_01900_, _01899_, _01898_);
  and (_26913_[2], _01900_, _22761_);
  and (_01901_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_01902_, _25781_, _25795_);
  or (_01903_, _01902_, _01901_);
  and (_26913_[3], _01903_, _22761_);
  and (_01904_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_01905_, _25781_, _25799_);
  or (_01906_, _01905_, _01904_);
  and (_26913_[4], _01906_, _22761_);
  and (_01907_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_01908_, _25781_, _25803_);
  or (_01909_, _01908_, _01907_);
  and (_26913_[5], _01909_, _22761_);
  and (_01910_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_01911_, _25781_, _25807_);
  or (_01912_, _01911_, _01910_);
  and (_26913_[6], _01912_, _22761_);
  and (_01913_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_01914_, _25781_, _25811_);
  or (_01915_, _01914_, _01913_);
  and (_26913_[7], _01915_, _22761_);
  and (_01916_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_01917_, _25781_, _25815_);
  or (_01919_, _01917_, _01916_);
  and (_26913_[8], _01919_, _22761_);
  and (_01920_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_01921_, _25781_, _25820_);
  or (_01922_, _01921_, _01920_);
  and (_26913_[9], _01922_, _22761_);
  and (_01923_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_01924_, _25781_, _25824_);
  or (_01925_, _01924_, _01923_);
  and (_26913_[10], _01925_, _22761_);
  and (_01926_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_01927_, _25781_, _25828_);
  or (_01928_, _01927_, _01926_);
  and (_26913_[11], _01928_, _22761_);
  and (_01929_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_01930_, _25781_, _25833_);
  or (_01931_, _01930_, _01929_);
  and (_26913_[12], _01931_, _22761_);
  and (_01932_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_01933_, _25781_, _25837_);
  or (_01934_, _01933_, _01932_);
  and (_26913_[13], _01934_, _22761_);
  and (_01935_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_01936_, _25781_, _25841_);
  or (_01937_, _01936_, _01935_);
  and (_26913_[14], _01937_, _22761_);
  or (_01938_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_01939_, _25845_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_01940_, _01939_, _22761_);
  and (_26913_[15], _01940_, _01938_);
  and (_01941_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01942_, _25781_, _25849_);
  or (_01943_, _01942_, _01941_);
  and (_26913_[16], _01943_, _22761_);
  and (_01944_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01945_, _25781_, _25855_);
  or (_01946_, _01945_, _01944_);
  and (_26913_[17], _01946_, _22761_);
  and (_01947_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01948_, _25781_, _25859_);
  or (_01949_, _01948_, _01947_);
  and (_26913_[18], _01949_, _22761_);
  and (_01950_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01951_, _25781_, _25863_);
  or (_01952_, _01951_, _01950_);
  and (_26913_[19], _01952_, _22761_);
  and (_01953_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01954_, _25781_, _25867_);
  or (_01955_, _01954_, _01953_);
  and (_26913_[20], _01955_, _22761_);
  and (_01956_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01957_, _25781_, _25871_);
  or (_01958_, _01957_, _01956_);
  and (_26913_[21], _01958_, _22761_);
  and (_01959_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01960_, _25781_, _25875_);
  or (_01961_, _01960_, _01959_);
  and (_26913_[22], _01961_, _22761_);
  or (_01962_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_01963_, _25845_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_01964_, _01963_, _22761_);
  and (_26913_[23], _01964_, _01962_);
  and (_01965_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01966_, _25781_, _25882_);
  or (_01967_, _01966_, _01965_);
  and (_26913_[24], _01967_, _22761_);
  and (_01968_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01969_, _25781_, _25888_);
  or (_01970_, _01969_, _01968_);
  and (_26913_[25], _01970_, _22761_);
  and (_01971_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01972_, _25781_, _25892_);
  or (_01973_, _01972_, _01971_);
  and (_26913_[26], _01973_, _22761_);
  and (_01974_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_01975_, _25845_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_01976_, _01975_, _01974_);
  and (_26913_[27], _01976_, _22761_);
  and (_01977_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_01978_, _25845_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_01979_, _01978_, _01977_);
  and (_26913_[28], _01979_, _22761_);
  and (_01980_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01981_, _25781_, _25903_);
  or (_01982_, _01981_, _01980_);
  and (_26913_[29], _01982_, _22761_);
  and (_01983_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01984_, _25781_, _25907_);
  or (_01985_, _01984_, _01983_);
  and (_26913_[30], _01985_, _22761_);
  and (_26870_[1], _26748_, _22761_);
  nor (_26896_[3], _00090_, rst);
  and (_01986_, _23843_, _23791_);
  and (_01987_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or (_22629_, _01987_, _01986_);
  and (_01988_, _24420_, _24459_);
  nor (_01989_, _24389_, _24368_);
  and (_01990_, _01989_, _24474_);
  and (_01991_, _01990_, _24346_);
  or (_01992_, _01991_, _26664_);
  or (_01993_, _26658_, _24480_);
  or (_01994_, _01993_, _01992_);
  or (_01995_, _01994_, _01988_);
  and (_01996_, _01989_, _24458_);
  and (_01997_, _24515_, _24317_);
  or (_01999_, _01997_, _01996_);
  or (_02000_, _01999_, _26697_);
  or (_02001_, _02000_, _24519_);
  and (_02002_, _24518_, _24489_);
  or (_02003_, _02002_, _26711_);
  or (_02004_, _02003_, _02001_);
  and (_02005_, _24491_, _24443_);
  and (_02006_, _02005_, _24486_);
  or (_02007_, _26694_, _02006_);
  nor (_02008_, _26729_, _24508_);
  not (_02009_, _02008_);
  or (_02010_, _02009_, _02007_);
  or (_02011_, _02010_, _02004_);
  or (_02012_, _02011_, _01995_);
  and (_02013_, _02012_, _22768_);
  and (_02014_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02015_, _02014_, _26822_);
  or (_02016_, _02015_, _02013_);
  and (_26880_[2], _02016_, _22761_);
  and (_02017_, _24558_, _23854_);
  not (_02018_, _02017_);
  and (_02019_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_02020_, _02017_, _23589_);
  or (_22630_, _02020_, _02019_);
  and (_02021_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_02022_, _02017_, _23755_);
  or (_22631_, _02022_, _02021_);
  and (_02023_, _24492_, _24486_);
  or (_02024_, _26596_, _02023_);
  and (_02025_, _24515_, _24321_);
  or (_02026_, _02025_, _26594_);
  or (_02027_, _02026_, _02009_);
  or (_02028_, _02027_, _02024_);
  and (_02029_, _00271_, _24470_);
  and (_02030_, _26664_, _24445_);
  or (_02031_, _02030_, _01991_);
  or (_02032_, _02031_, _02029_);
  or (_02033_, _26680_, _24507_);
  or (_02034_, _02033_, _26657_);
  and (_02035_, _24517_, _24466_);
  or (_02036_, _01993_, _02035_);
  or (_02037_, _02036_, _02034_);
  and (_02038_, _26692_, _24321_);
  or (_02039_, _02038_, _01999_);
  nor (_02040_, _24417_, _26587_);
  and (_02041_, _26595_, _24317_);
  or (_02042_, _02041_, _02040_);
  or (_02043_, _02042_, _02039_);
  or (_02044_, _02043_, _02007_);
  or (_02045_, _02044_, _02037_);
  or (_02046_, _02045_, _02032_);
  or (_02047_, _02046_, _02028_);
  and (_02048_, _02047_, _22768_);
  and (_02049_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02050_, _02049_, _26820_);
  or (_02052_, _02050_, _02048_);
  and (_26880_[1], _02052_, _22761_);
  nor (_02053_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_02054_, _02053_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not (_02055_, _02054_);
  or (_02056_, _02055_, _26568_);
  or (_02057_, _02054_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02058_, _02057_, _22761_);
  and (_26917_[0], _02058_, _02056_);
  or (_02059_, _02055_, _00408_);
  or (_02060_, _02054_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02061_, _02060_, _22761_);
  and (_26917_[1], _02061_, _02059_);
  or (_02062_, _02055_, _00484_);
  or (_02063_, _02054_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_02064_, _02063_, _22761_);
  and (_26917_[2], _02064_, _02062_);
  or (_02065_, _02055_, _00580_);
  or (_02066_, _02054_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_02067_, _02066_, _22761_);
  and (_26917_[3], _02067_, _02065_);
  and (_02069_, _23854_, _23599_);
  and (_02070_, _02069_, _23791_);
  not (_02071_, _02069_);
  and (_02072_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_22632_, _02072_, _02070_);
  and (_02073_, _25666_, _23926_);
  nand (_02074_, _02073_, _23585_);
  and (_02075_, _25702_, _25696_);
  not (_02076_, _02075_);
  and (_02077_, _25666_, _23993_);
  nor (_02078_, _02077_, _02076_);
  or (_02079_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_02080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_02081_, _02078_, _02080_);
  and (_02082_, _02081_, _02079_);
  or (_02083_, _02082_, _02073_);
  and (_02084_, _02083_, _22761_);
  and (_22633_, _02084_, _02074_);
  and (_22634_, t2ex_i, _22761_);
  and (_02086_, _24647_, _23875_);
  or (_02087_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_02088_, _02087_, _22761_);
  not (_02089_, _02086_);
  or (_02090_, _02089_, _23709_);
  and (_22635_, _02090_, _02088_);
  nand (_02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _22761_);
  nor (_22636_, _02091_, t2ex_i);
  and (_02092_, _01801_, _23849_);
  and (_02093_, _02092_, _23755_);
  not (_02095_, _02092_);
  and (_02096_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_27025_, _02096_, _02093_);
  nor (_02097_, t2_i, rst);
  and (_22637_, _02097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nor (_02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_02099_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _22761_);
  and (_02101_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_22638_, _02101_, _02099_);
  and (_02102_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_02103_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_22639_, _02103_, _02102_);
  and (_02104_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02105_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_22640_, _02105_, _02104_);
  and (_22641_, t2_i, _22761_);
  nor (_26869_[3], _24311_, rst);
  and (_02106_, _24080_, _23718_);
  and (_02107_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_22642_, _02107_, _02106_);
  and (_02108_, _02092_, _23635_);
  and (_02109_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_22643_, _02109_, _02108_);
  and (_02110_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_02111_, _25619_, _23676_);
  or (_22644_, _02111_, _02110_);
  and (_02112_, _02092_, _23589_);
  and (_02113_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_22645_, _02113_, _02112_);
  and (_22646_, _01829_, _24847_);
  and (_02114_, _24847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_02115_, _02114_, _24935_);
  and (_22647_, _02115_, _22761_);
  and (_02116_, _24881_, _24938_);
  and (_02117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _24850_);
  and (_02118_, _02117_, _24867_);
  or (_02119_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02120_, _02119_, _24873_);
  and (_02121_, _02120_, _24868_);
  or (_02122_, _25003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02123_, _02122_, _25006_);
  nand (_02124_, _02117_, _24876_);
  nand (_02125_, _02124_, _24873_);
  or (_02126_, _02125_, _02123_);
  and (_02127_, _02126_, _02121_);
  or (_02128_, _02127_, _02118_);
  and (_02129_, _02128_, _02116_);
  not (_02130_, _24903_);
  or (_02131_, _02130_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_02132_, _02119_, _24900_);
  and (_02133_, _02132_, _24895_);
  or (_02134_, _25020_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02135_, _02134_, _25019_);
  nand (_02137_, _02117_, _24889_);
  nand (_02138_, _02137_, _24900_);
  or (_02139_, _02138_, _02135_);
  and (_02140_, _02139_, _02133_);
  and (_02141_, _02117_, _24894_);
  or (_02142_, _02141_, _24903_);
  or (_02143_, _02142_, _02140_);
  and (_02144_, _02143_, _24933_);
  or (_02145_, _02144_, _24847_);
  and (_02146_, _02145_, _02131_);
  or (_02147_, _02146_, _02129_);
  and (_22648_, _02147_, _22761_);
  and (_02148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_02149_, _02148_, _24867_);
  or (_02150_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _24850_);
  or (_02151_, _02150_, _24873_);
  and (_02152_, _02151_, _24868_);
  or (_02154_, _24942_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02155_, _02154_, _24940_);
  nand (_02156_, _02148_, _24876_);
  nand (_02157_, _02156_, _24873_);
  or (_02158_, _02157_, _02155_);
  and (_02159_, _02158_, _02152_);
  or (_02160_, _02159_, _02149_);
  and (_02161_, _02160_, _02116_);
  or (_02162_, _02130_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_02163_, _02150_, _24900_);
  and (_02164_, _02163_, _24895_);
  or (_02165_, _24964_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02166_, _02165_, _24963_);
  nand (_02167_, _02148_, _24889_);
  nand (_02168_, _02167_, _24900_);
  or (_02169_, _02168_, _02166_);
  and (_02170_, _02169_, _02164_);
  and (_02171_, _02148_, _24894_);
  or (_02172_, _02171_, _24903_);
  or (_02173_, _02172_, _02170_);
  and (_02174_, _02173_, _24933_);
  or (_02175_, _02174_, _24847_);
  and (_02176_, _02175_, _02162_);
  or (_02177_, _02176_, _02161_);
  and (_22649_, _02177_, _22761_);
  and (_02178_, _24708_, _23919_);
  or (_02179_, _02178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_02180_, _02179_, _24716_);
  nand (_02181_, _02178_, _23522_);
  and (_02182_, _02181_, _02180_);
  nor (_02183_, _24716_, _23628_);
  or (_02184_, _02183_, _02182_);
  and (_22650_, _02184_, _22761_);
  and (_02185_, _24732_, _24634_);
  not (_02186_, _24634_);
  or (_02187_, _24728_, _02186_);
  or (_02188_, _02187_, _24641_);
  and (_02189_, _02188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_02190_, _02189_, _24674_);
  or (_02191_, _02190_, _02185_);
  nand (_02192_, _24648_, _23914_);
  and (_02193_, _02192_, _22761_);
  and (_22651_, _02193_, _02191_);
  and (_02194_, _23838_, _23798_);
  and (_02195_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or (_22652_, _02195_, _02194_);
  and (_02196_, _01802_, _23676_);
  and (_02197_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_22653_, _02197_, _02196_);
  and (_02198_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_02199_, _02017_, _23791_);
  or (_22654_, _02199_, _02198_);
  and (_02200_, _01801_, _23803_);
  and (_02201_, _02200_, _23589_);
  not (_02202_, _02200_);
  and (_02203_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_22655_, _02203_, _02201_);
  and (_02204_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_02205_, _02017_, _23718_);
  or (_22656_, _02205_, _02204_);
  and (_02206_, _02200_, _23755_);
  and (_02207_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_22657_, _02207_, _02206_);
  and (_02208_, _02200_, _23635_);
  and (_02209_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_22658_, _02209_, _02208_);
  and (_02210_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_02211_, _02017_, _23676_);
  or (_22659_, _02211_, _02210_);
  and (_02212_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_02213_, _02017_, _23982_);
  or (_22660_, _02213_, _02212_);
  and (_02214_, _02092_, _23791_);
  and (_02215_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_27024_, _02215_, _02214_);
  and (_02216_, _02092_, _23676_);
  and (_02217_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_22661_, _02217_, _02216_);
  and (_02218_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_02220_, _02017_, _23838_);
  or (_22662_, _02220_, _02218_);
  and (_02221_, _01801_, _23842_);
  and (_02222_, _02221_, _23589_);
  not (_02223_, _02221_);
  and (_02224_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_22663_, _02224_, _02222_);
  and (_02225_, _24541_, _23643_);
  and (_02226_, _02225_, _23838_);
  not (_02227_, _02225_);
  and (_02228_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_22664_, _02228_, _02226_);
  and (_02229_, _25536_, _23718_);
  and (_02230_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_22665_, _02230_, _02229_);
  and (_02231_, _02200_, _23676_);
  and (_02232_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_22666_, _02232_, _02231_);
  and (_02233_, _24558_, _23797_);
  not (_02234_, _02233_);
  and (_02235_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and (_02236_, _02233_, _23635_);
  or (_22667_, _02236_, _02235_);
  and (_02237_, _24768_, _24572_);
  and (_02238_, _02237_, _23838_);
  not (_02239_, _02237_);
  and (_02240_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_22668_, _02240_, _02238_);
  and (_02241_, _01988_, _24443_);
  and (_02242_, _26588_, _24321_);
  and (_02243_, _24418_, _26591_);
  or (_02244_, _02038_, _26572_);
  or (_02245_, _02244_, _02243_);
  or (_02246_, _02245_, _02242_);
  or (_02247_, _02246_, _02241_);
  or (_02248_, _26729_, _02035_);
  and (_02249_, _24517_, _24486_);
  and (_02250_, _24468_, _01989_);
  or (_02251_, _02250_, _02249_);
  or (_02252_, _02251_, _02248_);
  or (_02253_, _24536_, _01990_);
  or (_02254_, _24463_, _24449_);
  or (_02255_, _02254_, _02253_);
  or (_02256_, _26653_, _26688_);
  or (_02257_, _02256_, _02255_);
  or (_02259_, _02257_, _02252_);
  and (_02260_, _24499_, _24486_);
  not (_02261_, _26686_);
  or (_02262_, _02261_, _02260_);
  or (_02263_, _02262_, _26681_);
  and (_02264_, _26591_, _24321_);
  or (_02265_, _24508_, _02264_);
  or (_02266_, _02265_, _02263_);
  or (_02267_, _02266_, _02259_);
  or (_02268_, _02267_, _02247_);
  and (_02269_, _02268_, _22768_);
  and (_02271_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_02272_, _02271_, _26820_);
  or (_02273_, _02272_, _02269_);
  and (_26880_[0], _02273_, _22761_);
  and (_02274_, _02237_, _23791_);
  and (_02275_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_27156_, _02275_, _02274_);
  and (_02276_, _24571_, _23595_);
  and (_02277_, _02276_, _24768_);
  and (_02278_, _02277_, _23982_);
  not (_02279_, _02277_);
  and (_02280_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  or (_22669_, _02280_, _02278_);
  and (_02281_, _25742_, _23718_);
  and (_02282_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or (_22670_, _02282_, _02281_);
  and (_02283_, _02237_, _23676_);
  and (_02284_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_22671_, _02284_, _02283_);
  and (_02285_, _25742_, _23838_);
  and (_02286_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_22672_, _02286_, _02285_);
  and (_02287_, _25742_, _23982_);
  and (_02288_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or (_22673_, _02288_, _02287_);
  and (_02289_, _24572_, _24541_);
  and (_02290_, _02289_, _23755_);
  not (_02291_, _02289_);
  and (_02292_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or (_22674_, _02292_, _02290_);
  and (_02293_, _02289_, _23982_);
  and (_02294_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or (_22675_, _02294_, _02293_);
  and (_02295_, _02289_, _23718_);
  and (_02296_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or (_22676_, _02296_, _02295_);
  nand (_02297_, _23921_, _23748_);
  not (_02298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02299_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_02300_, _02299_, _24182_);
  and (_02301_, _24193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_02302_, _02301_, _23944_);
  and (_02303_, _23938_, _24146_);
  nand (_02304_, _02303_, _02302_);
  and (_02305_, _02304_, _24182_);
  nor (_02306_, _02305_, _02300_);
  and (_02307_, _02306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_02308_, _02307_, _02298_);
  and (_02309_, _02307_, _02298_);
  or (_02310_, _02309_, _02308_);
  or (_02311_, _02310_, _23921_);
  and (_02312_, _02311_, _23928_);
  and (_02313_, _02312_, _02297_);
  and (_02314_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_02315_, _02314_, _02313_);
  and (_22677_, _02315_, _22761_);
  and (_02316_, _02289_, _23791_);
  and (_02317_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or (_22678_, _02317_, _02316_);
  and (_02318_, _24572_, _24117_);
  and (_02319_, _02318_, _23755_);
  not (_02320_, _02318_);
  and (_02321_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_22679_, _02321_, _02319_);
  and (_02322_, _24768_, _24118_);
  and (_02323_, _02322_, _23589_);
  not (_02324_, _02322_);
  and (_02325_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_22680_, _02325_, _02323_);
  and (_02326_, _23641_, _23028_);
  and (_02327_, _02326_, _23982_);
  not (_02328_, _02326_);
  and (_02329_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_22681_, _02329_, _02327_);
  and (_02330_, _02326_, _23635_);
  and (_02331_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or (_27272_, _02331_, _02330_);
  and (_02332_, _02326_, _23755_);
  and (_02333_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or (_22682_, _02333_, _02332_);
  and (_02334_, _02318_, _23635_);
  and (_02335_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_22683_, _02335_, _02334_);
  and (_02336_, _02318_, _23838_);
  and (_02337_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_22684_, _02337_, _02336_);
  and (_02338_, _02318_, _23791_);
  and (_02339_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_22685_, _02339_, _02338_);
  and (_02340_, _02200_, _23838_);
  and (_02341_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_22686_, _02341_, _02340_);
  and (_02342_, _24572_, _23797_);
  and (_02343_, _02342_, _23589_);
  not (_02344_, _02342_);
  and (_02345_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_22687_, _02345_, _02343_);
  and (_02346_, _02200_, _23718_);
  and (_02347_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_22688_, _02347_, _02346_);
  and (_02348_, _02225_, _23635_);
  and (_02349_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_22689_, _02349_, _02348_);
  and (_02350_, _02200_, _23791_);
  and (_02351_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_22690_, _02351_, _02350_);
  or (_02352_, _02306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_02353_, _02307_, _23921_);
  and (_02354_, _02353_, _02352_);
  nor (_02355_, _23922_, _23628_);
  or (_02356_, _02355_, _02354_);
  and (_02357_, _02356_, _23928_);
  and (_02358_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_02359_, _02358_, _02357_);
  and (_22691_, _02359_, _22761_);
  nand (_02360_, _24385_, _22767_);
  or (_02361_, _22767_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_02362_, _02361_, _22761_);
  and (_26873_[5], _02362_, _02360_);
  not (_02363_, _22767_);
  or (_02364_, _24436_, _02363_);
  or (_02365_, _22767_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_02366_, _02365_, _22761_);
  and (_26873_[4], _02366_, _02364_);
  and (_26870_[0], _26674_, _22761_);
  or (_02367_, _24262_, _02363_);
  or (_02368_, _22767_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_02369_, _02368_, _22761_);
  and (_26873_[1], _02369_, _02367_);
  or (_26871_[0], _25616_, _24537_);
  and (_02370_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  and (_02371_, _02233_, _23589_);
  or (_22692_, _02371_, _02370_);
  and (_02372_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and (_02373_, _02233_, _23755_);
  or (_22693_, _02373_, _02372_);
  nor (_02374_, _23531_, _26382_);
  and (_02375_, _26387_, _23531_);
  or (_02376_, _02375_, _02374_);
  and (_22694_, _02376_, _22761_);
  and (_02377_, _23798_, _23718_);
  and (_02378_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or (_22695_, _02378_, _02377_);
  and (_02379_, _24118_, _23797_);
  and (_02380_, _02379_, _23676_);
  not (_02381_, _02379_);
  and (_02382_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_27229_, _02382_, _02380_);
  and (_02383_, _24572_, _23641_);
  and (_02384_, _02383_, _23589_);
  not (_02385_, _02383_);
  and (_02386_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or (_22696_, _02386_, _02384_);
  and (_02387_, _02221_, _23718_);
  and (_02388_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_26990_, _02388_, _02387_);
  and (_02389_, _02221_, _23791_);
  and (_02390_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_26989_, _02390_, _02389_);
  and (_02391_, _02225_, _23676_);
  and (_02392_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_22697_, _02392_, _02391_);
  nand (_02393_, _24340_, _22767_);
  or (_02394_, _22767_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_02395_, _02394_, _22761_);
  and (_26873_[7], _02395_, _02393_);
  and (_02396_, _02383_, _23755_);
  and (_02397_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or (_22698_, _02397_, _02396_);
  and (_02398_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and (_02399_, _02233_, _23791_);
  or (_22699_, _02399_, _02398_);
  and (_02400_, _02221_, _23635_);
  and (_02401_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_22700_, _02401_, _02400_);
  and (_02402_, _02221_, _23982_);
  and (_02403_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_22701_, _02403_, _02402_);
  and (_02404_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_02405_, _02233_, _23676_);
  or (_27063_, _02405_, _02404_);
  and (_02407_, _02221_, _23838_);
  and (_02408_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_26991_, _02408_, _02407_);
  nand (_02409_, _23921_, _23585_);
  and (_02410_, _02299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_02411_, _02410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_02412_, _02411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02413_, _02411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_02414_, _02413_, _02412_);
  and (_02415_, _02414_, _24147_);
  and (_02416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02418_, _02302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_02419_, _02418_, _23938_);
  and (_02420_, _02419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_02421_, _02420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02422_, _02420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_02423_, _02422_, _24192_);
  and (_02424_, _02423_, _02421_);
  or (_02425_, _02424_, _02416_);
  or (_02426_, _02425_, _02415_);
  or (_02427_, _02426_, _23921_);
  and (_02428_, _02427_, _23928_);
  and (_02429_, _02428_, _02409_);
  and (_02430_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02431_, _02430_, _02429_);
  and (_22702_, _02431_, _22761_);
  and (_02432_, _02383_, _23982_);
  and (_02434_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or (_22703_, _02434_, _02432_);
  and (_02436_, _23803_, _23643_);
  and (_02437_, _02436_, _23838_);
  not (_02438_, _02436_);
  and (_02439_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or (_22704_, _02439_, _02437_);
  and (_02440_, _02326_, _23718_);
  and (_02441_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_22705_, _02441_, _02440_);
  and (_02442_, _02383_, _23718_);
  and (_02443_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or (_22706_, _02443_, _02442_);
  and (_02444_, _23842_, _23643_);
  and (_02446_, _02444_, _23676_);
  not (_02447_, _02444_);
  and (_02449_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_22707_, _02449_, _02446_);
  and (_02450_, _24615_, _24117_);
  not (_02451_, _02450_);
  and (_02452_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and (_02453_, _02450_, _23589_);
  or (_22708_, _02453_, _02452_);
  and (_02454_, _02326_, _23838_);
  and (_02456_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or (_22710_, _02456_, _02454_);
  and (_02457_, _02326_, _23791_);
  and (_02458_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_27271_, _02458_, _02457_);
  and (_02459_, _24541_, _24118_);
  and (_02460_, _02459_, _23982_);
  not (_02462_, _02459_);
  and (_02463_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or (_27228_, _02463_, _02460_);
  and (_02465_, _24796_, _24633_);
  and (_02466_, _02465_, _24688_);
  nand (_02468_, _02466_, _23522_);
  or (_02469_, _02466_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_02471_, _25316_, _24714_);
  not (_02472_, _02471_);
  and (_02473_, _02472_, _02469_);
  and (_02474_, _02473_, _02468_);
  nor (_02475_, _02472_, _23748_);
  or (_02477_, _02475_, _02474_);
  and (_22711_, _02477_, _22761_);
  and (_02478_, _02465_, _23919_);
  and (_02479_, _02478_, _23522_);
  nor (_02480_, _02478_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_02481_, _02480_, _02479_);
  nand (_02482_, _02481_, _02472_);
  nand (_02483_, _02471_, _23628_);
  and (_02484_, _02483_, _22761_);
  and (_22712_, _02484_, _02482_);
  not (_02485_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02486_, _23985_, _23918_);
  nor (_02487_, _02486_, _02485_);
  or (_02488_, _02487_, _24732_);
  and (_02490_, _02488_, _02465_);
  nand (_02491_, _02486_, _24731_);
  nand (_02492_, _02465_, _02491_);
  and (_02493_, _02492_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02494_, _02493_, _02471_);
  or (_02495_, _02494_, _02490_);
  nand (_02496_, _02471_, _23914_);
  and (_02497_, _02496_, _22761_);
  and (_22713_, _02497_, _02495_);
  and (_02498_, _24636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_02499_, _02498_, _24635_);
  and (_02500_, _02499_, _02465_);
  nand (_02501_, _02465_, _23012_);
  and (_02502_, _02501_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_02503_, _02502_, _02471_);
  or (_02504_, _02503_, _02500_);
  nand (_02505_, _02471_, _23832_);
  and (_02506_, _02505_, _22761_);
  and (_22714_, _02506_, _02504_);
  not (_02508_, _23992_);
  nor (_02509_, _02508_, _23522_);
  not (_02510_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_02512_, _23992_, _02510_);
  nand (_02513_, _02512_, _02465_);
  or (_02514_, _02513_, _02509_);
  nor (_02516_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_02517_, _02516_);
  nor (_02518_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_02519_, _02518_, _02517_);
  and (_02520_, _02519_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_02521_, _02519_, _02510_);
  or (_02522_, _02521_, _02520_);
  or (_02524_, _02522_, _02465_);
  and (_02525_, _02524_, _02514_);
  or (_02526_, _02525_, _02471_);
  or (_02527_, _02472_, _23709_);
  and (_02528_, _02527_, _22761_);
  and (_22715_, _02528_, _02526_);
  or (_02530_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_02531_, _02530_, _02465_);
  not (_02532_, _23878_);
  nor (_02533_, _02532_, _23522_);
  nand (_02535_, _02532_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_02536_, _02535_, _02465_);
  or (_02537_, _02536_, _02533_);
  and (_02538_, _02537_, _02531_);
  or (_02539_, _02538_, _02471_);
  nand (_02540_, _02471_, _23784_);
  and (_02542_, _02540_, _22761_);
  and (_22716_, _02542_, _02539_);
  not (_02543_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_02544_, _02543_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_02545_, _02544_, _02516_);
  and (_02546_, _02545_, _02518_);
  or (_02547_, _02546_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02548_, _02547_, _02465_);
  and (_02549_, _24713_, _23812_);
  not (_02550_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02552_, _24713_, _02550_);
  nand (_02553_, _02552_, _02465_);
  or (_02554_, _02553_, _02549_);
  and (_02556_, _02554_, _02548_);
  or (_02557_, _02556_, _02471_);
  nand (_02558_, _02471_, _23669_);
  and (_02559_, _02558_, _22761_);
  and (_22717_, _02559_, _02557_);
  or (_02560_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_02561_, _02560_, _22761_);
  nand (_02562_, _02086_, _23748_);
  and (_22718_, _02562_, _02561_);
  or (_02563_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_02564_, _02563_, _22761_);
  nand (_02565_, _02086_, _23628_);
  and (_22719_, _02565_, _02564_);
  or (_02566_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_02567_, _02566_, _22761_);
  nand (_02568_, _02086_, _23832_);
  and (_22720_, _02568_, _02567_);
  or (_02570_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_02571_, _02570_, _22761_);
  nand (_02572_, _02086_, _23784_);
  and (_22721_, _02572_, _02571_);
  nand (_02573_, _02086_, _23669_);
  or (_02575_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_02576_, _02575_, _22761_);
  and (_22722_, _02576_, _02573_);
  not (_02578_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_02579_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_02580_, _02579_, _02516_);
  and (_02581_, _02517_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_02582_, _02581_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02583_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_02585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02586_, _02585_, _02583_);
  and (_02587_, _02586_, _02582_);
  nor (_02588_, _02587_, _02580_);
  nor (_02589_, _02588_, _02578_);
  and (_02590_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_02591_, _02590_, _02589_);
  and (_02592_, _25316_, _23883_);
  nor (_02593_, _02592_, _02591_);
  not (_02594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_02595_, _02594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_02596_, _02595_, _02517_);
  and (_02598_, _02596_, _02592_);
  or (_02599_, _02598_, _02593_);
  and (_22723_, _02599_, _22761_);
  and (_02601_, _02592_, _02517_);
  nand (_02602_, _02601_, _23585_);
  and (_02603_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  not (_02604_, _02588_);
  and (_02606_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_02607_, _02606_, _02603_);
  or (_02608_, _02607_, _02592_);
  and (_02609_, _02608_, _22761_);
  and (_22724_, _02609_, _02602_);
  not (_02610_, _23748_);
  and (_02611_, _02601_, _02610_);
  and (_02613_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_02614_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_02615_, _02614_, _02613_);
  nor (_02616_, _02615_, _02592_);
  not (_02618_, _23585_);
  and (_02619_, _02592_, _02516_);
  and (_02621_, _02619_, _02618_);
  or (_02622_, _02621_, _02616_);
  or (_02623_, _02622_, _02611_);
  and (_22725_, _02623_, _22761_);
  and (_02624_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_02625_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_02626_, _02625_, _02624_);
  nor (_02628_, _02626_, _02592_);
  not (_02629_, _23628_);
  and (_02630_, _02601_, _02629_);
  and (_02632_, _02619_, _02610_);
  or (_02633_, _02632_, _02630_);
  or (_02634_, _02633_, _02628_);
  and (_22726_, _02634_, _22761_);
  and (_02635_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02636_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_02638_, _02636_, _02635_);
  nor (_02639_, _02638_, _02592_);
  not (_02640_, _23914_);
  and (_02642_, _02601_, _02640_);
  or (_02643_, _02642_, _02639_);
  and (_02644_, _02619_, _02629_);
  or (_02645_, _02644_, _02643_);
  and (_22727_, _02645_, _22761_);
  and (_02646_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02647_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_02649_, _02647_, _02646_);
  nor (_02650_, _02649_, _02592_);
  not (_02651_, _23832_);
  and (_02652_, _02601_, _02651_);
  or (_02654_, _02652_, _02650_);
  and (_02655_, _02619_, _02640_);
  or (_02656_, _02655_, _02654_);
  and (_22728_, _02656_, _22761_);
  and (_02658_, _02619_, _02651_);
  and (_02659_, _02601_, _23709_);
  and (_02660_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_02662_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02663_, _02662_, _02660_);
  nor (_02664_, _02663_, _02592_);
  or (_02665_, _02664_, _02659_);
  or (_02666_, _02665_, _02658_);
  and (_22730_, _02666_, _22761_);
  and (_02667_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_02668_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_02669_, _02668_, _02667_);
  nor (_02670_, _02669_, _02592_);
  not (_02671_, _23784_);
  and (_02672_, _02601_, _02671_);
  and (_02673_, _02619_, _23709_);
  or (_02674_, _02673_, _02672_);
  or (_02675_, _02674_, _02670_);
  and (_22731_, _02675_, _22761_);
  and (_02676_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_02677_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02678_, _02677_, _02676_);
  nor (_02679_, _02678_, _02592_);
  and (_02680_, _02601_, _24763_);
  or (_02681_, _02680_, _02679_);
  and (_02682_, _02619_, _02671_);
  or (_02683_, _02682_, _02681_);
  and (_22732_, _02683_, _22761_);
  or (_02684_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_02685_, _02580_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_02686_, _02685_, _02587_);
  and (_02687_, _02686_, _02684_);
  nor (_02688_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor (_02689_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02690_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02691_, _02690_, _02689_);
  and (_02692_, _02691_, _02688_);
  nor (_02693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02695_, _02694_, _02693_);
  and (_02696_, _02695_, _02580_);
  and (_02697_, _02696_, _02692_);
  and (_02698_, _02697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_02699_, _02698_, _02687_);
  nor (_02700_, _02699_, _02592_);
  and (_02701_, _02619_, _24763_);
  or (_02702_, _02701_, _02700_);
  and (_22733_, _02702_, _22761_);
  not (_02703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_02704_, _02516_, _02703_);
  and (_02705_, _02704_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_02706_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_02707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _02706_);
  not (_02708_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02709_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _02708_);
  and (_02710_, _02709_, _02707_);
  and (_02711_, _02710_, _02705_);
  and (_02712_, _02703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02713_, _02516_, _02550_);
  and (_02714_, _02713_, _02712_);
  and (_02715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02716_, _02715_, _02517_);
  nor (_02717_, _02716_, _02714_);
  nor (_02718_, _02717_, _02705_);
  or (_02719_, _02718_, _02711_);
  and (_02720_, _02516_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02721_, _02720_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_02722_, _02721_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_02723_, _02722_, _02719_);
  nor (_02724_, _02721_, _02711_);
  or (_02725_, _02724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02726_, _02725_, _02100_);
  and (_02727_, _02726_, _02723_);
  or (_22734_, _02727_, _02099_);
  not (_02728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_02729_, _02724_);
  nor (_02730_, _02729_, _02718_);
  nor (_02731_, _02730_, _02728_);
  or (_02732_, _02731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_02733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _02728_);
  or (_02734_, _02733_, _02724_);
  and (_02735_, _02734_, _22761_);
  and (_22735_, _02735_, _02732_);
  and (_02736_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02737_, _02729_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not (_02738_, _02705_);
  nor (_02739_, _02710_, _02738_);
  and (_02740_, _02739_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_02741_, _02716_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nand (_02742_, _02741_, _02738_);
  nor (_02743_, _02742_, _02714_);
  nor (_02744_, _02743_, _02740_);
  nor (_02745_, _02744_, _02721_);
  or (_02746_, _02745_, _02737_);
  and (_02747_, _02746_, _02100_);
  or (_22736_, _02747_, _02736_);
  and (_02748_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and (_02749_, _02233_, _23838_);
  or (_22737_, _02749_, _02748_);
  and (_02750_, _01801_, _23854_);
  and (_02751_, _02750_, _23755_);
  not (_02752_, _02750_);
  and (_02753_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_22738_, _02753_, _02751_);
  and (_02754_, _02750_, _23635_);
  and (_02755_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_22739_, _02755_, _02754_);
  and (_02756_, _02750_, _23982_);
  and (_02757_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_22740_, _02757_, _02756_);
  and (_02758_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and (_02759_, _02233_, _23718_);
  or (_22741_, _02759_, _02758_);
  and (_02760_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  and (_02761_, _02450_, _23791_);
  or (_22742_, _02761_, _02760_);
  and (_02762_, _24768_, _24558_);
  not (_02763_, _02762_);
  and (_02764_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and (_02765_, _02762_, _23635_);
  or (_27062_, _02765_, _02764_);
  and (_02766_, _02750_, _23589_);
  and (_02767_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_22743_, _02767_, _02766_);
  and (_02768_, _01801_, _23797_);
  and (_02769_, _02768_, _23589_);
  not (_02770_, _02768_);
  and (_02771_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_22745_, _02771_, _02769_);
  and (_02772_, _02768_, _23755_);
  and (_02773_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_22746_, _02773_, _02772_);
  not (_02774_, _02730_);
  or (_02775_, _02774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_02776_, _02724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02777_, _02776_, _02100_);
  and (_02778_, _02777_, _02775_);
  or (_22747_, _02778_, _02104_);
  and (_02779_, _24572_, _24103_);
  and (_02780_, _02779_, _23718_);
  not (_02781_, _02779_);
  and (_02782_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_22748_, _02782_, _02780_);
  and (_02783_, _02779_, _23676_);
  and (_02784_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_22749_, _02784_, _02783_);
  and (_02785_, _02276_, _24117_);
  and (_02786_, _02785_, _23755_);
  not (_02787_, _02785_);
  and (_02788_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or (_22750_, _02788_, _02786_);
  and (_02789_, _02710_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_02790_, _02789_, _02717_);
  or (_02791_, _02790_, _02730_);
  and (_02792_, _02791_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02793_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _02728_);
  nand (_02794_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_02795_, _02794_, _02724_);
  or (_02796_, _02795_, _02793_);
  or (_02797_, _02796_, _02792_);
  and (_22751_, _02797_, _22761_);
  nor (_02798_, _02716_, _02705_);
  or (_02799_, _02798_, _02728_);
  or (_02800_, _02799_, _02708_);
  and (_02801_, _02705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02802_, _02801_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_02803_, _02802_, _22761_);
  and (_22752_, _02803_, _02800_);
  and (_02804_, _02459_, _23718_);
  and (_02805_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or (_27227_, _02805_, _02804_);
  and (_02806_, _02768_, _23635_);
  and (_02807_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_26946_, _02807_, _02806_);
  nand (_02808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22761_);
  nor (_02809_, _02808_, _02731_);
  or (_02810_, _02790_, _02729_);
  and (_02811_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_02812_, _02811_, _02810_);
  or (_22753_, _02812_, _02809_);
  and (_02813_, _02799_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_02814_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02815_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02816_, _02815_, _02814_);
  and (_02817_, _02816_, _02801_);
  or (_02818_, _02817_, _02813_);
  and (_22754_, _02818_, _22761_);
  and (_02819_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and (_02820_, _02762_, _23755_);
  or (_22755_, _02820_, _02819_);
  or (_02821_, _02582_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_02822_, _02582_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_02823_, _02822_, rst);
  nand (_02824_, _02823_, _02821_);
  nor (_22756_, _02824_, _02592_);
  and (_02825_, _02814_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02826_, _02825_, _02706_);
  and (_02827_, _02801_, _02826_);
  or (_02828_, _02827_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not (_02829_, rxd_i);
  nand (_02830_, _02827_, _02829_);
  and (_02831_, _02830_, _22761_);
  and (_22757_, _02831_, _02828_);
  or (_02832_, _02822_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_02833_, _02822_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02834_, _02833_, rst);
  nand (_02835_, _02834_, _02832_);
  nor (_22758_, _02835_, _02592_);
  nor (_02836_, _02833_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_02837_, _02833_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_02838_, _02837_, _02836_);
  nand (_02839_, _02838_, _22761_);
  nor (_22759_, _02839_, _02592_);
  and (_02840_, _24615_, _23649_);
  not (_02841_, _02840_);
  and (_02842_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  and (_02843_, _02840_, _23718_);
  or (_22760_, _02843_, _02842_);
  and (_02845_, _24768_, _23028_);
  and (_02847_, _02845_, _23791_);
  not (_02848_, _02845_);
  and (_02849_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_27275_, _02849_, _02847_);
  or (_02850_, _02731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_02851_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _02728_);
  or (_02852_, _02851_, _02724_);
  and (_02853_, _02852_, _22761_);
  and (_22766_, _02853_, _02850_);
  and (_02854_, _02750_, _23791_);
  and (_02855_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_26966_, _02855_, _02854_);
  and (_02856_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  and (_02857_, _02762_, _23791_);
  or (_27060_, _02857_, _02856_);
  and (_02858_, _24615_, _24541_);
  not (_02859_, _02858_);
  and (_02860_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and (_02861_, _02858_, _23676_);
  or (_22786_, _02861_, _02860_);
  and (_02862_, _24117_, _23028_);
  and (_02863_, _02862_, _23982_);
  not (_02864_, _02862_);
  and (_02865_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_22793_, _02865_, _02863_);
  and (_02866_, _02750_, _23676_);
  and (_02867_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_22806_, _02867_, _02866_);
  and (_02868_, _02799_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_02869_, _02825_, _02738_);
  or (_02870_, _02869_, _02868_);
  and (_02871_, _02814_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02872_, _02871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02873_, _02872_, _22761_);
  and (_22819_, _02873_, _02870_);
  and (_02874_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_22831_, _02874_, _02736_);
  and (_02875_, _24597_, _23838_);
  and (_02876_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or (_22845_, _02876_, _02875_);
  and (_02877_, _24118_, _23803_);
  and (_02878_, _02877_, _23755_);
  not (_02879_, _02877_);
  and (_02880_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_27233_, _02880_, _02878_);
  and (_02881_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02882_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_22851_, _02882_, _02881_);
  and (_02883_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02884_, _02883_, _02793_);
  and (_22859_, _02884_, _22761_);
  and (_02885_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and (_02886_, _02762_, _23838_);
  or (_27061_, _02886_, _02885_);
  and (_02887_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02888_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_22879_, _02888_, _02887_);
  and (_02889_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  and (_02890_, _02762_, _23718_);
  or (_22882_, _02890_, _02889_);
  and (_02891_, _02768_, _23791_);
  and (_02892_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_22888_, _02892_, _02891_);
  or (_02893_, _02731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02894_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _02728_);
  or (_02895_, _02894_, _02724_);
  and (_02896_, _02895_, _22761_);
  and (_22894_, _02896_, _02893_);
  or (_02897_, _02774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_02898_, _02724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02899_, _02898_, _02100_);
  and (_02900_, _02899_, _02897_);
  or (_22898_, _02900_, _02102_);
  or (_02901_, _02731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _02728_);
  or (_02903_, _02902_, _02724_);
  and (_02904_, _02903_, _22761_);
  and (_22901_, _02904_, _02901_);
  or (_02905_, _02731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _02728_);
  or (_02908_, _02906_, _02724_);
  and (_02909_, _02908_, _22761_);
  and (_22904_, _02909_, _02905_);
  and (_02910_, _02768_, _23676_);
  and (_02911_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_22907_, _02911_, _02910_);
  and (_02912_, _02444_, _23791_);
  and (_02913_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_22935_, _02913_, _02912_);
  and (_02914_, _24572_, _23594_);
  and (_02915_, _02914_, _23589_);
  not (_02916_, _02914_);
  and (_02917_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_22961_, _02917_, _02915_);
  and (_26869_[4], _24436_, _22761_);
  and (_02918_, _02914_, _23635_);
  and (_02919_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_23026_, _02919_, _02918_);
  and (_02920_, _02877_, _23589_);
  and (_02921_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_23036_, _02921_, _02920_);
  and (_02922_, _23864_, _23838_);
  and (_02923_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_23048_, _02923_, _02922_);
  and (_02924_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and (_02925_, _02450_, _23676_);
  or (_23053_, _02925_, _02924_);
  and (_02926_, _02768_, _23838_);
  and (_02927_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_23079_, _02927_, _02926_);
  and (_02928_, _02862_, _23635_);
  and (_02929_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_23085_, _02929_, _02928_);
  and (_02931_, _02862_, _23755_);
  and (_02932_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_23094_, _02932_, _02931_);
  and (_02933_, _02914_, _23838_);
  and (_02934_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_23097_, _02934_, _02933_);
  and (_02935_, _02914_, _23791_);
  and (_02936_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_27147_, _02936_, _02935_);
  and (_02937_, _24572_, _23863_);
  and (_02938_, _02937_, _23676_);
  not (_02939_, _02937_);
  and (_02940_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or (_27149_, _02940_, _02938_);
  and (_02941_, _02436_, _23589_);
  and (_02942_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or (_23144_, _02942_, _02941_);
  and (_02943_, _24573_, _23589_);
  and (_02945_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or (_23157_, _02945_, _02943_);
  and (_02947_, _01801_, _24768_);
  and (_02948_, _02947_, _23635_);
  not (_02950_, _02947_);
  and (_02951_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_23173_, _02951_, _02948_);
  and (_02953_, _02947_, _23982_);
  and (_02954_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_23186_, _02954_, _02953_);
  and (_02956_, _23864_, _23676_);
  and (_02957_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_23201_, _02957_, _02956_);
  and (_02958_, _02947_, _23838_);
  and (_02960_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_23204_, _02960_, _02958_);
  and (_02961_, _01416_, _01447_);
  and (_02962_, _02961_, _01487_);
  and (_02963_, _01440_, _01421_);
  or (_02964_, _02963_, _02962_);
  and (_02966_, _01439_, _01454_);
  nor (_02968_, _01549_, _02966_);
  or (_02969_, _01454_, _01405_);
  nand (_02970_, _02969_, _01476_);
  nand (_02971_, _02970_, _02968_);
  or (_02972_, _02971_, _02964_);
  or (_02974_, _01464_, _01504_);
  or (_02975_, _01525_, _01510_);
  or (_02976_, _02975_, _02974_);
  or (_02977_, _01526_, _01410_);
  or (_02978_, _02977_, _02976_);
  and (_02979_, _01440_, _01445_);
  and (_02980_, _01456_, _01406_);
  or (_02981_, _02980_, _02979_);
  and (_02982_, _01428_, _01412_);
  or (_02983_, _02982_, _01493_);
  and (_02984_, _01470_, _01451_);
  or (_02985_, _01557_, _02984_);
  or (_02986_, _02985_, _02983_);
  or (_02987_, _02986_, _02981_);
  or (_02988_, _02987_, _02978_);
  or (_02989_, _02988_, _02972_);
  and (_02990_, _02989_, _22769_);
  and (_02991_, _22764_, _22765_);
  and (_02993_, _02991_, _26569_);
  nor (_02994_, _02993_, _24526_);
  or (_02996_, _02994_, rst);
  or (_26872_[1], _02996_, _02990_);
  and (_02998_, _02947_, _23755_);
  and (_03000_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_23250_, _03000_, _02998_);
  and (_03001_, _24768_, _23599_);
  and (_03003_, _03001_, _23718_);
  not (_03004_, _03001_);
  and (_03005_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or (_27249_, _03005_, _03003_);
  and (_03006_, _24103_, _23643_);
  and (_03007_, _03006_, _23982_);
  not (_03008_, _03006_);
  and (_03009_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or (_23272_, _03009_, _03007_);
  and (_03010_, _01801_, _24541_);
  and (_03012_, _03010_, _23589_);
  not (_03013_, _03010_);
  and (_03014_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_23294_, _03014_, _03012_);
  and (_03015_, _24572_, _23803_);
  and (_03016_, _03015_, _23791_);
  not (_03017_, _03015_);
  and (_03018_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_23331_, _03018_, _03016_);
  and (_03019_, _03006_, _23755_);
  and (_03021_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or (_23336_, _03021_, _03019_);
  and (_03023_, _03006_, _23635_);
  and (_03024_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or (_23343_, _03024_, _03023_);
  and (_03025_, _02947_, _23791_);
  and (_03027_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_23357_, _03027_, _03025_);
  and (_03028_, _03010_, _23676_);
  and (_03029_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_23396_, _03029_, _03028_);
  and (_03030_, _03006_, _23718_);
  and (_03031_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or (_23400_, _03031_, _03030_);
  and (_03032_, _01801_, _24117_);
  and (_03033_, _03032_, _23589_);
  not (_03034_, _03032_);
  and (_03035_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_23421_, _03035_, _03033_);
  and (_03037_, _02069_, _23676_);
  and (_03038_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_27251_, _03038_, _03037_);
  and (_03039_, _03010_, _23838_);
  and (_03040_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_23450_, _03040_, _03039_);
  and (_03041_, _03015_, _23718_);
  and (_03042_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_23516_, _03042_, _03041_);
  and (_03043_, _24769_, _23635_);
  and (_03044_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or (_23539_, _03044_, _03043_);
  and (_03046_, _23594_, _23028_);
  and (_03047_, _03046_, _23635_);
  not (_03048_, _03046_);
  and (_03050_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_23559_, _03050_, _03047_);
  and (_03051_, _03046_, _23589_);
  and (_03052_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_23600_, _03052_, _03051_);
  nor (_03053_, _26727_, _26697_);
  not (_03054_, _26682_);
  nor (_03055_, _26714_, _03054_);
  and (_03056_, _03055_, _03053_);
  nor (_03057_, _00274_, _26585_);
  and (_03058_, _26609_, _24445_);
  nor (_03059_, _03058_, _26720_);
  and (_03061_, _03059_, _26696_);
  and (_03062_, _03061_, _03057_);
  and (_03063_, _03062_, _03056_);
  nor (_03064_, _03057_, _00224_);
  nor (_03065_, _03064_, _26575_);
  nor (_03066_, _03065_, _03063_);
  and (_26921_, _03066_, _22761_);
  and (_03067_, _25949_, _25523_);
  nand (_03068_, _03067_, _23585_);
  or (_03069_, _03067_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_03070_, _03069_, _22761_);
  and (_26883_[7], _03070_, _03068_);
  not (_03072_, _25950_);
  nor (_03073_, _03072_, _23585_);
  and (_03074_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03075_, _03074_, _25946_);
  or (_03076_, _03075_, _03073_);
  or (_03077_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03078_, _03077_, _22761_);
  and (_26884_[7], _03078_, _03076_);
  and (_03079_, _25956_, _25952_);
  or (_03080_, _03079_, _25946_);
  and (_03081_, _03080_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_03082_, _25956_, _23585_);
  not (_03083_, _25952_);
  and (_03084_, _03083_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_03085_, _03084_, _03082_);
  and (_03086_, _03085_, _25523_);
  or (_03087_, _03086_, _03081_);
  and (_26885_[7], _03087_, _22761_);
  and (_03088_, _25958_, _25523_);
  not (_03089_, _03088_);
  nor (_03090_, _03089_, _23585_);
  and (_03091_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_03092_, _03091_, _03090_);
  and (_26886_[7], _03092_, _22761_);
  and (_03093_, _25611_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_03094_, _25611_, _23585_);
  or (_03095_, _03094_, _03093_);
  and (_26887_[7], _03095_, _22761_);
  nor (_03096_, _25531_, _23585_);
  not (_03097_, _25528_);
  nand (_03098_, _25959_, _03097_);
  and (_03099_, _03098_, _25523_);
  not (_03100_, _03099_);
  and (_03101_, _03100_, _03080_);
  or (_03102_, _03101_, _03083_);
  and (_03103_, _03102_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand (_03104_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_03105_, _03104_, _25960_);
  or (_03106_, _03105_, _03103_);
  or (_03107_, _03106_, _03096_);
  and (_26888_[7], _03107_, _22761_);
  and (_03109_, _25965_, _25959_);
  or (_03110_, _03109_, _25946_);
  or (_03111_, _03110_, _03098_);
  and (_03112_, _03111_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_03113_, _25964_, _25523_);
  not (_03114_, _03113_);
  nor (_03115_, _03114_, _23585_);
  or (_03116_, _03115_, _03112_);
  and (_26889_[7], _03116_, _22761_);
  and (_03117_, _25963_, _25523_);
  and (_03118_, _03117_, _02618_);
  nand (_03119_, _03109_, _03079_);
  or (_03120_, _03119_, _25970_);
  and (_03121_, _03120_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_03122_, _03121_, _03118_);
  and (_26890_[7], _03122_, _22761_);
  and (_03124_, _25301_, _23676_);
  and (_03125_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_23675_, _03125_, _03124_);
  and (_03126_, _03010_, _23718_);
  and (_03127_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_23679_, _03127_, _03126_);
  and (_03128_, _02322_, _23982_);
  and (_03130_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_23686_, _03130_, _03128_);
  and (_03132_, _03010_, _23791_);
  and (_03133_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_23689_, _03133_, _03132_);
  and (_03134_, _23643_, _23594_);
  and (_03135_, _03134_, _23718_);
  not (_03136_, _03134_);
  and (_03137_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or (_23708_, _03137_, _03135_);
  and (_03138_, _03032_, _23676_);
  and (_03139_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_27292_, _03139_, _03138_);
  and (_03140_, _03032_, _23718_);
  and (_03141_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_23761_, _03141_, _03140_);
  and (_03142_, _03032_, _23791_);
  and (_03143_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_23764_, _03143_, _03142_);
  and (_03144_, _24089_, _23755_);
  and (_03145_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_27080_, _03145_, _03144_);
  and (_03147_, _03032_, _23635_);
  and (_03148_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_23856_, _03148_, _03147_);
  and (_03149_, _03032_, _23982_);
  and (_03150_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_23860_, _03150_, _03149_);
  and (_03151_, _24089_, _23589_);
  and (_03152_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_23905_, _03152_, _03151_);
  and (_03154_, _01801_, _23641_);
  and (_03155_, _03154_, _23791_);
  not (_03156_, _03154_);
  and (_03157_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_23912_, _03157_, _03155_);
  and (_03158_, _03001_, _23791_);
  and (_03159_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or (_23957_, _03159_, _03158_);
  and (_03160_, _03154_, _23838_);
  and (_03161_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_23960_, _03161_, _03160_);
  and (_03162_, _03154_, _23718_);
  and (_03163_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_23965_, _03163_, _03162_);
  and (_03165_, _03134_, _23635_);
  and (_03166_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or (_27081_, _03166_, _03165_);
  and (_03167_, _03134_, _23982_);
  and (_03168_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or (_23970_, _03168_, _03167_);
  and (_03169_, _03154_, _23635_);
  and (_03170_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_27270_, _03170_, _03169_);
  and (_03171_, _03154_, _23589_);
  and (_03173_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_24008_, _03173_, _03171_);
  and (_03174_, _03154_, _23755_);
  and (_03175_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_24014_, _03175_, _03174_);
  and (_03176_, _23843_, _23838_);
  and (_03177_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or (_24022_, _03177_, _03176_);
  and (_03178_, _03134_, _23589_);
  and (_03179_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or (_24060_, _03179_, _03178_);
  and (_03180_, _03134_, _23755_);
  and (_03181_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or (_24066_, _03181_, _03180_);
  and (_03183_, _24571_, _23650_);
  and (_03184_, _03183_, _24078_);
  not (_03185_, _03184_);
  and (_03187_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  and (_03188_, _03184_, _23718_);
  or (_24076_, _03188_, _03187_);
  and (_03189_, _01801_, _23863_);
  and (_03191_, _03189_, _23982_);
  not (_03192_, _03189_);
  and (_03193_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_24079_, _03193_, _03191_);
  and (_03195_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  and (_03196_, _03184_, _23791_);
  or (_24082_, _03196_, _03195_);
  and (_03198_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and (_03199_, _03184_, _23676_);
  or (_27124_, _03199_, _03198_);
  and (_03201_, _03189_, _23589_);
  and (_03202_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_24114_, _03202_, _03201_);
  and (_03203_, _03189_, _23755_);
  and (_03204_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_24143_, _03204_, _03203_);
  and (_03205_, _03183_, _23017_);
  not (_03206_, _03205_);
  and (_03207_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  and (_03208_, _03205_, _23982_);
  or (_27142_, _03208_, _03207_);
  and (_03210_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  and (_03211_, _03205_, _23635_);
  or (_24151_, _03211_, _03210_);
  and (_03212_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  and (_03213_, _03205_, _23589_);
  or (_24157_, _03213_, _03212_);
  and (_03214_, _01801_, _24103_);
  and (_03215_, _03214_, _23755_);
  not (_03216_, _03214_);
  and (_03217_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_24163_, _03217_, _03215_);
  and (_03218_, _03214_, _23635_);
  and (_03219_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_24167_, _03219_, _03218_);
  and (_03220_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  and (_03221_, _03184_, _23635_);
  or (_24173_, _03221_, _03220_);
  and (_03222_, _03214_, _23982_);
  and (_03223_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_24175_, _03223_, _03222_);
  and (_03225_, _03214_, _23838_);
  and (_03226_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_24177_, _03226_, _03225_);
  and (_03227_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and (_03228_, _03184_, _23982_);
  or (_24185_, _03228_, _03227_);
  and (_03229_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and (_03231_, _03184_, _23838_);
  or (_24188_, _03231_, _03229_);
  and (_03232_, _23642_, _22933_);
  and (_03233_, _03232_, _23023_);
  and (_03234_, _03233_, _24078_);
  and (_03235_, _03234_, _23755_);
  not (_03236_, _03234_);
  and (_03237_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or (_26988_, _03237_, _03235_);
  and (_03238_, _03189_, _23791_);
  and (_03239_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_24202_, _03239_, _03238_);
  and (_03241_, _02276_, _23849_);
  and (_03242_, _03241_, _23718_);
  not (_03244_, _03241_);
  and (_03245_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  or (_24205_, _03245_, _03242_);
  and (_03246_, _03189_, _23676_);
  and (_03247_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_24208_, _03247_, _03246_);
  and (_03248_, _03214_, _23589_);
  and (_03249_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_24212_, _03249_, _03248_);
  and (_03250_, _02276_, _23803_);
  and (_03251_, _03250_, _23838_);
  not (_03253_, _03250_);
  and (_03254_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  or (_24230_, _03254_, _03251_);
  and (_03255_, _03183_, _23649_);
  not (_03256_, _03255_);
  and (_03257_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_03259_, _03255_, _23718_);
  or (_24249_, _03259_, _03257_);
  and (_03260_, _02276_, _23641_);
  and (_03261_, _03260_, _23982_);
  not (_03262_, _03260_);
  and (_03263_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_24284_, _03263_, _03261_);
  and (_03264_, _02276_, _23863_);
  and (_03265_, _03264_, _23755_);
  not (_03266_, _03264_);
  and (_03267_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_24287_, _03267_, _03265_);
  and (_03269_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_03270_, _03255_, _23838_);
  or (_24290_, _03270_, _03269_);
  and (_03271_, _03264_, _23676_);
  and (_03272_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_24293_, _03272_, _03271_);
  and (_03273_, _01801_, _23594_);
  and (_03274_, _03273_, _23589_);
  not (_03275_, _03273_);
  and (_03276_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_24298_, _03276_, _03274_);
  and (_03277_, _02276_, _24103_);
  and (_03278_, _03277_, _23718_);
  not (_03279_, _03277_);
  and (_03280_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  or (_27182_, _03280_, _03278_);
  and (_03281_, _02276_, _23962_);
  and (_03282_, _03281_, _23838_);
  not (_03283_, _03281_);
  and (_03284_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_24312_, _03284_, _03282_);
  and (_03285_, _03046_, _23755_);
  and (_03286_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_24315_, _03286_, _03285_);
  and (_03287_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_03288_, _03255_, _23635_);
  or (_24320_, _03288_, _03287_);
  and (_03290_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_03291_, _03255_, _23589_);
  or (_24323_, _03291_, _03290_);
  and (_03292_, _03214_, _23791_);
  and (_03293_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_24326_, _03293_, _03292_);
  and (_03294_, _03214_, _23676_);
  and (_03295_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_24333_, _03295_, _03294_);
  and (_03296_, _24572_, _23849_);
  and (_03297_, _03296_, _23791_);
  not (_03298_, _03296_);
  and (_03299_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_24339_, _03299_, _03297_);
  and (_03300_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_03301_, _03255_, _23755_);
  or (_24342_, _03301_, _03300_);
  and (_03302_, _02276_, _23797_);
  and (_03303_, _03302_, _23718_);
  not (_03304_, _03302_);
  and (_03305_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  or (_24345_, _03305_, _03303_);
  and (_03306_, _25742_, _23635_);
  and (_03307_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_27268_, _03307_, _03306_);
  and (_03308_, _03273_, _23676_);
  and (_03309_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_24355_, _03309_, _03308_);
  and (_03310_, _03273_, _23718_);
  and (_03311_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_27226_, _03311_, _03310_);
  and (_03312_, _03273_, _23791_);
  and (_03313_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_24370_, _03313_, _03312_);
  and (_03314_, _03183_, _23594_);
  not (_03315_, _03314_);
  and (_03316_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_03317_, _03314_, _23589_);
  or (_24434_, _03317_, _03316_);
  and (_03318_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  and (_03319_, _03205_, _23838_);
  or (_24437_, _03319_, _03318_);
  and (_03320_, _03273_, _23982_);
  and (_03321_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_24442_, _03321_, _03320_);
  and (_03322_, _24572_, _23649_);
  and (_03323_, _03322_, _23791_);
  not (_03324_, _03322_);
  and (_03325_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_24444_, _03325_, _03323_);
  and (_03326_, _02276_, _23017_);
  and (_03327_, _03326_, _23791_);
  not (_03328_, _03326_);
  and (_03329_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_24455_, _03329_, _03327_);
  nor (_26869_[5], _24385_, rst);
  nor (_26869_[6], _24363_, rst);
  and (_03330_, _03322_, _23589_);
  and (_03331_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_24462_, _03331_, _03330_);
  and (_03332_, _03322_, _23982_);
  and (_03334_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_24467_, _03334_, _03332_);
  and (_03335_, _02276_, _23842_);
  and (_03336_, _03335_, _23791_);
  not (_03337_, _03335_);
  and (_03338_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_27192_, _03338_, _03336_);
  and (_03340_, _01801_, _23962_);
  and (_03341_, _03340_, _23982_);
  not (_03343_, _03340_);
  and (_03344_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_24477_, _03344_, _03341_);
  and (_03345_, _03322_, _23635_);
  and (_03346_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_27143_, _03346_, _03345_);
  and (_03348_, _02785_, _23838_);
  and (_03349_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  or (_27184_, _03349_, _03348_);
  and (_03350_, _03340_, _23838_);
  and (_03351_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_24498_, _03351_, _03350_);
  and (_03352_, _03340_, _23718_);
  and (_03353_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_24504_, _03353_, _03352_);
  and (_03354_, _02276_, _24541_);
  and (_03355_, _03354_, _23635_);
  not (_03356_, _03354_);
  and (_03357_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_24512_, _03357_, _03355_);
  and (_03358_, _24572_, _23017_);
  and (_03359_, _03358_, _23755_);
  not (_03360_, _03358_);
  and (_03361_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or (_24530_, _03361_, _03359_);
  and (_03362_, _03296_, _23635_);
  and (_03363_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_24532_, _03363_, _03362_);
  and (_03364_, _03340_, _23755_);
  and (_03365_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_24535_, _03365_, _03364_);
  and (_03367_, _03302_, _23755_);
  and (_03368_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  or (_24543_, _03368_, _03367_);
  and (_03369_, _03354_, _23838_);
  and (_03370_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_24548_, _03370_, _03369_);
  and (_03372_, _03340_, _23589_);
  and (_03373_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_24551_, _03373_, _03372_);
  and (_03374_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_03375_, _03314_, _23718_);
  or (_24553_, _03375_, _03374_);
  not (_03376_, _03067_);
  and (_03378_, _03376_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03379_, _03067_, _24763_);
  or (_03380_, _03379_, _03378_);
  and (_26883_[0], _03380_, _22761_);
  nand (_03381_, _03067_, _23784_);
  or (_03382_, _03067_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03383_, _03382_, _22761_);
  and (_26883_[1], _03383_, _03381_);
  or (_03384_, _03376_, _23709_);
  or (_03385_, _03067_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_03386_, _03385_, _22761_);
  and (_26883_[2], _03386_, _03384_);
  nand (_03388_, _03067_, _23832_);
  or (_03389_, _03067_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_03391_, _03389_, _22761_);
  and (_26883_[3], _03391_, _03388_);
  nand (_03392_, _03067_, _23914_);
  or (_03393_, _03067_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_03394_, _03393_, _22761_);
  and (_26883_[4], _03394_, _03392_);
  nand (_03395_, _03067_, _23628_);
  or (_03396_, _03067_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03397_, _03396_, _22761_);
  and (_26883_[5], _03397_, _03395_);
  nand (_03399_, _03067_, _23748_);
  or (_03400_, _03067_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03402_, _03400_, _22761_);
  and (_26883_[6], _03402_, _03399_);
  and (_03403_, _25950_, _24763_);
  and (_03404_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_03405_, _03404_, _25946_);
  or (_03406_, _03405_, _03403_);
  or (_03407_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_03408_, _03407_, _22761_);
  and (_26884_[0], _03408_, _03406_);
  nor (_03409_, _03072_, _23784_);
  and (_03410_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_03411_, _03410_, _25946_);
  or (_03412_, _03411_, _03409_);
  or (_03413_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03414_, _03413_, _22761_);
  and (_26884_[1], _03414_, _03412_);
  and (_03415_, _25950_, _23709_);
  and (_03416_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03417_, _03416_, _25946_);
  or (_03418_, _03417_, _03415_);
  or (_03420_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03421_, _03420_, _22761_);
  and (_26884_[2], _03421_, _03418_);
  nor (_03423_, _03072_, _23832_);
  and (_03424_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03425_, _03424_, _25946_);
  or (_03426_, _03425_, _03423_);
  or (_03427_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03429_, _03427_, _22761_);
  and (_26884_[3], _03429_, _03426_);
  nor (_03430_, _03072_, _23914_);
  and (_03431_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_03432_, _03431_, _25946_);
  or (_03433_, _03432_, _03430_);
  or (_03434_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_03435_, _03434_, _22761_);
  and (_26884_[4], _03435_, _03433_);
  nor (_03436_, _03072_, _23628_);
  and (_03437_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_03438_, _03437_, _25946_);
  or (_03439_, _03438_, _03436_);
  or (_03440_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_03441_, _03440_, _22761_);
  and (_26884_[5], _03441_, _03439_);
  nor (_03442_, _03072_, _23748_);
  and (_03443_, _03072_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03445_, _03443_, _25946_);
  or (_03446_, _03445_, _03442_);
  or (_03447_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03448_, _03447_, _22761_);
  and (_26884_[6], _03448_, _03446_);
  and (_03449_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_03450_, _03314_, _23791_);
  or (_24589_, _03450_, _03449_);
  nor (_03452_, _25952_, _25946_);
  or (_03453_, _03452_, _03080_);
  and (_03454_, _03453_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_03455_, _25946_, _23669_);
  and (_03456_, _03455_, _25955_);
  or (_03457_, _03456_, _03454_);
  and (_26885_[0], _03457_, _22761_);
  and (_03459_, _03453_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_03460_, _25955_, _25523_);
  and (_03461_, _03460_, _02671_);
  or (_03462_, _03461_, _03459_);
  and (_26885_[1], _03462_, _22761_);
  and (_03463_, _03453_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_03464_, _03460_, _23709_);
  or (_03466_, _03464_, _03463_);
  and (_26885_[2], _03466_, _22761_);
  and (_03467_, _03453_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_03469_, _03460_, _02651_);
  or (_03470_, _03469_, _03467_);
  and (_26885_[3], _03470_, _22761_);
  and (_03471_, _03453_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_03472_, _03460_, _02640_);
  or (_03473_, _03472_, _03471_);
  and (_26885_[4], _03473_, _22761_);
  and (_03474_, _03453_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_03475_, _03460_, _02629_);
  or (_03476_, _03475_, _03474_);
  and (_26885_[5], _03476_, _22761_);
  and (_03477_, _03453_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_03478_, _03460_, _02610_);
  or (_03479_, _03478_, _03477_);
  and (_26885_[6], _03479_, _22761_);
  and (_03480_, _03088_, _24763_);
  and (_03482_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_03483_, _03482_, _03480_);
  and (_26886_[0], _03483_, _22761_);
  nor (_03485_, _03089_, _23784_);
  and (_03486_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_03487_, _03486_, _03485_);
  and (_26886_[1], _03487_, _22761_);
  and (_03489_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_03490_, _03088_, _23709_);
  or (_03491_, _03490_, _03489_);
  and (_26886_[2], _03491_, _22761_);
  and (_03492_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_03493_, _03089_, _23832_);
  or (_03494_, _03493_, _03492_);
  and (_26886_[3], _03494_, _22761_);
  nor (_03495_, _03089_, _23914_);
  and (_03496_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_03497_, _03496_, _03495_);
  and (_26886_[4], _03497_, _22761_);
  nor (_03498_, _03089_, _23628_);
  and (_03499_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_03501_, _03499_, _03498_);
  and (_26886_[5], _03501_, _22761_);
  nor (_03503_, _03089_, _23748_);
  and (_03504_, _03089_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03505_, _03504_, _03503_);
  and (_26886_[6], _03505_, _22761_);
  or (_03506_, _25961_, _25946_);
  or (_03507_, _03506_, _25949_);
  and (_03508_, _03507_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or (_03509_, _25958_, _25955_);
  or (_03510_, _03509_, _25950_);
  and (_03511_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_03512_, _03511_, _03510_);
  or (_03513_, _03512_, _25751_);
  or (_03514_, _03513_, _03508_);
  and (_26887_[0], _03514_, _22761_);
  and (_03515_, _03507_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_03516_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_03517_, _03516_, _03510_);
  or (_03518_, _03517_, _25749_);
  or (_03519_, _03518_, _03515_);
  and (_26887_[1], _03519_, _22761_);
  and (_03521_, _25611_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_03522_, _25609_, _23709_);
  or (_03524_, _03522_, _03521_);
  and (_26887_[2], _03524_, _22761_);
  and (_03525_, _25611_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_03526_, _03525_, _26109_);
  and (_26887_[3], _03526_, _22761_);
  and (_03527_, _25611_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or (_03528_, _03527_, _25910_);
  and (_26887_[4], _03528_, _22761_);
  nor (_03529_, _25611_, _23628_);
  and (_03530_, _25611_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_03531_, _03530_, _03529_);
  and (_26887_[5], _03531_, _22761_);
  and (_03532_, _25611_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_03533_, _03532_, _25617_);
  and (_26887_[6], _03533_, _22761_);
  and (_03534_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_03535_, _03314_, _23676_);
  or (_24609_, _03535_, _03534_);
  and (_03536_, _03102_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand (_03537_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_03538_, _03537_, _25960_);
  and (_03539_, _25529_, _24763_);
  or (_03540_, _03539_, _03538_);
  or (_03541_, _03540_, _03536_);
  and (_26888_[0], _03541_, _22761_);
  and (_03543_, _03102_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nand (_03544_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_03545_, _03544_, _25960_);
  nor (_03546_, _25531_, _23784_);
  or (_03547_, _03546_, _03545_);
  or (_03548_, _03547_, _03543_);
  and (_26888_[1], _03548_, _22761_);
  and (_03549_, _25529_, _23709_);
  and (_03550_, _03102_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nand (_03552_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_03553_, _03552_, _25960_);
  or (_03554_, _03553_, _03550_);
  or (_03555_, _03554_, _03549_);
  and (_26888_[2], _03555_, _22761_);
  nor (_03556_, _25531_, _23832_);
  and (_03557_, _25531_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or (_03558_, _03557_, _03556_);
  and (_26888_[3], _03558_, _22761_);
  nor (_03560_, _25531_, _23914_);
  and (_03562_, _03102_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nand (_03563_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_03564_, _03563_, _25960_);
  or (_03565_, _03564_, _03562_);
  or (_03566_, _03565_, _03560_);
  and (_26888_[4], _03566_, _22761_);
  nor (_03567_, _25531_, _23628_);
  and (_03568_, _03101_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nand (_03569_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_03570_, _03569_, _25961_);
  or (_03571_, _03570_, _03568_);
  or (_03572_, _03571_, _03567_);
  and (_26888_[5], _03572_, _22761_);
  nor (_03573_, _25531_, _23748_);
  and (_03574_, _03102_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nand (_03576_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_03577_, _03576_, _25960_);
  or (_03579_, _03577_, _03574_);
  or (_03580_, _03579_, _03573_);
  and (_26888_[6], _03580_, _22761_);
  and (_03582_, _03113_, _24763_);
  or (_03583_, _03110_, _03099_);
  and (_03584_, _03583_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or (_03586_, _03584_, _03582_);
  and (_26889_[0], _03586_, _22761_);
  nor (_03587_, _03114_, _23784_);
  and (_03588_, _03583_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  or (_03589_, _03588_, _03587_);
  and (_26889_[1], _03589_, _22761_);
  and (_03591_, _03113_, _23709_);
  and (_03592_, _03114_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_03593_, _03592_, _03591_);
  and (_26889_[2], _03593_, _22761_);
  and (_03594_, _03114_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_03595_, _03114_, _23832_);
  or (_03596_, _03595_, _03594_);
  and (_26889_[3], _03596_, _22761_);
  nor (_03597_, _03114_, _23914_);
  and (_03599_, _03583_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or (_03600_, _03599_, _03597_);
  and (_26889_[4], _03600_, _22761_);
  nor (_03601_, _03114_, _23628_);
  and (_03602_, _03583_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_03603_, _03602_, _03601_);
  and (_26889_[5], _03603_, _22761_);
  nor (_03604_, _03114_, _23748_);
  and (_03605_, _03583_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_03606_, _03605_, _03604_);
  and (_26889_[6], _03606_, _22761_);
  or (_03607_, _03509_, _03083_);
  or (_03608_, _25970_, _03607_);
  and (_03609_, _03608_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_03610_, _25966_, _25608_);
  and (_03611_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03612_, _03611_, _03610_);
  and (_03613_, _03117_, _24763_);
  or (_03614_, _03613_, _03612_);
  or (_03615_, _03614_, _03609_);
  and (_26890_[0], _03615_, _22761_);
  and (_03616_, _03608_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_03617_, _25523_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_03618_, _03617_, _03610_);
  and (_03619_, _03117_, _02671_);
  or (_03620_, _03619_, _03618_);
  or (_03621_, _03620_, _03616_);
  and (_26890_[1], _03621_, _22761_);
  and (_03622_, _03117_, _23709_);
  and (_03623_, _03120_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_03624_, _03623_, _03622_);
  and (_26890_[2], _03624_, _22761_);
  or (_03625_, _03608_, _03610_);
  and (_03626_, _03625_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_03627_, _03117_, _02651_);
  or (_03628_, _03627_, _03626_);
  and (_26890_[3], _03628_, _22761_);
  and (_03629_, _03625_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_03630_, _03117_, _02640_);
  or (_03631_, _03630_, _03629_);
  and (_26890_[4], _03631_, _22761_);
  and (_03632_, _03625_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_03633_, _03117_, _02629_);
  or (_03634_, _03633_, _03632_);
  and (_26890_[5], _03634_, _22761_);
  and (_03635_, _03117_, _02610_);
  and (_03636_, _03610_, _25523_);
  or (_03637_, _03636_, _03608_);
  and (_03638_, _03637_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_03639_, _03638_, _03635_);
  and (_26890_[6], _03639_, _22761_);
  and (_03641_, _24615_, _23803_);
  not (_03643_, _03641_);
  and (_03644_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  and (_03645_, _03641_, _23755_);
  or (_24781_, _03645_, _03644_);
  and (_03646_, _03001_, _23982_);
  and (_03647_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or (_24878_, _03647_, _03646_);
  and (_03648_, _01801_, _24078_);
  and (_03650_, _03648_, _23755_);
  not (_03651_, _03648_);
  and (_03652_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_25007_, _03652_, _03650_);
  and (_03653_, _03250_, _23982_);
  and (_03654_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  or (_25057_, _03654_, _03653_);
  and (_03655_, _03001_, _23755_);
  and (_03656_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or (_25062_, _03656_, _03655_);
  and (_03657_, _24615_, _23863_);
  not (_03658_, _03657_);
  and (_03659_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_03660_, _03657_, _23589_);
  or (_25065_, _03660_, _03659_);
  and (_03662_, _03001_, _23635_);
  and (_03663_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or (_27250_, _03663_, _03662_);
  and (_03664_, _03648_, _23589_);
  and (_03665_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_25096_, _03665_, _03664_);
  and (_03666_, _02277_, _23676_);
  and (_03667_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or (_25112_, _03667_, _03666_);
  not (_03669_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03670_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_03671_, _03670_, _03669_);
  and (_03672_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _22761_);
  and (_27318_, _03672_, _03671_);
  nor (_03674_, _03671_, rst);
  nand (_03675_, _03670_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03677_, _03670_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03678_, _03677_, _03675_);
  and (_27319_[3], _03678_, _03674_);
  and (_03679_, _00144_, _26838_);
  and (_03680_, _03679_, _00106_);
  nor (_03681_, _00029_, _00067_);
  and (_03682_, _03681_, _03680_);
  and (_03683_, _03682_, _00296_);
  nor (_03684_, _03683_, _00152_);
  nor (_03685_, _00196_, _00176_);
  and (_03686_, _03685_, _02618_);
  or (_03687_, _03686_, _00214_);
  and (_03688_, _00196_, _00176_);
  and (_03690_, _03688_, _02640_);
  not (_03691_, _00196_);
  and (_03692_, _03691_, _00176_);
  and (_03694_, _03692_, _02629_);
  nor (_03695_, _03691_, _00176_);
  and (_03696_, _03695_, _02610_);
  or (_03697_, _03696_, _03694_);
  or (_03698_, _03697_, _03690_);
  or (_03699_, _03698_, _03687_);
  not (_03700_, _00214_);
  and (_03701_, _03685_, _02651_);
  or (_03702_, _03701_, _03700_);
  and (_03703_, _03688_, _24763_);
  and (_03704_, _03692_, _02671_);
  and (_03705_, _03695_, _23709_);
  or (_03706_, _03705_, _03704_);
  or (_03707_, _03706_, _03703_);
  or (_03708_, _03707_, _03702_);
  nand (_03709_, _03708_, _03699_);
  nor (_03710_, _03709_, _03684_);
  not (_03711_, _00067_);
  and (_03712_, _00029_, _03711_);
  not (_03713_, _00144_);
  and (_03714_, _00106_, _26838_);
  and (_03715_, _03714_, _03713_);
  and (_03716_, _03715_, _03712_);
  not (_03717_, _00299_);
  nand (_03718_, _03717_, _26568_);
  nor (_03719_, _24713_, _23275_);
  nor (_03720_, _03719_, _02549_);
  and (_03721_, _00303_, _00300_);
  not (_03722_, _03721_);
  nor (_03723_, _03722_, _03720_);
  and (_03724_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03725_, _03724_, _00292_);
  nor (_03726_, _03725_, _03723_);
  nand (_03727_, _03726_, _03718_);
  and (_03728_, _00950_, _00292_);
  not (_03729_, _03728_);
  and (_03730_, _03729_, _03727_);
  nand (_03731_, _00408_, _03717_);
  nor (_03732_, _23878_, _23245_);
  nor (_03733_, _03732_, _02533_);
  nor (_03734_, _03733_, _03722_);
  and (_03735_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03736_, _03735_, _00292_);
  nor (_03737_, _03736_, _03734_);
  nand (_03738_, _03737_, _03731_);
  and (_03740_, _01011_, _00292_);
  not (_03742_, _03740_);
  and (_03743_, _03742_, _03738_);
  or (_03744_, _03743_, _03730_);
  nand (_03745_, _03743_, _03730_);
  nand (_03746_, _03745_, _03744_);
  nand (_03747_, _00484_, _03717_);
  nor (_03749_, _23992_, _23214_);
  nor (_03750_, _03749_, _02509_);
  nor (_03752_, _03750_, _03722_);
  and (_03753_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03754_, _03753_, _00292_);
  nor (_03755_, _03754_, _03752_);
  nand (_03756_, _03755_, _03747_);
  and (_03757_, _01071_, _00292_);
  not (_03758_, _03757_);
  nand (_03759_, _03758_, _03756_);
  nand (_03760_, _00580_, _03717_);
  nor (_03761_, _23925_, _23181_);
  nor (_03763_, _03761_, _24635_);
  nor (_03764_, _03763_, _03722_);
  and (_03766_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_03767_, _03766_, _03764_);
  and (_03769_, _03767_, _00293_);
  and (_03770_, _03769_, _03760_);
  and (_03772_, _01138_, _00292_);
  nor (_03773_, _03772_, _03770_);
  nand (_03774_, _03773_, _03759_);
  or (_03775_, _03773_, _03759_);
  and (_03776_, _03775_, _03774_);
  nand (_03777_, _03776_, _03746_);
  or (_03778_, _03776_, _03746_);
  nand (_03779_, _03778_, _03777_);
  and (_03780_, _00647_, _03717_);
  nor (_03781_, _23986_, _23149_);
  or (_03782_, _03781_, _24732_);
  and (_03783_, _03782_, _03721_);
  and (_03785_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03787_, _03785_, _00292_);
  or (_03789_, _03787_, _03783_);
  or (_03790_, _03789_, _03780_);
  or (_03791_, _01228_, _00293_);
  and (_03792_, _03791_, _03790_);
  and (_03793_, _00708_, _03717_);
  nand (_03794_, _23919_, _23522_);
  or (_03795_, _23919_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03796_, _03795_, _03721_);
  and (_03797_, _03796_, _03794_);
  and (_03798_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03799_, _03798_, _00292_);
  or (_03800_, _03799_, _03797_);
  or (_03801_, _03800_, _03793_);
  or (_03802_, _01300_, _00293_);
  and (_03803_, _03802_, _03801_);
  or (_03804_, _03803_, _03792_);
  nand (_03805_, _03803_, _03792_);
  nand (_03806_, _03805_, _03804_);
  or (_03808_, _00791_, _00299_);
  not (_03809_, _24688_);
  nor (_03810_, _03809_, _23522_);
  nor (_03811_, _24688_, _23369_);
  nor (_03812_, _03811_, _03810_);
  nor (_03814_, _03812_, _03722_);
  and (_03816_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03817_, _03816_, _00292_);
  nor (_03819_, _03817_, _03814_);
  and (_03821_, _03819_, _03808_);
  and (_03822_, _01377_, _00292_);
  or (_03823_, _03822_, _03821_);
  and (_03824_, _00874_, _03717_);
  not (_03825_, _24671_);
  nor (_03826_, _03825_, _23522_);
  nor (_03827_, _24671_, _23084_);
  or (_03828_, _03827_, _03826_);
  and (_03829_, _03828_, _03721_);
  and (_03830_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03831_, _03830_, _00292_);
  or (_03832_, _03831_, _03829_);
  or (_03833_, _03832_, _03824_);
  nor (_03834_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_03836_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_03837_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _03836_);
  nor (_03838_, _03837_, _03834_);
  nor (_03839_, _03838_, _01335_);
  and (_03840_, _03838_, _01335_);
  or (_03841_, _03840_, _03839_);
  and (_03843_, _03841_, _23037_);
  or (_03844_, _26524_, _26484_);
  and (_03846_, _03844_, _26526_);
  and (_03847_, _03846_, _23531_);
  and (_03848_, _01280_, _23404_);
  and (_03849_, _03848_, _23373_);
  nor (_03850_, _03849_, _01352_);
  or (_03852_, _03850_, _01362_);
  nand (_03853_, _03852_, _23090_);
  or (_03854_, _03852_, _23090_);
  and (_03855_, _03854_, _23543_);
  and (_03857_, _03855_, _03853_);
  and (_03858_, _23468_, _23401_);
  or (_03859_, _03858_, _00930_);
  and (_03860_, _03859_, _23568_);
  and (_03861_, _23509_, _23552_);
  nor (_03862_, _26552_, _23090_);
  and (_03863_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or (_03864_, _03863_, _03862_);
  or (_03865_, _03864_, _03861_);
  or (_03866_, _03865_, _03860_);
  or (_03867_, _03866_, _03857_);
  or (_03868_, _03867_, _03847_);
  or (_03869_, _03868_, _03843_);
  or (_03871_, _03869_, _00293_);
  and (_03872_, _03871_, _03833_);
  or (_03874_, _03872_, _03823_);
  nand (_03875_, _03872_, _03823_);
  and (_03876_, _03875_, _03874_);
  nand (_03877_, _03876_, _03806_);
  or (_03878_, _03876_, _03806_);
  nand (_03879_, _03878_, _03877_);
  nand (_03880_, _03879_, _03779_);
  or (_03881_, _03879_, _03779_);
  nand (_03882_, _03881_, _03880_);
  nand (_03883_, _03882_, _00214_);
  or (_03884_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03885_, _03884_, _03688_);
  and (_03886_, _03885_, _03883_);
  and (_03887_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03888_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03889_, _03888_, _03887_);
  and (_03890_, _03889_, _03700_);
  nor (_03891_, _00214_, _00569_);
  and (_03892_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03893_, _03892_, _03891_);
  and (_03894_, _03893_, _03695_);
  and (_03895_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03896_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03897_, _03896_, _03895_);
  and (_03898_, _03897_, _00214_);
  or (_03899_, _03898_, _03894_);
  or (_03900_, _03899_, _03890_);
  or (_03901_, _03900_, _03886_);
  and (_03902_, _03901_, _03716_);
  and (_03903_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_03905_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03907_, _03905_, _03903_);
  and (_03908_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03909_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03910_, _03909_, _03908_);
  or (_03911_, _03910_, _03907_);
  and (_03912_, _03911_, _00214_);
  and (_03914_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03915_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03916_, _03915_, _03914_);
  and (_03917_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03918_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03919_, _03918_, _03917_);
  or (_03920_, _03919_, _03916_);
  and (_03921_, _03920_, _03700_);
  or (_03922_, _03921_, _03912_);
  and (_03923_, _03922_, _03680_);
  and (_03924_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03925_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_03927_, _03925_, _03924_);
  and (_03928_, _03927_, _03688_);
  and (_03929_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03930_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03931_, _03930_, _03929_);
  and (_03932_, _03931_, _03685_);
  or (_03934_, _03932_, _03928_);
  and (_03935_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03937_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03938_, _03937_, _03935_);
  and (_03939_, _03938_, _03695_);
  and (_03940_, _03700_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_03941_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03942_, _03941_, _03940_);
  and (_03943_, _03942_, _03692_);
  or (_03944_, _03943_, _03939_);
  or (_03945_, _03944_, _03934_);
  and (_03946_, _03945_, _03715_);
  or (_03947_, _03946_, _03923_);
  and (_03949_, _03947_, _03681_);
  nor (_03950_, _00144_, _00106_);
  and (_03951_, _03950_, _26838_);
  not (_03952_, _00029_);
  and (_03954_, _03952_, _00067_);
  and (_03955_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_03956_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_03958_, _03956_, _03955_);
  and (_03960_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_03961_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03963_, _03961_, _03960_);
  or (_03964_, _03963_, _03958_);
  and (_03965_, _03964_, _03954_);
  and (_03966_, _00029_, _00067_);
  and (_03967_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_03968_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03969_, _03968_, _03967_);
  and (_03971_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_03972_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03973_, _03972_, _03971_);
  or (_03974_, _03973_, _03969_);
  and (_03975_, _03974_, _03966_);
  or (_03976_, _03975_, _03965_);
  and (_03977_, _03976_, _00214_);
  and (_03978_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03979_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_03980_, _03979_, _03978_);
  and (_03981_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03982_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_03983_, _03982_, _03981_);
  or (_03984_, _03983_, _03980_);
  and (_03985_, _03984_, _03954_);
  and (_03986_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_03987_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_03988_, _03987_, _03986_);
  and (_03989_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_03990_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_03991_, _03990_, _03989_);
  or (_03992_, _03991_, _03988_);
  and (_03993_, _03992_, _03966_);
  or (_03994_, _03993_, _03985_);
  and (_03996_, _03994_, _03700_);
  or (_03997_, _03996_, _03977_);
  and (_03998_, _03997_, _03951_);
  or (_04000_, _03998_, _03949_);
  and (_04001_, _00220_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not (_04002_, _00106_);
  and (_04003_, _03679_, _04002_);
  and (_04004_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_04005_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_04006_, _04005_, _04004_);
  and (_04007_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04009_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_04010_, _04009_, _04007_);
  or (_04011_, _04010_, _04006_);
  and (_04012_, _04011_, _00214_);
  and (_04013_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_04014_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_04015_, _04014_, _04013_);
  and (_04016_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04017_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_04018_, _04017_, _04016_);
  or (_04019_, _04018_, _04015_);
  and (_04020_, _04019_, _03700_);
  or (_04022_, _04020_, _04012_);
  and (_04023_, _04022_, _03954_);
  and (_04025_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_04026_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_04027_, _04026_, _04025_);
  and (_04028_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_04030_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_04031_, _04030_, _04028_);
  or (_04033_, _04031_, _04027_);
  and (_04034_, _04033_, _00214_);
  and (_04035_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_04036_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_04037_, _04036_, _04035_);
  and (_04039_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_04040_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_04042_, _04040_, _04039_);
  or (_04043_, _04042_, _04037_);
  and (_04045_, _04043_, _03700_);
  or (_04046_, _04045_, _04034_);
  and (_04048_, _04046_, _03966_);
  or (_04049_, _04048_, _04023_);
  and (_04051_, _04049_, _04003_);
  or (_04052_, _04051_, _04001_);
  or (_04054_, _04052_, _04000_);
  not (_04055_, _26658_);
  not (_04056_, _01997_);
  and (_04057_, _24474_, _24451_);
  nor (_04059_, _04057_, _01996_);
  and (_04061_, _04059_, _04056_);
  and (_04062_, _04061_, _04055_);
  and (_04064_, _04062_, _26705_);
  not (_04065_, _26739_);
  and (_04066_, _04065_, _26708_);
  and (_04067_, _04066_, _04064_);
  and (_04068_, _24466_, _24460_);
  not (_04069_, _04068_);
  and (_04070_, _26577_, _24517_);
  and (_04071_, _24466_, _24453_);
  nor (_04072_, _04071_, _04070_);
  and (_04073_, _04072_, _04069_);
  and (_04074_, _04073_, _02008_);
  and (_04075_, _04074_, _04067_);
  and (_04076_, _04075_, _26700_);
  nor (_04077_, _04076_, _26576_);
  or (_04078_, _04077_, p0_in[1]);
  not (_04079_, _04077_);
  or (_04080_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_04081_, _04080_, _04078_);
  and (_04083_, _04081_, _03692_);
  or (_04085_, _04077_, p0_in[3]);
  or (_04086_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_04088_, _04086_, _04085_);
  and (_04089_, _04088_, _03685_);
  or (_04091_, _04089_, _04083_);
  nor (_04092_, _04077_, p0_in[0]);
  and (_04093_, _04077_, _25445_);
  nor (_04095_, _04093_, _04092_);
  and (_04096_, _04095_, _03688_);
  or (_04097_, _04077_, p0_in[2]);
  or (_04098_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_04100_, _04098_, _04097_);
  and (_04101_, _04100_, _03695_);
  or (_04103_, _04101_, _04096_);
  or (_04104_, _04103_, _04091_);
  and (_04105_, _04104_, _03680_);
  or (_04106_, _04077_, p1_in[3]);
  or (_04107_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_04108_, _04107_, _04106_);
  and (_04109_, _04108_, _03685_);
  or (_04111_, _04077_, p1_in[1]);
  or (_04112_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_04114_, _04112_, _04111_);
  and (_04115_, _04114_, _03692_);
  or (_04116_, _04115_, _04109_);
  or (_04118_, _04077_, p1_in[2]);
  or (_04119_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_04121_, _04119_, _04118_);
  and (_04122_, _04121_, _03695_);
  nor (_04123_, _04077_, p1_in[0]);
  and (_04124_, _04077_, _25364_);
  nor (_04126_, _04124_, _04123_);
  and (_04128_, _04126_, _03688_);
  or (_04129_, _04128_, _04122_);
  or (_04130_, _04129_, _04116_);
  and (_04131_, _04130_, _03715_);
  or (_04132_, _04131_, _04105_);
  and (_04134_, _04132_, _00214_);
  or (_04136_, _04077_, p1_in[6]);
  or (_04138_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_04139_, _04138_, _04136_);
  and (_04140_, _04139_, _03695_);
  or (_04141_, _04077_, p1_in[4]);
  or (_04142_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_04143_, _04142_, _04141_);
  and (_04145_, _04143_, _03688_);
  or (_04146_, _04145_, _04140_);
  or (_04147_, _04077_, p1_in[7]);
  or (_04148_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_04149_, _04148_, _04147_);
  and (_04150_, _04149_, _03685_);
  or (_04151_, _04077_, p1_in[5]);
  or (_04152_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_04153_, _04152_, _04151_);
  and (_04154_, _04153_, _03692_);
  or (_04155_, _04154_, _04150_);
  or (_04156_, _04155_, _04146_);
  and (_04157_, _04156_, _03715_);
  or (_04158_, _04077_, p0_in[5]);
  or (_04159_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_04160_, _04159_, _04158_);
  and (_04161_, _04160_, _03692_);
  or (_04162_, _04077_, p0_in[7]);
  or (_04163_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_04165_, _04163_, _04162_);
  and (_04166_, _04165_, _03685_);
  or (_04167_, _04166_, _04161_);
  or (_04168_, _04077_, p0_in[4]);
  or (_04169_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_04170_, _04169_, _04168_);
  and (_04171_, _04170_, _03688_);
  or (_04172_, _04077_, p0_in[6]);
  or (_04174_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_04175_, _04174_, _04172_);
  and (_04177_, _04175_, _03695_);
  or (_04178_, _04177_, _04171_);
  or (_04179_, _04178_, _04167_);
  and (_04180_, _04179_, _03680_);
  or (_04181_, _04180_, _04157_);
  and (_04182_, _04181_, _03700_);
  or (_04183_, _04182_, _04134_);
  and (_04184_, _04183_, _03966_);
  and (_04186_, _04003_, _03712_);
  nand (_04187_, _03712_, _00144_);
  nand (_04188_, _04187_, _03714_);
  and (_04190_, _26838_, _00067_);
  nand (_04191_, _04190_, _04002_);
  and (_04193_, _04191_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nand (_04194_, _04193_, _04188_);
  nor (_04195_, _04194_, _04186_);
  and (_04196_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_04197_, _04196_, _00214_);
  and (_04199_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04200_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_04202_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_04203_, _04202_, _04200_);
  or (_04204_, _04203_, _04199_);
  or (_04205_, _04204_, _04197_);
  and (_04206_, _03695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_04207_, _04206_, _03700_);
  and (_04208_, _03692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_04210_, _03688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_04211_, _03685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_04212_, _04211_, _04210_);
  or (_04214_, _04212_, _04208_);
  or (_04215_, _04214_, _04207_);
  and (_04216_, _04215_, _04205_);
  and (_04217_, _04216_, _04186_);
  or (_04219_, _04077_, p2_in[7]);
  or (_04220_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_04222_, _04220_, _04219_);
  and (_04223_, _04222_, _03700_);
  or (_04224_, _04077_, p2_in[3]);
  or (_04226_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_04227_, _04226_, _04224_);
  and (_04228_, _04227_, _00214_);
  or (_04229_, _04228_, _04223_);
  and (_04230_, _04229_, _03685_);
  or (_04231_, _04077_, p2_in[6]);
  or (_04232_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_04234_, _04232_, _04231_);
  and (_04235_, _04234_, _03700_);
  or (_04237_, _04077_, p2_in[2]);
  or (_04238_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_04239_, _04238_, _04237_);
  and (_04240_, _04239_, _00214_);
  or (_04241_, _04240_, _04235_);
  and (_04242_, _04241_, _03695_);
  or (_04243_, _04242_, _04230_);
  or (_04245_, _04077_, p2_in[4]);
  or (_04246_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_04247_, _04246_, _04245_);
  and (_04248_, _04247_, _03700_);
  nor (_04250_, _04077_, p2_in[0]);
  and (_04251_, _04077_, _25284_);
  nor (_04252_, _04251_, _04250_);
  and (_04253_, _04252_, _00214_);
  or (_04254_, _04253_, _04248_);
  and (_04255_, _04254_, _03688_);
  or (_04256_, _04077_, p2_in[5]);
  or (_04257_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_04258_, _04257_, _04256_);
  and (_04259_, _04258_, _03700_);
  or (_04260_, _04077_, p2_in[1]);
  or (_04261_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_04262_, _04261_, _04260_);
  and (_04263_, _04262_, _00214_);
  or (_04264_, _04263_, _04259_);
  and (_04265_, _04264_, _03692_);
  or (_04266_, _04265_, _04255_);
  or (_04267_, _04266_, _04243_);
  and (_04268_, _04267_, _03680_);
  or (_04269_, _04077_, p3_in[7]);
  or (_04270_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_04271_, _04270_, _04269_);
  and (_04272_, _04271_, _03700_);
  or (_04273_, _04077_, p3_in[3]);
  or (_04274_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_04276_, _04274_, _04273_);
  and (_04277_, _04276_, _00214_);
  or (_04278_, _04277_, _04272_);
  and (_04279_, _04278_, _03685_);
  or (_04280_, _04077_, p3_in[6]);
  or (_04282_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_04284_, _04282_, _04280_);
  and (_04285_, _04284_, _03700_);
  or (_04287_, _04077_, p3_in[2]);
  or (_04289_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_04290_, _04289_, _04287_);
  and (_04291_, _04290_, _00214_);
  or (_04293_, _04291_, _04285_);
  and (_04294_, _04293_, _03695_);
  or (_04295_, _04294_, _04279_);
  or (_04296_, _04077_, p3_in[4]);
  or (_04297_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_04299_, _04297_, _04296_);
  and (_04300_, _04299_, _03700_);
  nor (_04302_, _04077_, p3_in[0]);
  and (_04303_, _04077_, _25167_);
  nor (_04304_, _04303_, _04302_);
  and (_04305_, _04304_, _00214_);
  or (_04306_, _04305_, _04300_);
  and (_04308_, _04306_, _03688_);
  or (_04309_, _04077_, p3_in[5]);
  or (_04310_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_04312_, _04310_, _04309_);
  and (_04313_, _04312_, _03700_);
  or (_04314_, _04077_, p3_in[1]);
  or (_04315_, _04079_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_04316_, _04315_, _04314_);
  and (_04318_, _04316_, _00214_);
  or (_04319_, _04318_, _04313_);
  and (_04321_, _04319_, _03692_);
  or (_04323_, _04321_, _04308_);
  or (_04325_, _04323_, _04295_);
  and (_04326_, _04325_, _03715_);
  or (_04327_, _04326_, _04268_);
  and (_04329_, _04327_, _03954_);
  or (_04330_, _04329_, _04217_);
  or (_04332_, _04330_, _04195_);
  or (_04334_, _04332_, _04184_);
  or (_04335_, _04334_, _04054_);
  or (_04336_, _04335_, _03902_);
  nand (_04337_, _04001_, _23522_);
  and (_04338_, _04337_, _03684_);
  and (_04339_, _04338_, _04336_);
  or (_04340_, _04339_, _03710_);
  and (_27320_, _04340_, _22761_);
  and (_04341_, _00214_, _00106_);
  and (_04342_, _04341_, _03688_);
  and (_04343_, _03681_, _03679_);
  and (_04344_, _04343_, _04342_);
  and (_04345_, _04344_, _00296_);
  not (_04347_, _24706_);
  and (_04348_, _03685_, _03700_);
  nor (_04349_, _04348_, _04347_);
  and (_04350_, _04349_, _00150_);
  nor (_04351_, _04350_, _04345_);
  and (_04352_, _04351_, _00223_);
  and (_04353_, _00295_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_04355_, _03966_, _03679_);
  and (_04356_, _04355_, _03685_);
  and (_04357_, _04356_, _04341_);
  and (_04358_, _04357_, _04353_);
  not (_04359_, _04358_);
  not (_04360_, _26838_);
  nor (_04361_, _04360_, _00067_);
  and (_04362_, _00029_, _03713_);
  and (_04363_, _04362_, _04361_);
  and (_04364_, _04363_, _04342_);
  and (_04365_, _04364_, _00312_);
  and (_04366_, _04344_, _00292_);
  nor (_04367_, _04366_, _04365_);
  and (_04368_, _04367_, _04359_);
  nor (_04369_, _04368_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_04370_, _04369_);
  and (_04371_, _04370_, _04352_);
  and (_04372_, _04355_, _03695_);
  and (_04374_, _04372_, _04341_);
  and (_04375_, _04374_, _04353_);
  or (_04376_, _04375_, rst);
  nor (_27321_, _04376_, _04371_);
  nor (_04378_, _00029_, _00144_);
  and (_04379_, _04378_, _04361_);
  and (_04381_, _04379_, _04342_);
  nor (_04382_, _03700_, _00106_);
  and (_04383_, _04382_, _03688_);
  and (_04384_, _04362_, _04190_);
  and (_04385_, _04384_, _04383_);
  and (_04386_, _04355_, _03692_);
  and (_04387_, _04386_, _04341_);
  or (_04388_, _04387_, _04385_);
  nor (_04390_, _04388_, _04381_);
  and (_04391_, _04382_, _03685_);
  and (_04393_, _04391_, _04355_);
  and (_04394_, _04382_, _03692_);
  and (_04395_, _04394_, _04355_);
  nor (_04397_, _04395_, _04393_);
  and (_04398_, _04382_, _04372_);
  and (_04400_, _04348_, _00106_);
  and (_04401_, _04378_, _04190_);
  and (_04402_, _04401_, _04400_);
  nor (_04403_, _04402_, _04398_);
  and (_04405_, _04403_, _04397_);
  and (_04406_, _04405_, _04390_);
  or (_04407_, _04343_, _04190_);
  or (_04408_, _04407_, _04363_);
  nand (_04409_, _04408_, _04342_);
  nor (_04410_, _04374_, _04357_);
  and (_04411_, _03712_, _03679_);
  and (_04413_, _04411_, _04383_);
  nor (_04414_, _00214_, _00106_);
  and (_04415_, _04414_, _03692_);
  and (_04416_, _04415_, _04411_);
  and (_04418_, _04414_, _03688_);
  and (_04419_, _04418_, _04411_);
  or (_04421_, _04419_, _04416_);
  nor (_04422_, _04421_, _04413_);
  and (_04423_, _04422_, _04410_);
  and (_04424_, _04423_, _04409_);
  and (_04425_, _03954_, _03679_);
  and (_04426_, _04425_, _04383_);
  and (_04427_, _04382_, _03695_);
  and (_04428_, _04427_, _04411_);
  not (_04429_, _04428_);
  and (_04430_, _04383_, _04355_);
  and (_04432_, _04391_, _04411_);
  nor (_04433_, _04432_, _04430_);
  nand (_04434_, _04433_, _04429_);
  nor (_04435_, _04434_, _04426_);
  and (_04436_, _04418_, _04355_);
  and (_04437_, _04415_, _04355_);
  nor (_04439_, _04437_, _04436_);
  and (_04440_, _04394_, _04384_);
  and (_04442_, _04400_, _04355_);
  nor (_04443_, _04442_, _04440_);
  and (_04444_, _04443_, _04439_);
  and (_04446_, _04444_, _04435_);
  and (_04447_, _04446_, _04424_);
  and (_04448_, _04447_, _04406_);
  not (_04449_, _04448_);
  and (_04450_, _04449_, _04371_);
  not (_04451_, _04450_);
  and (_04452_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_04453_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_04454_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_04455_, _04454_, _04453_);
  and (_04456_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_04457_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_04458_, _04457_, _04456_);
  or (_04459_, _04458_, _04455_);
  and (_04460_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_04461_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_04463_, _04461_, _04460_);
  and (_04464_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_04465_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_04466_, _04465_, _04464_);
  or (_04467_, _04466_, _04463_);
  or (_04468_, _04467_, _04459_);
  and (_04469_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_04470_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_04472_, _04470_, _04469_);
  and (_04473_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_04474_, _04427_, _04355_);
  and (_04476_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_04477_, _04476_, _04473_);
  or (_04479_, _04477_, _04472_);
  and (_04480_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_04481_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_04483_, _04481_, _04480_);
  and (_04484_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_04486_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_04487_, _04486_, _04484_);
  or (_04488_, _04487_, _04483_);
  or (_04489_, _04488_, _04479_);
  or (_04491_, _04489_, _04468_);
  and (_04493_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_04494_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_04496_, _04494_, _04493_);
  and (_04497_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_04499_, _04341_, _03692_);
  and (_04500_, _04499_, _04355_);
  and (_04501_, _04500_, _26794_);
  or (_04502_, _04501_, _04497_);
  or (_04504_, _04502_, _04496_);
  and (_04505_, _04425_, _04342_);
  and (_04506_, _04505_, _04222_);
  and (_04507_, _04401_, _04342_);
  and (_04508_, _04507_, _04271_);
  or (_04509_, _04508_, _04506_);
  and (_04510_, _04355_, _04342_);
  and (_04511_, _04510_, _04165_);
  and (_04512_, _04384_, _04342_);
  and (_04513_, _04512_, _04149_);
  or (_04514_, _04513_, _04511_);
  or (_04515_, _04514_, _04509_);
  or (_04516_, _04515_, _04504_);
  and (_04517_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_04518_, _04364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_04519_, _04518_, _04517_);
  or (_04520_, _04519_, _04516_);
  or (_04521_, _04520_, _04491_);
  and (_04522_, _04521_, _04371_);
  or (_04524_, _04522_, _04375_);
  or (_04525_, _04524_, _04452_);
  not (_04526_, _04375_);
  or (_04527_, _04526_, _00874_);
  and (_04528_, _04527_, _22761_);
  and (_27322_[7], _04528_, _04525_);
  and (_04529_, _02785_, _23982_);
  and (_04530_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or (_25225_, _04530_, _04529_);
  and (_04532_, _02276_, _24078_);
  and (_04533_, _04532_, _23589_);
  not (_04535_, _04532_);
  and (_04537_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_25229_, _04537_, _04533_);
  and (_04538_, _03302_, _23589_);
  and (_04539_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or (_25232_, _04539_, _04538_);
  and (_04541_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_04542_, _03314_, _23635_);
  or (_25287_, _04542_, _04541_);
  and (_04544_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_04545_, _03314_, _23982_);
  or (_25293_, _04545_, _04544_);
  and (_04547_, _03340_, _23676_);
  and (_04549_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_27207_, _04549_, _04547_);
  and (_04551_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_04552_, _03314_, _23838_);
  or (_25300_, _04552_, _04551_);
  and (_04554_, _25742_, _23755_);
  and (_04556_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or (_27269_, _04556_, _04554_);
  and (_04557_, _03183_, _23962_);
  not (_04558_, _04557_);
  and (_04559_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  and (_04560_, _04557_, _23791_);
  or (_25318_, _04560_, _04559_);
  and (_04561_, _03648_, _23718_);
  and (_04562_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_25326_, _04562_, _04561_);
  and (_04563_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  and (_04564_, _04557_, _23838_);
  or (_25330_, _04564_, _04563_);
  and (_04565_, _03648_, _23791_);
  and (_04566_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_25347_, _04566_, _04565_);
  and (_04568_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and (_04569_, _04557_, _23718_);
  or (_25350_, _04569_, _04568_);
  and (_04570_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and (_04571_, _04557_, _23635_);
  or (_25393_, _04571_, _04570_);
  and (_04572_, _03648_, _23982_);
  and (_04573_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_25396_, _04573_, _04572_);
  and (_04576_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  and (_04578_, _04557_, _23589_);
  or (_25404_, _04578_, _04576_);
  and (_04579_, _03648_, _23838_);
  and (_04580_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_27112_, _04580_, _04579_);
  and (_04582_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  and (_04583_, _04557_, _23755_);
  or (_25421_, _04583_, _04582_);
  and (_04584_, _23652_, _23635_);
  and (_04585_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_25427_, _04585_, _04584_);
  or (_04587_, _03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_25439_, _04587_, _03395_);
  and (_04588_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  and (_04589_, _03184_, _23589_);
  or (_25460_, _04589_, _04588_);
  or (_04591_, _03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_25475_, _04591_, _03068_);
  and (_04592_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and (_04593_, _02762_, _23676_);
  or (_25480_, _04593_, _04592_);
  and (_04595_, _24615_, _23017_);
  not (_04596_, _04595_);
  and (_04597_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and (_04598_, _04595_, _23676_);
  or (_25490_, _04598_, _04597_);
  and (_04599_, _24615_, _23849_);
  not (_04601_, _04599_);
  and (_04602_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and (_04603_, _04599_, _23589_);
  or (_25500_, _04603_, _04602_);
  and (_04604_, _03376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_26923_, _04604_, _03379_);
  and (_04606_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_04608_, _04595_, _23838_);
  or (_25511_, _04608_, _04606_);
  or (_04609_, _03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_25514_, _04609_, _03388_);
  or (_04612_, _03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_26924_, _04612_, _03384_);
  and (_04613_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_04614_, _04595_, _23718_);
  or (_25524_, _04614_, _04613_);
  and (_04615_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_04617_, _04595_, _23791_);
  or (_25527_, _04617_, _04615_);
  and (_04619_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  and (_04621_, _04599_, _23718_);
  or (_25545_, _04621_, _04619_);
  not (_04622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_04623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not (_04624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_04625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_04626_, _04625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_04627_, _04626_, _04624_);
  nor (_04629_, _02594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04630_, _04629_, _04627_);
  nor (_04631_, _04630_, _04623_);
  nand (_04632_, _04631_, _04622_);
  nor (_04633_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_04634_, _04633_, _04631_);
  nand (_04635_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_04636_, _04635_, _04634_);
  and (_04637_, _04636_, _22761_);
  and (_25557_, _04637_, _04632_);
  not (_04638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and (_04639_, _02586_, _04638_);
  and (_04640_, _04639_, _02695_);
  and (_04641_, _04640_, _02692_);
  nand (_04642_, _04641_, _02581_);
  not (_04643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_04644_, _02697_, _04643_);
  and (_04645_, _04644_, _04642_);
  or (_04646_, _04645_, _02592_);
  and (_25560_, _04646_, _22761_);
  and (_25563_, _04634_, _22761_);
  and (_04649_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  and (_04650_, _04599_, _23635_);
  or (_25567_, _04650_, _04649_);
  and (_04651_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  and (_04652_, _04599_, _23982_);
  or (_25623_, _04652_, _04651_);
  and (_04653_, _02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or (_04654_, _04653_, _02592_);
  and (_04655_, _02592_, _02594_);
  nor (_04656_, _04655_, rst);
  and (_25624_, _04656_, _04654_);
  nand (_04657_, _02837_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or (_04658_, _02837_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_04659_, _04658_, _22761_);
  nand (_04660_, _04659_, _04657_);
  nor (_25626_, _04660_, _02592_);
  not (_04661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_04662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_04663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04664_, _04626_, _04663_);
  or (_04665_, _04664_, _04629_);
  nor (_04667_, _04665_, _04662_);
  nand (_04668_, _04667_, _04661_);
  nor (_04670_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_04671_, _04670_, _04667_);
  nand (_04672_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_04673_, _04672_, _04671_);
  and (_04674_, _04673_, _22761_);
  and (_25645_, _04674_, _04668_);
  and (_25649_, _04671_, _22761_);
  not (_04675_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_04676_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _02485_);
  not (_04677_, _04676_);
  nor (_04678_, _02516_, _02728_);
  and (_04679_, _04678_, _04677_);
  and (_04681_, _04679_, _02738_);
  nor (_04682_, _04681_, _04675_);
  and (_04683_, _04681_, rxd_i);
  or (_04684_, _04683_, rst);
  or (_25684_, _04684_, _04682_);
  or (_04686_, _02724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_04687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_04688_, _04687_, _02516_);
  or (_04689_, _04688_, _02705_);
  nand (_04690_, _04689_, _04686_);
  nand (_25686_, _04690_, _02100_);
  and (_04692_, _24541_, _23599_);
  and (_04693_, _04692_, _23982_);
  not (_04695_, _04692_);
  and (_04696_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_25698_, _04696_, _04693_);
  and (_04698_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_04699_, _04595_, _23755_);
  or (_25714_, _04699_, _04698_);
  and (_04700_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and (_04701_, _04595_, _23635_);
  or (_25719_, _04701_, _04700_);
  and (_04702_, _24080_, _23676_);
  and (_04703_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_25726_, _04703_, _04702_);
  and (_04704_, _24572_, _23962_);
  and (_04705_, _04704_, _23755_);
  not (_04706_, _04704_);
  and (_04707_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or (_25737_, _04707_, _04705_);
  and (_04708_, _24777_, _23755_);
  and (_04709_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or (_25747_, _04709_, _04708_);
  and (_04710_, _02862_, _23791_);
  and (_04711_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_25757_, _04711_, _04710_);
  and (_04712_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_04713_, _03255_, _23676_);
  or (_27123_, _04713_, _04712_);
  and (_04714_, _02342_, _23676_);
  and (_04715_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_25831_, _04715_, _04714_);
  and (_04717_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_04718_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_04719_, _22770_, _04718_);
  or (_04720_, _04719_, _04717_);
  and (_26891_[15], _04720_, _22761_);
  or (_04722_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand (_04724_, _22770_, _04718_);
  and (_04726_, _04724_, _22761_);
  and (_26892_[15], _04726_, _04722_);
  and (_04727_, _24769_, _23791_);
  and (_04728_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or (_25851_, _04728_, _04727_);
  and (_04730_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_04731_, _03255_, _23791_);
  or (_25854_, _04731_, _04730_);
  and (_04733_, _23650_, _23642_);
  and (_04734_, _04733_, _23842_);
  not (_04735_, _04734_);
  and (_04736_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  and (_04737_, _04734_, _23838_);
  or (_25884_, _04737_, _04736_);
  nand (_04739_, _02077_, _23585_);
  not (_04740_, _02073_);
  and (_04741_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_04742_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_04743_, _04742_, _04741_);
  or (_04744_, _04743_, _02077_);
  and (_04746_, _04744_, _04740_);
  and (_04747_, _04746_, _04739_);
  and (_04749_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_04750_, _04749_, _04747_);
  and (_25886_, _04750_, _22761_);
  and (_04751_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  and (_04752_, _04734_, _23718_);
  or (_25894_, _04752_, _04751_);
  and (_04753_, _04692_, _23755_);
  and (_04754_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_25912_, _04754_, _04753_);
  and (_04756_, _24558_, _24078_);
  not (_04757_, _04756_);
  and (_04758_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_04759_, _04756_, _23589_);
  or (_25919_, _04759_, _04758_);
  and (_04761_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_04763_, _04756_, _23676_);
  or (_27040_, _04763_, _04761_);
  and (_04764_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_04765_, _04756_, _23791_);
  or (_25931_, _04765_, _04764_);
  and (_04766_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_04767_, _04756_, _23838_);
  or (_27041_, _04767_, _04766_);
  and (_04769_, _03354_, _23718_);
  and (_04771_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_25939_, _04771_, _04769_);
  and (_04772_, _02277_, _23838_);
  and (_04773_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or (_25944_, _04773_, _04772_);
  and (_04774_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_04775_, _04756_, _23982_);
  or (_25947_, _04775_, _04774_);
  and (_04776_, _04733_, _23803_);
  not (_04777_, _04776_);
  and (_04778_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_04779_, _04776_, _23982_);
  or (_25951_, _04779_, _04778_);
  and (_04780_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_04781_, _04776_, _23635_);
  or (_25954_, _04781_, _04780_);
  and (_04783_, _02277_, _23791_);
  and (_04785_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  or (_25957_, _04785_, _04783_);
  and (_04786_, _02277_, _23589_);
  and (_04787_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or (_25962_, _04787_, _04786_);
  and (_04789_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_04790_, _04776_, _23589_);
  or (_27034_, _04790_, _04789_);
  and (_04792_, _04733_, _23849_);
  not (_04793_, _04792_);
  and (_04794_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_04795_, _04792_, _23676_);
  or (_25969_, _04795_, _04794_);
  and (_04796_, _03354_, _23982_);
  and (_04797_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_25973_, _04797_, _04796_);
  and (_04798_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_04799_, _04792_, _23838_);
  or (_25982_, _04799_, _04798_);
  and (_04800_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_04801_, _04792_, _23982_);
  or (_25992_, _04801_, _04800_);
  and (_04802_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_04803_, _04792_, _23755_);
  or (_25998_, _04803_, _04802_);
  and (_04804_, _03302_, _23791_);
  and (_04805_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or (_26007_, _04805_, _04804_);
  and (_04807_, _03302_, _23635_);
  and (_04808_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  or (_26009_, _04808_, _04807_);
  and (_04810_, _04733_, _23017_);
  not (_04811_, _04810_);
  and (_04812_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and (_04813_, _04810_, _23718_);
  or (_26012_, _04813_, _04812_);
  and (_04814_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  and (_04815_, _04810_, _23838_);
  or (_27035_, _04815_, _04814_);
  nor (_27319_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_04816_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_04817_, _03670_, rst);
  and (_27319_[1], _04817_, _04816_);
  nor (_04818_, _03670_, _03669_);
  or (_04819_, _04818_, _03671_);
  and (_04820_, _03675_, _22761_);
  and (_27319_[2], _04820_, _04819_);
  and (_04822_, _03302_, _23982_);
  and (_04823_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or (_26031_, _04823_, _04822_);
  not (_04824_, _04371_);
  nand (_04825_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_04826_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_04827_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_04828_, _04827_, _04826_);
  and (_04829_, _04828_, _04825_);
  nand (_04830_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_04831_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_04832_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_04833_, _04832_, _04831_);
  and (_04834_, _04833_, _04830_);
  and (_04835_, _04834_, _04829_);
  nand (_04836_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_04837_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_04838_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_04839_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_04840_, _04839_, _04838_);
  and (_04841_, _04840_, _04837_);
  and (_04842_, _04841_, _04836_);
  nand (_04843_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand (_04844_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_04845_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_04846_, _04845_, _04844_);
  and (_04847_, _04846_, _04843_);
  nand (_04848_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_04849_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_04850_, _04849_, _04848_);
  and (_04851_, _04850_, _04847_);
  nand (_04852_, _04510_, _04095_);
  nand (_04853_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nand (_04854_, _04512_, _04126_);
  and (_04855_, _04854_, _04853_);
  and (_04856_, _04855_, _04852_);
  nand (_04857_, _04387_, _00188_);
  nand (_04858_, _04505_, _04252_);
  nand (_04859_, _04507_, _04304_);
  and (_04860_, _04859_, _04858_);
  and (_04861_, _04860_, _04857_);
  and (_04863_, _04861_, _04856_);
  and (_04864_, _04863_, _04851_);
  and (_04865_, _04864_, _04842_);
  and (_04866_, _04865_, _04835_);
  not (_04867_, _04364_);
  or (_04868_, _04867_, _03882_);
  nand (_04869_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand (_04870_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_04871_, _04870_, _04869_);
  nand (_04873_, _04398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_04874_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_04875_, _04874_, _04873_);
  and (_04876_, _04875_, _04871_);
  and (_04878_, _04876_, _04868_);
  and (_04879_, _04878_, _04866_);
  nor (_04880_, _04879_, _04824_);
  nand (_04881_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_04882_, _04881_, _04526_);
  or (_04883_, _04882_, _04880_);
  or (_04884_, _04526_, _26568_);
  and (_04886_, _04884_, _22761_);
  and (_27322_[0], _04886_, _04883_);
  and (_04887_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_04888_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_04889_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_04890_, _04889_, _04888_);
  and (_04892_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_04893_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_04894_, _04893_, _04892_);
  or (_04895_, _04894_, _04890_);
  and (_04896_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04897_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_04898_, _04897_, _04896_);
  and (_04899_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_04901_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_04902_, _04901_, _04899_);
  or (_04904_, _04902_, _04898_);
  or (_04905_, _04904_, _04895_);
  and (_04906_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_04907_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_04908_, _04907_, _04906_);
  and (_04909_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_04910_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_04911_, _04910_, _04909_);
  or (_04912_, _04911_, _04908_);
  and (_04913_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_04915_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_04916_, _04915_, _04913_);
  and (_04917_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_04918_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_04919_, _04918_, _04917_);
  or (_04920_, _04919_, _04916_);
  or (_04921_, _04920_, _04912_);
  or (_04922_, _04921_, _04905_);
  and (_04923_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_04924_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_04925_, _04924_, _04923_);
  and (_04926_, _04387_, _00170_);
  and (_04928_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_04929_, _04928_, _04926_);
  or (_04930_, _04929_, _04925_);
  and (_04931_, _04512_, _04114_);
  and (_04932_, _04510_, _04081_);
  or (_04933_, _04932_, _04931_);
  and (_04935_, _04505_, _04262_);
  and (_04936_, _04507_, _04316_);
  or (_04937_, _04936_, _04935_);
  or (_04938_, _04937_, _04933_);
  or (_04939_, _04938_, _04930_);
  and (_04940_, _04364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_04942_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_04944_, _04942_, _04940_);
  or (_04945_, _04944_, _04939_);
  nor (_04946_, _04945_, _04922_);
  nor (_04947_, _04946_, _04824_);
  or (_04948_, _04947_, _04375_);
  or (_04949_, _04948_, _04887_);
  or (_04950_, _04526_, _00408_);
  and (_04951_, _04950_, _22761_);
  and (_27322_[1], _04951_, _04949_);
  and (_04952_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_04953_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_04954_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_04955_, _04954_, _04953_);
  and (_04956_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04957_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_04958_, _04957_, _04956_);
  or (_04959_, _04958_, _04955_);
  and (_04960_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_04961_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_04962_, _04961_, _04960_);
  and (_04963_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_04964_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_04965_, _04964_, _04963_);
  or (_04966_, _04965_, _04962_);
  or (_04967_, _04966_, _04959_);
  and (_04968_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_04969_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_04970_, _04969_, _04968_);
  and (_04971_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_04972_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_04973_, _04972_, _04971_);
  or (_04974_, _04973_, _04970_);
  and (_04975_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_04976_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_04977_, _04976_, _04975_);
  and (_04978_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_04979_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_04980_, _04979_, _04978_);
  or (_04981_, _04980_, _04977_);
  or (_04983_, _04981_, _04974_);
  or (_04984_, _04983_, _04967_);
  and (_04985_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_04987_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_04988_, _04987_, _04985_);
  and (_04989_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_04990_, _04500_, _00211_);
  or (_04992_, _04990_, _04989_);
  or (_04993_, _04992_, _04988_);
  and (_04994_, _04505_, _04239_);
  and (_04995_, _04507_, _04290_);
  or (_04996_, _04995_, _04994_);
  and (_04998_, _04510_, _04100_);
  and (_05000_, _04512_, _04121_);
  or (_05001_, _05000_, _04998_);
  or (_05002_, _05001_, _04996_);
  or (_05004_, _05002_, _04993_);
  and (_05005_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_05006_, _04364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_05007_, _05006_, _05005_);
  or (_05008_, _05007_, _05004_);
  or (_05009_, _05008_, _04984_);
  and (_05010_, _05009_, _04371_);
  or (_05011_, _05010_, _04375_);
  or (_05012_, _05011_, _04952_);
  or (_05013_, _04526_, _00484_);
  and (_05014_, _05013_, _22761_);
  and (_27322_[2], _05014_, _05012_);
  and (_05016_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_05017_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_05018_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_05019_, _05018_, _05017_);
  and (_05020_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_05021_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_05022_, _05021_, _05020_);
  or (_05023_, _05022_, _05019_);
  and (_05025_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_05026_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_05027_, _05026_, _05025_);
  and (_05028_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_05029_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_05030_, _05029_, _05028_);
  or (_05031_, _05030_, _05027_);
  or (_05032_, _05031_, _05023_);
  and (_05034_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_05035_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_05037_, _05035_, _05034_);
  and (_05038_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_05039_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_05040_, _05039_, _05038_);
  or (_05042_, _05040_, _05037_);
  and (_05043_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_05044_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_05045_, _05044_, _05043_);
  and (_05046_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_05047_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_05048_, _05047_, _05046_);
  or (_05049_, _05048_, _05045_);
  or (_05050_, _05049_, _05042_);
  or (_05051_, _05050_, _05032_);
  and (_05052_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_05054_, _04364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_05055_, _05054_, _05052_);
  and (_05056_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_05057_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_05058_, _05057_, _05056_);
  and (_05059_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_05060_, _04500_, _00099_);
  or (_05061_, _05060_, _05059_);
  or (_05062_, _05061_, _05058_);
  and (_05063_, _04505_, _04227_);
  and (_05064_, _04507_, _04276_);
  or (_05065_, _05064_, _05063_);
  and (_05066_, _04512_, _04108_);
  and (_05067_, _04510_, _04088_);
  or (_05068_, _05067_, _05066_);
  or (_05069_, _05068_, _05065_);
  or (_05070_, _05069_, _05062_);
  or (_05072_, _05070_, _05055_);
  or (_05073_, _05072_, _05051_);
  and (_05074_, _05073_, _04371_);
  or (_05076_, _05074_, _04375_);
  or (_05077_, _05076_, _05016_);
  or (_05078_, _04526_, _00580_);
  and (_05079_, _05078_, _22761_);
  and (_27322_[3], _05079_, _05077_);
  and (_05080_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_05081_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_05082_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_05083_, _05082_, _05081_);
  and (_05084_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_05085_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_05087_, _05085_, _05084_);
  or (_05088_, _05087_, _05083_);
  and (_05090_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_05091_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_05092_, _05091_, _05090_);
  and (_05093_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_05095_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_05096_, _05095_, _05093_);
  or (_05097_, _05096_, _05092_);
  or (_05099_, _05097_, _05088_);
  and (_05100_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_05101_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or (_05102_, _05101_, _05100_);
  and (_05103_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_05104_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_05105_, _05104_, _05103_);
  or (_05106_, _05105_, _05102_);
  and (_05108_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_05109_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_05110_, _05109_, _05108_);
  and (_05111_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_05113_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_05115_, _05113_, _05111_);
  or (_05117_, _05115_, _05110_);
  or (_05119_, _05117_, _05106_);
  or (_05120_, _05119_, _05099_);
  and (_05122_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_05123_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_05124_, _05123_, _05122_);
  and (_05125_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_05126_, _00116_);
  and (_05127_, _04500_, _05126_);
  or (_05128_, _05127_, _05125_);
  or (_05129_, _05128_, _05124_);
  and (_05130_, _04505_, _04247_);
  and (_05131_, _04507_, _04299_);
  or (_05133_, _05131_, _05130_);
  and (_05134_, _04512_, _04143_);
  and (_05135_, _04510_, _04170_);
  or (_05137_, _05135_, _05134_);
  or (_05138_, _05137_, _05133_);
  or (_05140_, _05138_, _05129_);
  and (_05141_, _04364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_05142_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_05143_, _05142_, _05141_);
  or (_05144_, _05143_, _05140_);
  or (_05145_, _05144_, _05120_);
  and (_05146_, _05145_, _04371_);
  or (_05147_, _05146_, _04375_);
  or (_05148_, _05147_, _05080_);
  or (_05149_, _04526_, _00647_);
  and (_05151_, _05149_, _22761_);
  and (_27322_[4], _05151_, _05148_);
  and (_05152_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_05153_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_05154_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_05155_, _05154_, _05153_);
  and (_05156_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_05157_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_05158_, _05157_, _05156_);
  or (_05159_, _05158_, _05155_);
  and (_05160_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_05161_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_05162_, _05161_, _05160_);
  and (_05163_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_05164_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_05165_, _05164_, _05163_);
  or (_05166_, _05165_, _05162_);
  or (_05167_, _05166_, _05159_);
  and (_05168_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_05169_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_05170_, _05169_, _05168_);
  and (_05171_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_05172_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_05173_, _05172_, _05171_);
  or (_05175_, _05173_, _05170_);
  and (_05176_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_05177_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_05178_, _05177_, _05176_);
  and (_05179_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_05180_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_05181_, _05180_, _05179_);
  or (_05182_, _05181_, _05178_);
  or (_05183_, _05182_, _05175_);
  or (_05184_, _05183_, _05167_);
  and (_05185_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_05186_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_05187_, _05186_, _05185_);
  and (_05188_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_05189_, _00001_);
  and (_05190_, _04500_, _05189_);
  or (_05191_, _05190_, _05188_);
  or (_05193_, _05191_, _05187_);
  and (_05194_, _04505_, _04258_);
  and (_05195_, _04507_, _04312_);
  or (_05196_, _05195_, _05194_);
  and (_05197_, _04512_, _04153_);
  and (_05198_, _04510_, _04160_);
  or (_05199_, _05198_, _05197_);
  or (_05200_, _05199_, _05196_);
  or (_05201_, _05200_, _05193_);
  and (_05202_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_05203_, _04364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_05204_, _05203_, _05202_);
  or (_05205_, _05204_, _05201_);
  or (_05206_, _05205_, _05184_);
  and (_05207_, _05206_, _04371_);
  or (_05208_, _05207_, _04375_);
  or (_05210_, _05208_, _05152_);
  or (_05211_, _04526_, _00708_);
  and (_05212_, _05211_, _22761_);
  and (_27322_[5], _05212_, _05210_);
  and (_05213_, _04451_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_05214_, _04416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_05215_, _04428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_05216_, _05215_, _05214_);
  and (_05217_, _04413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_05218_, _04419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_05219_, _05218_, _05217_);
  or (_05220_, _05219_, _05216_);
  and (_05221_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_05222_, _04402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_05223_, _05222_, _05221_);
  and (_05225_, _04432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_05226_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_05227_, _05226_, _05225_);
  or (_05228_, _05227_, _05223_);
  or (_05229_, _05228_, _05220_);
  and (_05230_, _04393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_05232_, _04395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or (_05234_, _05232_, _05230_);
  and (_05235_, _04437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_05236_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_05237_, _05236_, _05235_);
  or (_05238_, _05237_, _05234_);
  and (_05239_, _04440_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_05240_, _04385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_05241_, _05240_, _05239_);
  and (_05242_, _04442_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_05244_, _04436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_05245_, _05244_, _05242_);
  or (_05246_, _05245_, _05241_);
  or (_05247_, _05246_, _05238_);
  or (_05248_, _05247_, _05229_);
  and (_05249_, _04381_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_05250_, _00041_);
  and (_05251_, _04387_, _05250_);
  or (_05252_, _05251_, _05249_);
  and (_05253_, _04357_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_05254_, _04374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_05255_, _05254_, _05253_);
  or (_05256_, _05255_, _05252_);
  and (_05257_, _04510_, _04175_);
  and (_05258_, _04512_, _04139_);
  or (_05259_, _05258_, _05257_);
  and (_05260_, _04505_, _04234_);
  and (_05261_, _04507_, _04284_);
  or (_05262_, _05261_, _05260_);
  or (_05263_, _05262_, _05259_);
  or (_05264_, _05263_, _05256_);
  and (_05265_, _04364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_05266_, _04344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_05267_, _05266_, _05265_);
  or (_05268_, _05267_, _05264_);
  or (_05269_, _05268_, _05248_);
  and (_05270_, _05269_, _04371_);
  or (_05271_, _05270_, _04375_);
  or (_05272_, _05271_, _05213_);
  nand (_05273_, _04375_, _00791_);
  and (_05274_, _05273_, _22761_);
  and (_27322_[6], _05274_, _05272_);
  and (_05276_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  and (_05278_, _04810_, _23635_);
  or (_26043_, _05278_, _05276_);
  and (_05280_, _02379_, _23718_);
  and (_05281_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_26525_, _05281_, _05280_);
  and (_05282_, _04704_, _23838_);
  and (_05283_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or (_26527_, _05283_, _05282_);
  and (_05284_, _02862_, _23718_);
  and (_05286_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_27273_, _05286_, _05284_);
  and (_05287_, \oc8051_top_1.oc8051_sfr1.wait_data , _22761_);
  and (_05288_, _05287_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_05289_, _26656_, _24515_);
  or (_05290_, _05289_, _24391_);
  and (_05291_, _05290_, _00271_);
  and (_05292_, _24458_, _24515_);
  or (_05293_, _05292_, _26617_);
  or (_05294_, _24449_, _02243_);
  nor (_05295_, _05294_, _05293_);
  nand (_05296_, _05295_, _26715_);
  or (_05297_, _05296_, _02032_);
  or (_05298_, _05297_, _05291_);
  nor (_05299_, _26595_, _24517_);
  nor (_05300_, _05299_, _24417_);
  not (_05301_, _03053_);
  or (_05302_, _05301_, _02249_);
  or (_05303_, _05302_, _05300_);
  or (_05304_, _05303_, _02241_);
  and (_05305_, _26584_, _24321_);
  or (_05306_, _05305_, _26594_);
  and (_05307_, _24471_, _24486_);
  or (_05308_, _26725_, _05307_);
  or (_05309_, _03054_, _05308_);
  or (_05311_, _05309_, _02264_);
  or (_05312_, _05311_, _05306_);
  or (_05313_, _05312_, _05304_);
  or (_05314_, _05313_, _05298_);
  and (_05315_, _05314_, _25615_);
  or (_26879_[0], _05315_, _05288_);
  and (_05316_, _02862_, _23838_);
  and (_05317_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_26573_, _05317_, _05316_);
  and (_05318_, _02444_, _23718_);
  and (_05319_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_26586_, _05319_, _05318_);
  and (_05320_, _04704_, _23718_);
  and (_05321_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or (_26613_, _05321_, _05320_);
  and (_05322_, _23595_, _23027_);
  and (_05323_, _05322_, _24768_);
  and (_05324_, _05323_, _23718_);
  not (_05325_, _05323_);
  and (_05326_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or (_26649_, _05326_, _05324_);
  and (_05327_, _04704_, _23676_);
  and (_05328_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or (_26669_, _05328_, _05327_);
  and (_05329_, _24572_, _24078_);
  and (_05330_, _05329_, _23589_);
  not (_05331_, _05329_);
  and (_05332_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or (_26678_, _05332_, _05330_);
  and (_05333_, _05329_, _23982_);
  and (_05334_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or (_26684_, _05334_, _05333_);
  and (_05335_, _05329_, _23838_);
  and (_05336_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or (_26704_, _05336_, _05335_);
  and (_05338_, _05329_, _23791_);
  and (_05339_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or (_26734_, _05339_, _05338_);
  and (_05341_, _24542_, _23982_);
  and (_05342_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_26738_, _05342_, _05341_);
  and (_05343_, _24542_, _23838_);
  and (_05344_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_26763_, _05344_, _05343_);
  and (_05345_, _02937_, _23589_);
  and (_05346_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or (_26793_, _05346_, _05345_);
  and (_05347_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  and (_05348_, _04810_, _23589_);
  or (_26808_, _05348_, _05347_);
  nand (_05349_, _03066_, _04360_);
  or (_05350_, _05349_, _00144_);
  or (_05351_, _03066_, _00176_);
  nand (_05352_, _05351_, _05350_);
  and (_05353_, _05352_, _22967_);
  nor (_05354_, _05352_, _22967_);
  nor (_05355_, _05354_, _05353_);
  not (_05356_, _23024_);
  and (_05357_, _05349_, _03711_);
  nor (_05358_, _05357_, _05356_);
  and (_05359_, _05357_, _05356_);
  nor (_05360_, _05359_, _05358_);
  and (_05361_, _05349_, _03713_);
  nor (_05362_, _05361_, _23804_);
  and (_05363_, _05349_, _00029_);
  nor (_05364_, _05363_, _23021_);
  nor (_05365_, _05364_, _05362_);
  and (_05367_, _05365_, _05360_);
  and (_05368_, _05367_, _05355_);
  not (_05369_, _23014_);
  nor (_05371_, _05349_, _00029_);
  nor (_05372_, _03066_, _00214_);
  nor (_05373_, _05372_, _05371_);
  nor (_05374_, _05373_, _05369_);
  and (_05375_, _05373_, _05369_);
  nor (_05376_, _05375_, _05374_);
  and (_05377_, _05349_, _00106_);
  nor (_05378_, _05349_, _03711_);
  nor (_05379_, _05378_, _05377_);
  and (_05380_, _05379_, _22985_);
  nor (_05381_, _05379_, _22985_);
  or (_05382_, _05381_, _05380_);
  not (_05384_, _05382_);
  and (_05385_, _05384_, _05376_);
  or (_05386_, _05349_, _00106_);
  or (_05387_, _03066_, _00196_);
  nand (_05388_, _05387_, _05386_);
  and (_05389_, _05388_, _22928_);
  nor (_05390_, _05388_, _22928_);
  nor (_05391_, _05390_, _05389_);
  and (_05392_, _05363_, _23021_);
  not (_05393_, _05392_);
  nor (_05394_, _26841_, _22934_);
  not (_05395_, _05394_);
  and (_05396_, _05361_, _23804_);
  nor (_05397_, _05396_, _05395_);
  and (_05398_, _05397_, _05393_);
  and (_05399_, _05398_, _05391_);
  and (_05400_, _05399_, _05385_);
  and (_05401_, _05400_, _05368_);
  and (_26919_, _05401_, _22761_);
  and (_26920_[7], _23588_, _22761_);
  nor (_26922_[2], _00214_, rst);
  and (_05402_, _03015_, _23589_);
  and (_05403_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_00049_, _05403_, _05402_);
  and (_05404_, _03296_, _23982_);
  and (_05405_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_00051_, _05405_, _05404_);
  and (_05407_, _24558_, _23649_);
  not (_05408_, _05407_);
  and (_05409_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and (_05410_, _05407_, _23676_);
  or (_27039_, _05410_, _05409_);
  and (_05411_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  and (_05412_, _05407_, _23718_);
  or (_00071_, _05412_, _05411_);
  and (_05413_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and (_05414_, _05407_, _23982_);
  or (_00077_, _05414_, _05413_);
  and (_05415_, _03358_, _23791_);
  and (_05416_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or (_00079_, _05416_, _05415_);
  and (_05417_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  and (_05418_, _05407_, _23635_);
  or (_00085_, _05418_, _05417_);
  and (_05420_, _24558_, _23962_);
  not (_05421_, _05420_);
  and (_05423_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_05424_, _05420_, _23676_);
  or (_00134_, _05424_, _05423_);
  and (_05425_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_05426_, _05420_, _23718_);
  or (_00139_, _05426_, _05425_);
  and (_05427_, _03296_, _23589_);
  and (_05428_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_00142_, _05428_, _05427_);
  and (_05430_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_05431_, _05420_, _23982_);
  or (_27042_, _05431_, _05430_);
  and (_05433_, _03358_, _23635_);
  and (_05434_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or (_27169_, _05434_, _05433_);
  and (_05435_, _03358_, _23838_);
  and (_05436_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or (_00154_, _05436_, _05435_);
  and (_05437_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_05438_, _05420_, _23635_);
  or (_00157_, _05438_, _05437_);
  and (_05439_, _24558_, _23594_);
  not (_05440_, _05439_);
  and (_05441_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and (_05442_, _05439_, _23791_);
  or (_00162_, _05442_, _05441_);
  and (_05443_, _04692_, _23635_);
  and (_05444_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_00164_, _05444_, _05443_);
  and (_05445_, _02276_, _23649_);
  and (_05446_, _05445_, _23838_);
  not (_05447_, _05445_);
  and (_05448_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  or (_00167_, _05448_, _05446_);
  and (_26920_[0], _23674_, _22761_);
  and (_26920_[1], _23790_, _22761_);
  and (_26920_[2], _23717_, _22761_);
  and (_26920_[3], _23837_, _22761_);
  and (_26920_[4], _23981_, _22761_);
  and (_26920_[5], _23634_, _22761_);
  and (_26920_[6], _23754_, _22761_);
  and (_05449_, _05445_, _23589_);
  and (_05450_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or (_00243_, _05450_, _05449_);
  nor (_26922_[0], _00196_, rst);
  nor (_26922_[1], _00176_, rst);
  and (_05451_, _02937_, _23755_);
  and (_05452_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or (_00266_, _05452_, _05451_);
  nor (_05453_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_05454_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01853_);
  nor (_05455_, _05454_, _05453_);
  not (_05456_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_05457_, _00607_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_05458_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01853_);
  nor (_05459_, _05458_, _05457_);
  and (_05460_, _05459_, _05456_);
  nor (_05461_, _05459_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05462_, _05461_, _05460_);
  not (_05463_, _05462_);
  nor (_05464_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_05465_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01853_);
  nor (_05466_, _05465_, _05464_);
  not (_05468_, _05466_);
  nor (_05469_, _00528_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_05470_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01853_);
  nor (_05471_, _05470_, _05469_);
  and (_05473_, _05471_, _05468_);
  nand (_05474_, _05473_, _05463_);
  and (_05475_, _05474_, _05455_);
  nor (_05477_, _05471_, _05468_);
  not (_05478_, _05477_);
  not (_05479_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_05480_, _05459_, _05479_);
  and (_05481_, _05459_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05482_, _05481_, _05480_);
  nor (_05483_, _05482_, _05478_);
  and (_05484_, _05471_, _05466_);
  not (_05485_, _05484_);
  nor (_05486_, _05459_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_05487_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05488_, _05459_, _05487_);
  or (_05489_, _05488_, _05486_);
  nor (_05490_, _05489_, _05485_);
  nor (_05492_, _05490_, _05483_);
  not (_05493_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05495_, _05459_, _05493_);
  nor (_05496_, _05459_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_05497_, _05471_, _05466_);
  not (_05498_, _05497_);
  or (_05499_, _05498_, _05496_);
  or (_05500_, _05499_, _05495_);
  and (_05501_, _05500_, _05492_);
  and (_05502_, _05501_, _05475_);
  nor (_05503_, _05459_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_05504_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05505_, _05459_, _05504_);
  or (_05507_, _05505_, _05503_);
  nor (_05508_, _05507_, _05485_);
  nor (_05509_, _05508_, _05455_);
  and (_05510_, _05459_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not (_05511_, _05459_);
  and (_05513_, _05511_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_05514_, _05513_, _05510_);
  not (_05515_, _05514_);
  nand (_05517_, _05515_, _05473_);
  and (_05518_, _05459_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_05519_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05521_, _05459_, _05519_);
  nor (_05522_, _05521_, _05518_);
  nor (_05523_, _05522_, _05478_);
  nor (_05524_, _05459_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_05525_, _05524_);
  not (_05526_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05528_, _05459_, _05526_);
  nor (_05529_, _05528_, _05498_);
  and (_05530_, _05529_, _05525_);
  nor (_05532_, _05530_, _05523_);
  and (_05533_, _05532_, _05517_);
  and (_05534_, _05533_, _05509_);
  nor (_05536_, _05534_, _05502_);
  not (_05537_, _05536_);
  and (_05538_, _05537_, word_in[7]);
  not (_05539_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_05541_, _05455_, _05539_);
  or (_05542_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_05543_, _05542_, _05541_);
  and (_05544_, _05543_, _05497_);
  or (_05545_, _05544_, _05459_);
  not (_05546_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_05547_, _05455_, _05546_);
  or (_05548_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_05549_, _05548_, _05547_);
  and (_05550_, _05549_, _05484_);
  not (_05551_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_05552_, _05455_, _05551_);
  or (_05553_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_05554_, _05553_, _05552_);
  and (_05555_, _05554_, _05473_);
  not (_05556_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_05557_, _05455_, _05556_);
  or (_05558_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_05559_, _05558_, _05557_);
  and (_05560_, _05559_, _05477_);
  or (_05561_, _05560_, _05555_);
  or (_05562_, _05561_, _05550_);
  or (_05563_, _05562_, _05545_);
  not (_05564_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_05565_, _05455_, _05564_);
  or (_05566_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05567_, _05566_, _05565_);
  and (_05568_, _05567_, _05497_);
  or (_05569_, _05568_, _05511_);
  not (_05570_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_05571_, _05455_, _05570_);
  or (_05573_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_05574_, _05573_, _05571_);
  and (_05575_, _05574_, _05473_);
  not (_05576_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_05577_, _05455_, _05576_);
  or (_05578_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_05580_, _05578_, _05577_);
  and (_05582_, _05580_, _05484_);
  or (_05583_, _05582_, _05575_);
  not (_05584_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_05585_, _05455_, _05584_);
  or (_05586_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_05588_, _05586_, _05585_);
  and (_05589_, _05588_, _05477_);
  or (_05590_, _05589_, _05583_);
  or (_05591_, _05590_, _05569_);
  and (_05592_, _05591_, _05563_);
  and (_05593_, _05592_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _05593_, _05538_);
  not (_05594_, _05455_);
  and (_05595_, _05466_, _05594_);
  not (_05596_, _05595_);
  and (_05597_, _05466_, _05455_);
  and (_05598_, _05597_, _05471_);
  nor (_05599_, _05597_, _05471_);
  nor (_05600_, _05599_, _05598_);
  not (_05601_, _05600_);
  nor (_05602_, _05601_, _05489_);
  nor (_05603_, _05598_, _05511_);
  and (_05604_, _05598_, _05511_);
  nor (_05605_, _05604_, _05603_);
  and (_05606_, _05605_, _05601_);
  and (_05607_, _05606_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_05608_, _05605_, _05600_);
  and (_05609_, _05608_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05610_, _05609_, _05607_);
  nor (_05611_, _05610_, _05602_);
  nor (_05612_, _05611_, _05596_);
  nor (_05613_, _05466_, _05455_);
  not (_05614_, _05613_);
  nor (_05615_, _05601_, _05462_);
  and (_05616_, _05606_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05617_, _05608_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_05618_, _05617_, _05616_);
  nor (_05619_, _05618_, _05615_);
  nor (_05620_, _05619_, _05614_);
  nor (_05621_, _05620_, _05612_);
  and (_05622_, _05468_, _05455_);
  not (_05623_, _05622_);
  nor (_05624_, _05601_, _05507_);
  and (_05625_, _05606_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_05626_, _05608_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05627_, _05626_, _05625_);
  nor (_05628_, _05627_, _05624_);
  nor (_05630_, _05628_, _05623_);
  not (_05631_, _05597_);
  nor (_05632_, _05601_, _05514_);
  and (_05633_, _05606_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05634_, _05608_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05635_, _05634_, _05633_);
  nor (_05636_, _05635_, _05632_);
  nor (_05637_, _05636_, _05631_);
  nor (_05638_, _05637_, _05630_);
  and (_05639_, _05638_, _05621_);
  or (_05640_, _05613_, _05597_);
  not (_05641_, _05640_);
  not (_05642_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_05643_, _05455_, _05642_);
  or (_05644_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_05645_, _05644_, _05643_);
  and (_05646_, _05645_, _05641_);
  not (_05647_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_05648_, _05455_, _05647_);
  or (_05649_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_05650_, _05649_, _05648_);
  and (_05651_, _05650_, _05640_);
  or (_05653_, _05651_, _05646_);
  and (_05654_, _05653_, _05608_);
  not (_05655_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_05656_, _05455_, _05655_);
  or (_05657_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_05659_, _05657_, _05656_);
  and (_05660_, _05659_, _05641_);
  not (_05661_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_05662_, _05455_, _05661_);
  or (_05663_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_05665_, _05663_, _05662_);
  and (_05666_, _05665_, _05640_);
  or (_05668_, _05666_, _05660_);
  and (_05669_, _05668_, _05606_);
  and (_05670_, _05600_, _05511_);
  not (_05671_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_05673_, _05455_, _05671_);
  or (_05674_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_05675_, _05674_, _05673_);
  and (_05676_, _05675_, _05641_);
  not (_05677_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_05678_, _05455_, _05677_);
  or (_05679_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_05680_, _05679_, _05678_);
  and (_05681_, _05680_, _05640_);
  or (_05682_, _05681_, _05676_);
  and (_05683_, _05682_, _05670_);
  and (_05684_, _05600_, _05459_);
  not (_05685_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_05686_, _05455_, _05685_);
  or (_05687_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_05688_, _05687_, _05686_);
  and (_05689_, _05688_, _05641_);
  not (_05690_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_05691_, _05455_, _05690_);
  or (_05692_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_05693_, _05692_, _05691_);
  and (_05694_, _05693_, _05640_);
  or (_05695_, _05694_, _05689_);
  and (_05696_, _05695_, _05684_);
  or (_05697_, _05696_, _05683_);
  or (_05698_, _05697_, _05669_);
  nor (_05699_, _05698_, _05654_);
  nor (_05700_, _05699_, _05639_);
  and (_05701_, _05639_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _05701_, _05700_);
  nor (_05703_, _05497_, _05484_);
  and (_05704_, _05484_, _05511_);
  and (_05705_, _05485_, _05459_);
  or (_05706_, _05705_, _05704_);
  nor (_05707_, _05706_, _05703_);
  and (_05708_, _05707_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_05709_, _05703_);
  and (_05710_, _05706_, _05709_);
  and (_05712_, _05710_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05714_, _05709_, _05489_);
  or (_05715_, _05714_, _05712_);
  nor (_05717_, _05715_, _05708_);
  nor (_05718_, _05717_, _05623_);
  not (_05719_, _05718_);
  nor (_05720_, _05709_, _05514_);
  and (_05721_, _05707_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05723_, _05710_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05724_, _05723_, _05721_);
  or (_05726_, _05724_, _05720_);
  nand (_05727_, _05726_, _05595_);
  and (_05728_, _05727_, _05719_);
  and (_05730_, _05707_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_05732_, _05730_);
  nor (_05733_, _05709_, _05507_);
  and (_05735_, _05710_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05736_, _05735_, _05733_);
  and (_05738_, _05736_, _05732_);
  nor (_05739_, _05738_, _05614_);
  nor (_05740_, _05709_, _05462_);
  and (_05741_, _05710_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05743_, _05707_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05744_, _05743_, _05741_);
  nor (_05746_, _05744_, _05740_);
  nor (_05747_, _05746_, _05631_);
  nor (_05749_, _05747_, _05739_);
  and (_05750_, _05749_, _05728_);
  and (_05751_, _05750_, word_in[23]);
  and (_05752_, _05549_, _05473_);
  and (_05753_, _05543_, _05484_);
  or (_05754_, _05753_, _05752_);
  and (_05755_, _05554_, _05477_);
  and (_05756_, _05559_, _05497_);
  or (_05757_, _05756_, _05755_);
  or (_05758_, _05757_, _05754_);
  or (_05759_, _05758_, _05706_);
  not (_05760_, _05706_);
  and (_05761_, _05580_, _05473_);
  and (_05762_, _05588_, _05497_);
  or (_05763_, _05762_, _05761_);
  and (_05764_, _05574_, _05477_);
  and (_05765_, _05567_, _05511_);
  or (_05766_, _05765_, _05764_);
  or (_05767_, _05766_, _05763_);
  or (_05768_, _05767_, _05760_);
  nand (_05769_, _05768_, _05759_);
  nor (_05770_, _05769_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _05770_, _05751_);
  and (_05771_, _05598_, _05459_);
  and (_05772_, _05771_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05773_, _05614_, _05471_);
  not (_05774_, _05773_);
  nand (_05775_, _05614_, _05471_);
  and (_05776_, _05775_, _05774_);
  not (_05777_, _05776_);
  nor (_05778_, _05777_, _05507_);
  nor (_05779_, _05775_, _05459_);
  and (_05780_, _05775_, _05459_);
  nor (_05781_, _05780_, _05779_);
  nor (_05782_, _05781_, _05776_);
  and (_05783_, _05782_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05784_, _05783_, _05778_);
  nor (_05785_, _05784_, _05631_);
  nor (_05786_, _05777_, _05514_);
  and (_05787_, _05781_, _05777_);
  and (_05788_, _05787_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05789_, _05782_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05790_, _05789_, _05788_);
  or (_05791_, _05790_, _05786_);
  and (_05792_, _05791_, _05622_);
  or (_05793_, _05792_, _05785_);
  nor (_05794_, _05793_, _05772_);
  nor (_05795_, _05777_, _05462_);
  and (_05796_, _05787_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05797_, _05782_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_05798_, _05797_, _05796_);
  nor (_05799_, _05798_, _05795_);
  or (_05800_, _05799_, _05596_);
  and (_05801_, _05773_, _05480_);
  nor (_05802_, _05777_, _05489_);
  and (_05803_, _05782_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05804_, _05803_, _05802_);
  nor (_05805_, _05804_, _05614_);
  nor (_05806_, _05805_, _05801_);
  and (_05807_, _05806_, _05800_);
  and (_05808_, _05807_, _05794_);
  and (_05809_, _05665_, _05641_);
  and (_05810_, _05659_, _05640_);
  or (_05811_, _05810_, _05809_);
  and (_05813_, _05811_, _05787_);
  and (_05814_, _05650_, _05641_);
  and (_05815_, _05645_, _05640_);
  or (_05816_, _05815_, _05814_);
  and (_05817_, _05816_, _05782_);
  and (_05819_, _05776_, _05511_);
  and (_05820_, _05680_, _05641_);
  and (_05821_, _05675_, _05640_);
  or (_05822_, _05821_, _05820_);
  and (_05823_, _05822_, _05819_);
  and (_05824_, _05693_, _05641_);
  and (_05825_, _05688_, _05640_);
  or (_05826_, _05825_, _05824_);
  and (_05827_, _05780_, _05774_);
  and (_05829_, _05827_, _05826_);
  or (_05831_, _05829_, _05823_);
  or (_05832_, _05831_, _05817_);
  nor (_05833_, _05832_, _05813_);
  nor (_05834_, _05833_, _05808_);
  and (_05835_, _05808_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _05835_, _05834_);
  and (_05836_, _04532_, _23755_);
  and (_05838_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_00414_, _05838_, _05836_);
  and (_05839_, _05471_, _05459_);
  or (_05840_, _05839_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_26851_[15], _05840_, _22761_);
  and (_05842_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and (_05843_, _05439_, _23838_);
  or (_00460_, _05843_, _05842_);
  and (_05845_, _05613_, _05839_);
  and (_05846_, _05808_, _22761_);
  and (_05847_, _05846_, _05845_);
  not (_05848_, _05847_);
  and (_05849_, _05750_, _22761_);
  and (_05850_, _05849_, _05703_);
  and (_05851_, _05850_, _05706_);
  and (_05852_, _05851_, _05622_);
  and (_05853_, _05639_, _22761_);
  and (_05854_, _05853_, _05595_);
  and (_05855_, _05854_, _05684_);
  and (_05856_, _05502_, _22761_);
  and (_05857_, _05856_, _05466_);
  nor (_05858_, _05536_, rst);
  and (_05860_, _05858_, _05839_);
  and (_05861_, _05860_, _05857_);
  and (_05862_, _05858_, word_in[7]);
  and (_05864_, _05862_, _05861_);
  nor (_05865_, _05861_, _05576_);
  nor (_05866_, _05865_, _05864_);
  nor (_05867_, _05866_, _05855_);
  and (_05869_, _05855_, word_in[15]);
  nor (_05870_, _05869_, _05867_);
  nor (_05871_, _05870_, _05852_);
  and (_05872_, _05849_, word_in[23]);
  and (_05874_, _05872_, _05852_);
  or (_05875_, _05874_, _05871_);
  and (_05876_, _05875_, _05848_);
  and (_05877_, _05847_, word_in[31]);
  or (_26858_[7], _05877_, _05876_);
  or (_05879_, _05787_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_26868_, _05879_, _22761_);
  and (_05881_, _02277_, _23755_);
  and (_05882_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or (_00515_, _05882_, _05881_);
  and (_05884_, _05787_, _05595_);
  not (_05885_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05886_, _05498_, _05459_);
  not (_05887_, _05886_);
  nor (_05888_, _05887_, _05771_);
  nand (_05889_, _05888_, _05885_);
  or (_05890_, _05889_, _05884_);
  and (_26851_[1], _05890_, _22761_);
  and (_05891_, _05819_, _05595_);
  nor (_05892_, _05891_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_05893_, _05888_, _05892_);
  and (_26851_[2], _05893_, _22761_);
  not (_05894_, _05606_);
  and (_05895_, _05819_, _05597_);
  or (_05896_, _05471_, _05459_);
  or (_05898_, _05896_, _05595_);
  and (_05899_, _05898_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05900_, _05899_, _05895_);
  and (_05901_, _05900_, _05894_);
  and (_05903_, _05497_, _05480_);
  or (_05904_, _05903_, _05891_);
  or (_05906_, _05904_, _05901_);
  and (_05907_, _05906_, _05888_);
  or (_05908_, _05903_, _05900_);
  and (_05909_, _05908_, _05771_);
  or (_05911_, _05909_, _05887_);
  or (_05912_, _05911_, _05907_);
  and (_26851_[3], _05912_, _22761_);
  and (_05913_, _05471_, _05511_);
  and (_05914_, _05613_, _05913_);
  or (_05916_, _05914_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05917_, _05916_, _05896_);
  or (_05918_, _05917_, _05895_);
  and (_05919_, _05918_, _05894_);
  and (_05920_, _05916_, _05771_);
  and (_05921_, _05622_, _05819_);
  and (_05922_, _05773_, _05511_);
  and (_05923_, _05922_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_05924_, _05923_, _05921_);
  or (_05925_, _05924_, _05920_);
  or (_05926_, _05925_, _05891_);
  or (_05928_, _05926_, _05919_);
  and (_26851_[4], _05928_, _22761_);
  or (_05930_, _05779_, _05603_);
  or (_05931_, _05930_, _05771_);
  or (_05932_, _05484_, _05459_);
  or (_05933_, _05914_, _05895_);
  or (_05934_, _05933_, _05932_);
  and (_05935_, _05934_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05936_, _05891_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05938_, _05622_, _05913_);
  and (_05939_, _05887_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05940_, _05939_, _05938_);
  or (_05941_, _05940_, _05936_);
  or (_05943_, _05941_, _05935_);
  and (_05944_, _05943_, _05931_);
  and (_05945_, _05921_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05946_, _05922_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05947_, _05946_, _05891_);
  or (_05948_, _05947_, _05945_);
  or (_05950_, _05948_, _05914_);
  or (_05951_, _05950_, _05895_);
  or (_05952_, _05951_, _05944_);
  and (_26851_[5], _05952_, _22761_);
  and (_05953_, _02277_, _23635_);
  and (_05954_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or (_00741_, _05954_, _05953_);
  and (_05955_, _05595_, _05913_);
  or (_05956_, _05955_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_05957_, _05956_, _05931_);
  and (_05958_, _05957_, _05932_);
  and (_05959_, _05933_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05960_, _05959_, _05938_);
  or (_05961_, _05960_, _05958_);
  and (_05962_, _05961_, _05930_);
  and (_05963_, _05956_, _05771_);
  and (_05964_, _05891_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_05965_, _05887_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05966_, _05965_, _05895_);
  or (_05967_, _05966_, _05964_);
  or (_05968_, _05967_, _05914_);
  or (_05970_, _05968_, _05963_);
  or (_05971_, _05970_, _05962_);
  and (_26851_[6], _05971_, _22761_);
  and (_05972_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  and (_05973_, _03641_, _23589_);
  or (_00808_, _05973_, _05972_);
  and (_05974_, _25517_, _23676_);
  and (_05975_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_00823_, _05975_, _05974_);
  and (_05976_, _05459_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05977_, _05819_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05978_, _05922_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_05979_, _05978_, _05914_);
  or (_05980_, _05979_, _05977_);
  or (_05981_, _05980_, _05955_);
  or (_05983_, _05981_, _05976_);
  or (_05985_, _05983_, _05938_);
  or (_05986_, _05985_, _05604_);
  and (_26851_[7], _05986_, _22761_);
  and (_05988_, _25517_, _23718_);
  and (_05990_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_00854_, _05990_, _05988_);
  and (_05991_, _25517_, _23791_);
  and (_05993_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_00898_, _05993_, _05991_);
  or (_05994_, _05819_, _05782_);
  or (_05996_, _05994_, _05922_);
  nor (_05997_, _05996_, _05526_);
  and (_05999_, _05773_, _05459_);
  and (_06000_, _05914_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_06001_, _05896_, _05526_);
  or (_06002_, _06001_, _05604_);
  or (_06003_, _06002_, _05938_);
  or (_06004_, _06003_, _06000_);
  or (_06006_, _06004_, _05999_);
  or (_06007_, _06006_, _05955_);
  or (_06008_, _06007_, _05997_);
  and (_26851_[8], _06008_, _22761_);
  and (_06009_, _23643_, _23017_);
  and (_06010_, _06009_, _23791_);
  not (_06011_, _06009_);
  and (_06012_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_00913_, _06012_, _06010_);
  and (_06013_, _05938_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_06014_, _05819_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_06015_, _06014_, _06013_);
  and (_06016_, _05827_, _05622_);
  or (_06017_, _06016_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_06018_, _05774_, _05603_);
  and (_06019_, _06018_, _06017_);
  and (_06020_, _06019_, _05485_);
  or (_06021_, _06020_, _05773_);
  and (_06022_, _06021_, _05459_);
  and (_06023_, _05704_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_06025_, _06019_, _06023_);
  and (_06026_, _06025_, _05884_);
  and (_06027_, _05773_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_06029_, _06027_, _05598_);
  and (_06030_, _06029_, _05511_);
  and (_06031_, _06017_, _05771_);
  or (_06033_, _06031_, _05955_);
  or (_06035_, _06033_, _06030_);
  or (_06036_, _06035_, _06026_);
  or (_06037_, _06036_, _06022_);
  or (_06038_, _06037_, _06015_);
  and (_26851_[9], _06038_, _22761_);
  and (_06040_, _24615_, _23842_);
  not (_06041_, _06040_);
  and (_06042_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_06043_, _06040_, _23755_);
  or (_27119_, _06043_, _06042_);
  and (_06044_, _24118_, _23849_);
  and (_06045_, _06044_, _23791_);
  not (_06046_, _06044_);
  and (_06047_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_01039_, _06047_, _06045_);
  and (_06049_, _05498_, _05459_);
  and (_06051_, _06016_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_06052_, _05599_);
  and (_06053_, _06052_, _05518_);
  and (_06054_, _05922_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_06055_, _06054_, _06053_);
  or (_06056_, _06055_, _06051_);
  and (_06057_, _05780_, _05595_);
  or (_06058_, _05999_, _05604_);
  and (_06059_, _06058_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_06061_, _06059_, _06057_);
  or (_06062_, _06061_, _06056_);
  and (_06063_, _05641_, _05819_);
  or (_06064_, _05670_, _06063_);
  and (_06065_, _06064_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_06066_, _06065_, _06062_);
  and (_06067_, _06066_, _06049_);
  and (_06069_, _05703_, _05511_);
  and (_06070_, _06069_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_06071_, _05955_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_06073_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_06074_, _05886_, _06073_);
  or (_06075_, _06074_, _05604_);
  or (_06076_, _06075_, _06071_);
  or (_06077_, _06076_, _06016_);
  or (_06078_, _06077_, _06070_);
  or (_06079_, _06078_, _05999_);
  or (_06080_, _06079_, _06067_);
  and (_26851_[10], _06080_, _22761_);
  and (_06081_, _23962_, _23028_);
  and (_06082_, _06081_, _23755_);
  not (_06083_, _06081_);
  and (_06084_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or (_01070_, _06084_, _06082_);
  and (_06085_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_06086_, _24616_, _23755_);
  or (_01092_, _06086_, _06085_);
  and (_06088_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_06089_, _06040_, _23589_);
  or (_01095_, _06089_, _06088_);
  nand (_06090_, _25711_, _23585_);
  and (_06092_, _25691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_06093_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_06094_, _06093_, _02080_);
  nor (_06095_, _06094_, _25691_);
  or (_06097_, _06095_, _25699_);
  or (_06098_, _06097_, _06092_);
  nor (_06099_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_06100_, _06099_, _25667_);
  and (_06101_, _06100_, _06098_);
  nor (_06103_, _25711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_06104_, _06103_, _25712_);
  or (_06106_, _06104_, _06101_);
  and (_06107_, _06106_, _22761_);
  and (_01097_, _06107_, _06090_);
  and (_06108_, _06081_, _23589_);
  and (_06110_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or (_01116_, _06110_, _06108_);
  not (_06111_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_06112_, _06049_, _06111_);
  or (_06113_, _05999_, _06016_);
  and (_06114_, _05780_, _05597_);
  and (_06115_, _05839_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_06117_, _06115_, _06114_);
  or (_06118_, _06117_, _06113_);
  or (_06120_, _06118_, _06057_);
  or (_06121_, _06120_, _06112_);
  and (_26851_[11], _06121_, _22761_);
  and (_06123_, _02465_, _24671_);
  nand (_06124_, _06123_, _23522_);
  or (_06125_, _06123_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_06126_, _06125_, _02472_);
  and (_06127_, _06126_, _06124_);
  nor (_06129_, _02472_, _23585_);
  or (_06130_, _06129_, _06127_);
  and (_01176_, _06130_, _22761_);
  or (_06131_, _02869_, _02799_);
  and (_06132_, _06131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_06133_, _06132_, _02827_);
  and (_01184_, _06133_, _22761_);
  nor (_01186_, _04625_, rst);
  and (_06136_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_06137_, _02100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_01202_, _06137_, _06136_);
  and (_06138_, _05614_, _05839_);
  and (_06139_, _06138_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_06140_, _05996_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_06142_, _06140_, _05827_);
  or (_06143_, _06142_, _06139_);
  and (_26851_[12], _06143_, _22761_);
  or (_06144_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_06146_, _06144_, _22761_);
  and (_06147_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_06148_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_06149_, _06148_, rxd_i);
  or (_06150_, _06149_, _06147_);
  and (_06151_, _06150_, _02711_);
  and (_06152_, _02730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_06154_, _06152_, _06151_);
  and (_06155_, _02721_, rxd_i);
  or (_06156_, _06155_, _02728_);
  or (_06157_, _06156_, _06154_);
  and (_01217_, _06157_, _06146_);
  and (_06158_, _03046_, _23718_);
  and (_06159_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_01221_, _06159_, _06158_);
  and (_06161_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  and (_06162_, _03641_, _23718_);
  or (_01242_, _06162_, _06161_);
  not (_06164_, _25667_);
  nor (_06165_, _06164_, _23585_);
  and (_06166_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_06168_, _06166_, _25674_);
  and (_06169_, _06168_, _25701_);
  nand (_06171_, _25681_, _25674_);
  and (_06172_, _06171_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_06174_, _06171_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_06175_, _06174_, _25699_);
  or (_06176_, _06175_, _06172_);
  or (_06177_, _06176_, _06169_);
  nor (_06178_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_06179_, _06178_, _25667_);
  and (_06181_, _06179_, _06177_);
  or (_06183_, _06181_, _25711_);
  or (_06184_, _06183_, _06165_);
  or (_06185_, _25716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_06186_, _06185_, _22761_);
  and (_01248_, _06186_, _06184_);
  not (_06187_, _25695_);
  and (_06188_, _25712_, _25674_);
  and (_06189_, _06188_, _06187_);
  not (_06190_, _06189_);
  or (_06191_, _06190_, _25701_);
  or (_06192_, _06189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_06193_, _06192_, _22761_);
  and (_01256_, _06193_, _06191_);
  or (_06194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_06195_, _00308_, _24797_);
  or (_06196_, _06195_, _06194_);
  nand (_06197_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_06198_, _06197_, _06195_);
  or (_06200_, _06198_, _03826_);
  and (_06201_, _06200_, _06196_);
  and (_06202_, _25666_, _24714_);
  or (_06203_, _06202_, _06201_);
  nand (_06204_, _06202_, _23585_);
  and (_06205_, _06204_, _22761_);
  and (_01259_, _06205_, _06203_);
  not (_06207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor (_06208_, _25712_, _06207_);
  nor (_06209_, _25699_, _06187_);
  and (_06210_, _06209_, _25701_);
  and (_06211_, _06210_, _06188_);
  or (_06212_, _06211_, _06208_);
  and (_01261_, _06212_, _22761_);
  and (_06214_, _02815_, _02707_);
  and (_06215_, _02801_, _06214_);
  nand (_06216_, _06215_, _02829_);
  or (_06217_, _06215_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_06218_, _06217_, _22761_);
  and (_01265_, _06218_, _06216_);
  or (_06220_, _04675_, rxd_i);
  nand (_06222_, _06220_, _02715_);
  or (_06223_, _02716_, _02704_);
  and (_06224_, _06223_, _06222_);
  or (_06225_, _02720_, _02705_);
  or (_06227_, _06225_, _02714_);
  or (_06228_, _06227_, _06224_);
  and (_01269_, _06228_, _02100_);
  or (_06229_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_06230_, _06229_, _22761_);
  nand (_06231_, _02086_, _23585_);
  and (_01277_, _06231_, _06230_);
  not (_06233_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_06234_, _02586_, _06233_);
  or (_06235_, _06234_, _04641_);
  and (_06236_, _06235_, _02582_);
  nand (_06238_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_06239_, _06238_, _02581_);
  nor (_06240_, _06239_, _06236_);
  nor (_06241_, _06240_, _02580_);
  or (_06242_, _06241_, _02697_);
  nand (_06243_, _06242_, _22761_);
  nor (_01279_, _06243_, _02592_);
  and (_06244_, _03046_, _23791_);
  and (_06245_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_01283_, _06245_, _06244_);
  and (_06246_, _05706_, _05703_);
  or (_06247_, _06246_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_26851_[13], _06247_, _22761_);
  and (_06248_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  and (_06250_, _03641_, _23791_);
  or (_01310_, _06250_, _06248_);
  and (_06251_, _06081_, _23791_);
  and (_06253_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_01354_, _06253_, _06251_);
  or (_06254_, _05684_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_26851_[14], _06254_, _22761_);
  and (_06255_, _24572_, _23854_);
  and (_06256_, _06255_, _23589_);
  not (_06257_, _06255_);
  and (_06258_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or (_27161_, _06258_, _06256_);
  and (_06259_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_06260_, _24616_, _23718_);
  or (_01364_, _06260_, _06259_);
  and (_06261_, _06081_, _23676_);
  and (_06262_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or (_01367_, _06262_, _06261_);
  and (_06264_, _05322_, _23854_);
  and (_06265_, _06264_, _23982_);
  not (_06267_, _06264_);
  and (_06268_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_01371_, _06268_, _06265_);
  and (_06269_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_06270_, _24616_, _23791_);
  or (_01382_, _06270_, _06269_);
  and (_06271_, _03001_, _23676_);
  and (_06273_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or (_01407_, _06273_, _06271_);
  and (_06274_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_06275_, _03657_, _23791_);
  or (_01423_, _06275_, _06274_);
  and (_06276_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and (_06277_, _03657_, _23676_);
  or (_01431_, _06277_, _06276_);
  and (_06279_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and (_06280_, _05439_, _23982_);
  or (_01494_, _06280_, _06279_);
  and (_06281_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and (_06282_, _05439_, _23755_);
  or (_01500_, _06282_, _06281_);
  and (_06283_, _03281_, _23791_);
  and (_06284_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_27180_, _06284_, _06283_);
  and (_06285_, _03281_, _23589_);
  and (_06286_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_01518_, _06286_, _06285_);
  and (_06288_, _03281_, _23635_);
  and (_06289_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_01520_, _06289_, _06288_);
  and (_06290_, _02276_, _23594_);
  and (_06292_, _06290_, _23838_);
  not (_06293_, _06290_);
  and (_06294_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  or (_01523_, _06294_, _06292_);
  and (_06296_, _24558_, _24103_);
  not (_06298_, _06296_);
  and (_06299_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  and (_06300_, _06296_, _23791_);
  or (_01566_, _06300_, _06299_);
  and (_06301_, _02459_, _23755_);
  and (_06302_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or (_01568_, _06302_, _06301_);
  and (_06303_, _06290_, _23589_);
  and (_06304_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or (_27181_, _06304_, _06303_);
  and (_06305_, _03234_, _23589_);
  and (_06306_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or (_01618_, _06306_, _06305_);
  and (_06307_, _03264_, _23838_);
  and (_06308_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_01633_, _06308_, _06307_);
  and (_06309_, _02785_, _23718_);
  and (_06310_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  or (_01659_, _06310_, _06309_);
  and (_06311_, _05849_, _05884_);
  not (_06312_, _06311_);
  and (_06313_, _05853_, _05771_);
  not (_06315_, _06313_);
  and (_06316_, _05858_, _05466_);
  nor (_06317_, _06316_, _05856_);
  and (_06318_, _05858_, _05896_);
  not (_06320_, _06318_);
  and (_06322_, _06320_, _06317_);
  and (_06323_, _06322_, _05858_);
  and (_06325_, _06323_, word_in[0]);
  not (_06326_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_06327_, _06323_, _06326_);
  or (_06328_, _06327_, _06325_);
  and (_06329_, _06328_, _06315_);
  and (_06330_, _06313_, word_in[8]);
  or (_06331_, _06330_, _06329_);
  and (_06332_, _06331_, _06312_);
  and (_06334_, _05622_, _05839_);
  and (_06335_, _05846_, _06334_);
  and (_06336_, _05849_, word_in[16]);
  and (_06337_, _06336_, _05884_);
  or (_06338_, _06337_, _06335_);
  or (_06339_, _06338_, _06332_);
  not (_06340_, _06335_);
  or (_06341_, _06340_, word_in[24]);
  and (_26852_[0], _06341_, _06339_);
  and (_06342_, _03260_, _23589_);
  and (_06343_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_01677_, _06343_, _06342_);
  not (_06344_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_06345_, _06323_, _06344_);
  and (_06346_, _05858_, word_in[1]);
  and (_06347_, _06346_, _06322_);
  or (_06348_, _06347_, _06345_);
  or (_06350_, _06348_, _06313_);
  or (_06351_, _06315_, word_in[9]);
  and (_06352_, _06351_, _06312_);
  and (_06353_, _06352_, _06350_);
  and (_06355_, _06311_, word_in[17]);
  or (_06356_, _06355_, _06353_);
  and (_06357_, _06356_, _06340_);
  and (_06358_, _06335_, word_in[25]);
  or (_26852_[1], _06358_, _06357_);
  or (_06359_, _06315_, word_in[10]);
  and (_06360_, _06359_, _06312_);
  not (_06361_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_06362_, _06323_, _06361_);
  and (_06363_, _06323_, word_in[2]);
  or (_06364_, _06363_, _06362_);
  or (_06366_, _06364_, _06313_);
  and (_06367_, _06366_, _06360_);
  and (_06368_, _06311_, word_in[18]);
  or (_06369_, _06368_, _06335_);
  or (_06370_, _06369_, _06367_);
  or (_06371_, _06340_, word_in[26]);
  and (_26852_[2], _06371_, _06370_);
  and (_06373_, _02276_, _23854_);
  and (_06375_, _06373_, _23838_);
  not (_06376_, _06373_);
  and (_06377_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_01684_, _06377_, _06375_);
  or (_06379_, _06315_, word_in[11]);
  and (_06380_, _06379_, _06312_);
  and (_06381_, _06323_, word_in[3]);
  not (_06383_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_06384_, _06323_, _06383_);
  or (_06386_, _06384_, _06381_);
  or (_06387_, _06386_, _06313_);
  and (_06388_, _06387_, _06380_);
  and (_06390_, _06311_, word_in[19]);
  or (_06391_, _06390_, _06335_);
  or (_06393_, _06391_, _06388_);
  or (_06395_, _06340_, word_in[27]);
  and (_26852_[3], _06395_, _06393_);
  and (_06396_, _06311_, word_in[20]);
  or (_06397_, _06315_, word_in[12]);
  and (_06398_, _06397_, _06312_);
  not (_06399_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_06401_, _06323_, _06399_);
  and (_06402_, _06323_, word_in[4]);
  or (_06403_, _06402_, _06401_);
  or (_06404_, _06403_, _06313_);
  and (_06406_, _06404_, _06398_);
  or (_06407_, _06406_, _06396_);
  and (_06408_, _06407_, _06340_);
  and (_06409_, _06335_, word_in[28]);
  or (_26852_[4], _06409_, _06408_);
  and (_06410_, _06373_, _23791_);
  and (_06411_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_01690_, _06411_, _06410_);
  and (_06412_, _05846_, word_in[29]);
  and (_06413_, _06412_, _06335_);
  or (_06414_, _06315_, word_in[13]);
  and (_06415_, _06414_, _06312_);
  and (_06416_, _06323_, word_in[5]);
  not (_06417_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_06418_, _06323_, _06417_);
  or (_06419_, _06418_, _06416_);
  or (_06420_, _06419_, _06313_);
  and (_06421_, _06420_, _06415_);
  and (_06422_, _06311_, word_in[21]);
  or (_06423_, _06422_, _06421_);
  and (_06424_, _06423_, _06340_);
  or (_26852_[5], _06424_, _06413_);
  or (_06425_, _06315_, word_in[14]);
  and (_06426_, _06425_, _06312_);
  not (_06427_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_06428_, _06323_, _06427_);
  and (_06429_, _06323_, word_in[6]);
  or (_06430_, _06429_, _06428_);
  or (_06431_, _06430_, _06313_);
  and (_06432_, _06431_, _06426_);
  and (_06434_, _06311_, word_in[22]);
  or (_06436_, _06434_, _06335_);
  or (_06438_, _06436_, _06432_);
  or (_06439_, _06340_, word_in[30]);
  and (_26852_[6], _06439_, _06438_);
  or (_06441_, _06340_, word_in[31]);
  nor (_06443_, _06323_, _05661_);
  and (_06444_, _06323_, _05862_);
  or (_06445_, _06444_, _06443_);
  or (_06446_, _06445_, _06313_);
  or (_06448_, _06315_, word_in[15]);
  and (_06449_, _06448_, _06312_);
  and (_06451_, _06449_, _06446_);
  and (_06452_, _06311_, word_in[23]);
  or (_06454_, _06452_, _06335_);
  or (_06455_, _06454_, _06451_);
  and (_26852_[7], _06455_, _06441_);
  and (_06457_, _03335_, _23676_);
  and (_06458_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_27191_, _06458_, _06457_);
  and (_06460_, _06373_, _23755_);
  and (_06462_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_01711_, _06462_, _06460_);
  and (_06464_, _03335_, _23755_);
  and (_06466_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_01718_, _06466_, _06464_);
  and (_06467_, _03335_, _23838_);
  and (_06469_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_01731_, _06469_, _06467_);
  and (_06470_, _03326_, _23676_);
  and (_06471_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_01758_, _06471_, _06470_);
  and (_06472_, _05846_, _05884_);
  not (_06474_, _06472_);
  and (_06475_, _05853_, _05613_);
  and (_06476_, _06475_, _05606_);
  not (_06477_, _06476_);
  not (_06478_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_06479_, _05856_, _05468_);
  and (_06480_, _06479_, _06320_);
  nor (_06481_, _06480_, _06478_);
  and (_06482_, _05858_, word_in[0]);
  and (_06484_, _06480_, _06482_);
  or (_06485_, _06484_, _06481_);
  and (_06486_, _06485_, _06477_);
  and (_06487_, _05849_, _05597_);
  and (_06488_, _06487_, _05707_);
  and (_06489_, _06476_, word_in[8]);
  or (_06490_, _06489_, _06488_);
  or (_06491_, _06490_, _06486_);
  not (_06492_, _06488_);
  or (_06493_, _06492_, _06336_);
  and (_06494_, _06493_, _06491_);
  and (_06495_, _06494_, _06474_);
  and (_06496_, _06472_, word_in[24]);
  or (_26859_[0], _06496_, _06495_);
  and (_06497_, _03326_, _23589_);
  and (_06499_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_27196_, _06499_, _06497_);
  and (_06500_, _05849_, word_in[17]);
  or (_06501_, _06492_, _06500_);
  not (_06502_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_06504_, _06480_, _06502_);
  and (_06505_, _06480_, _06346_);
  or (_06506_, _06505_, _06504_);
  and (_06507_, _06506_, _06477_);
  and (_06508_, _06476_, word_in[9]);
  or (_06509_, _06508_, _06488_);
  or (_06510_, _06509_, _06507_);
  and (_06511_, _06510_, _06501_);
  and (_06512_, _06511_, _06474_);
  and (_06513_, _06472_, word_in[25]);
  or (_26859_[1], _06513_, _06512_);
  and (_06514_, _05849_, word_in[18]);
  or (_06515_, _06492_, _06514_);
  not (_06516_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_06517_, _06480_, _06516_);
  and (_06519_, _05858_, word_in[2]);
  and (_06521_, _06480_, _06519_);
  or (_06522_, _06521_, _06517_);
  and (_06524_, _06522_, _06477_);
  and (_06525_, _06476_, word_in[10]);
  or (_06527_, _06525_, _06488_);
  or (_06528_, _06527_, _06524_);
  and (_06529_, _06528_, _06515_);
  and (_06530_, _06529_, _06474_);
  and (_06531_, _06472_, word_in[26]);
  or (_26859_[2], _06531_, _06530_);
  and (_06532_, _03326_, _23635_);
  and (_06533_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_01779_, _06533_, _06532_);
  and (_06534_, _05849_, word_in[19]);
  or (_06535_, _06492_, _06534_);
  not (_06536_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_06537_, _06480_, _06536_);
  and (_06538_, _05858_, word_in[3]);
  and (_06539_, _06480_, _06538_);
  or (_06540_, _06539_, _06537_);
  and (_06541_, _06540_, _06477_);
  and (_06542_, _06476_, word_in[11]);
  or (_06543_, _06542_, _06488_);
  or (_06544_, _06543_, _06541_);
  and (_06546_, _06544_, _06535_);
  and (_06547_, _06546_, _06474_);
  and (_06548_, _06472_, word_in[27]);
  or (_26859_[3], _06548_, _06547_);
  and (_06549_, _05849_, word_in[20]);
  or (_06550_, _06492_, _06549_);
  not (_06551_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_06552_, _06480_, _06551_);
  and (_06554_, _05858_, word_in[4]);
  and (_06555_, _06480_, _06554_);
  or (_06557_, _06555_, _06552_);
  and (_06558_, _06557_, _06477_);
  and (_06560_, _06476_, word_in[12]);
  or (_06561_, _06560_, _06488_);
  or (_06562_, _06561_, _06558_);
  and (_06563_, _06562_, _06550_);
  and (_06564_, _06563_, _06474_);
  and (_06565_, _06472_, word_in[28]);
  or (_26859_[4], _06565_, _06564_);
  and (_06566_, _05849_, word_in[21]);
  or (_06567_, _06492_, _06566_);
  not (_06568_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_06569_, _06480_, _06568_);
  and (_06570_, _05858_, word_in[5]);
  and (_06571_, _06480_, _06570_);
  or (_06572_, _06571_, _06569_);
  and (_06573_, _06572_, _06477_);
  and (_06574_, _06476_, word_in[13]);
  or (_06575_, _06574_, _06488_);
  or (_06576_, _06575_, _06573_);
  and (_06577_, _06576_, _06567_);
  and (_06578_, _06577_, _06474_);
  and (_06579_, _06472_, word_in[29]);
  or (_26859_[5], _06579_, _06578_);
  and (_06580_, _05849_, word_in[22]);
  or (_06581_, _06492_, _06580_);
  not (_06582_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_06583_, _06480_, _06582_);
  and (_06585_, _05858_, word_in[6]);
  and (_06586_, _06480_, _06585_);
  or (_06587_, _06586_, _06583_);
  and (_06588_, _06587_, _06477_);
  and (_06589_, _06476_, word_in[14]);
  or (_06590_, _06589_, _06488_);
  or (_06591_, _06590_, _06588_);
  and (_06593_, _06591_, _06581_);
  and (_06594_, _06593_, _06474_);
  and (_06595_, _06472_, word_in[30]);
  or (_26859_[6], _06595_, _06594_);
  or (_06596_, _06492_, _05872_);
  nor (_06597_, _06480_, _05539_);
  and (_06598_, _06480_, _05862_);
  or (_06599_, _06598_, _06597_);
  and (_06600_, _06599_, _06477_);
  and (_06601_, _06476_, word_in[15]);
  or (_06602_, _06601_, _06488_);
  or (_06603_, _06602_, _06600_);
  and (_06604_, _06603_, _06596_);
  and (_06605_, _06604_, _06474_);
  and (_06606_, _06472_, word_in[31]);
  or (_26859_[7], _06606_, _06605_);
  and (_06607_, _05846_, _05597_);
  and (_06608_, _06607_, _05787_);
  and (_06609_, _05849_, _05613_);
  and (_06610_, _06609_, _05707_);
  not (_06611_, _06610_);
  or (_06612_, _06611_, _06336_);
  and (_06613_, _05853_, _05622_);
  and (_06614_, _06613_, _05606_);
  not (_06615_, _06614_);
  not (_06616_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not (_06617_, _05856_);
  and (_06618_, _06316_, _06617_);
  and (_06620_, _06618_, _06320_);
  nor (_06621_, _06620_, _06616_);
  and (_06622_, _06620_, _06482_);
  or (_06623_, _06622_, _06621_);
  and (_06624_, _06623_, _06615_);
  and (_06625_, _06614_, word_in[8]);
  or (_06626_, _06625_, _06610_);
  or (_06627_, _06626_, _06624_);
  and (_06628_, _06627_, _06612_);
  or (_06629_, _06628_, _06608_);
  not (_06630_, _06608_);
  or (_06631_, _06630_, word_in[24]);
  and (_26860_[0], _06631_, _06629_);
  or (_06632_, _06611_, _06500_);
  not (_06633_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_06634_, _06620_, _06633_);
  and (_06635_, _06620_, _06346_);
  or (_06636_, _06635_, _06634_);
  and (_06637_, _06636_, _06615_);
  and (_06638_, _06614_, word_in[9]);
  or (_06639_, _06638_, _06610_);
  or (_06640_, _06639_, _06637_);
  and (_06642_, _06640_, _06632_);
  or (_06644_, _06642_, _06608_);
  or (_06645_, _06630_, word_in[25]);
  and (_26860_[1], _06645_, _06644_);
  or (_06646_, _06611_, _06514_);
  not (_06647_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_06648_, _06620_, _06647_);
  and (_06649_, _06620_, _06519_);
  or (_06651_, _06649_, _06648_);
  and (_06652_, _06651_, _06615_);
  and (_06653_, _06614_, word_in[10]);
  or (_06654_, _06653_, _06610_);
  or (_06655_, _06654_, _06652_);
  and (_06656_, _06655_, _06646_);
  or (_06658_, _06656_, _06608_);
  or (_06659_, _06630_, word_in[26]);
  and (_26860_[2], _06659_, _06658_);
  or (_06660_, _06611_, _06534_);
  not (_06661_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_06662_, _06620_, _06661_);
  and (_06663_, _06620_, _06538_);
  or (_06664_, _06663_, _06662_);
  and (_06665_, _06664_, _06615_);
  and (_06666_, _06614_, word_in[11]);
  or (_06667_, _06666_, _06610_);
  or (_06668_, _06667_, _06665_);
  and (_06669_, _06668_, _06660_);
  or (_06670_, _06669_, _06608_);
  or (_06671_, _06630_, word_in[27]);
  and (_26860_[3], _06671_, _06670_);
  not (_06672_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_06673_, _06620_, _06672_);
  and (_06674_, _06620_, _06554_);
  or (_06675_, _06674_, _06673_);
  and (_06676_, _06675_, _06615_);
  and (_06677_, _06614_, word_in[12]);
  or (_06678_, _06677_, _06610_);
  or (_06679_, _06678_, _06676_);
  or (_06680_, _06611_, _06549_);
  and (_06681_, _06680_, _06679_);
  or (_06682_, _06681_, _06608_);
  or (_06683_, _06630_, word_in[28]);
  and (_26860_[4], _06683_, _06682_);
  or (_06684_, _06611_, _06566_);
  not (_06685_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_06686_, _06620_, _06685_);
  and (_06687_, _06620_, _06570_);
  or (_06688_, _06687_, _06686_);
  and (_06690_, _06688_, _06615_);
  and (_06691_, _06614_, word_in[13]);
  or (_06692_, _06691_, _06610_);
  or (_06693_, _06692_, _06690_);
  and (_06694_, _06693_, _06684_);
  or (_06695_, _06694_, _06608_);
  or (_06696_, _06630_, word_in[29]);
  and (_26860_[5], _06696_, _06695_);
  and (_06697_, _23755_, _23029_);
  and (_06699_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or (_01856_, _06699_, _06697_);
  or (_06701_, _06611_, _06580_);
  not (_06702_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_06703_, _06620_, _06702_);
  and (_06704_, _06620_, _06585_);
  or (_06705_, _06704_, _06703_);
  and (_06706_, _06705_, _06615_);
  and (_06707_, _06614_, word_in[14]);
  or (_06708_, _06707_, _06610_);
  or (_06709_, _06708_, _06706_);
  and (_06710_, _06709_, _06701_);
  or (_06711_, _06710_, _06608_);
  or (_06712_, _06630_, word_in[30]);
  and (_26860_[6], _06712_, _06711_);
  or (_06714_, _06611_, _05872_);
  nor (_06715_, _06620_, _05655_);
  and (_06716_, _06620_, _05862_);
  or (_06718_, _06716_, _06715_);
  and (_06719_, _06718_, _06615_);
  and (_06720_, _06614_, word_in[15]);
  or (_06721_, _06720_, _06610_);
  or (_06723_, _06721_, _06719_);
  and (_06724_, _06723_, _06714_);
  or (_06725_, _06724_, _06608_);
  or (_06726_, _06630_, word_in[31]);
  and (_26860_[7], _06726_, _06725_);
  and (_06727_, _05846_, _05922_);
  not (_06728_, _06727_);
  and (_06729_, _05854_, _05606_);
  not (_06730_, _06729_);
  not (_06731_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_06732_, _06320_, _05857_);
  nor (_06733_, _06732_, _06731_);
  and (_06734_, _06732_, _06482_);
  or (_06735_, _06734_, _06733_);
  and (_06736_, _06735_, _06730_);
  and (_06737_, _05849_, _05622_);
  and (_06738_, _06737_, _05707_);
  and (_06739_, _06729_, word_in[8]);
  or (_06740_, _06739_, _06738_);
  or (_06742_, _06740_, _06736_);
  not (_06743_, _06738_);
  or (_06745_, _06743_, _06336_);
  and (_06746_, _06745_, _06742_);
  and (_06747_, _06746_, _06728_);
  and (_06748_, _06727_, word_in[24]);
  or (_26861_[0], _06748_, _06747_);
  or (_06749_, _06743_, _06500_);
  not (_06751_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_06752_, _06732_, _06751_);
  and (_06753_, _06732_, _06346_);
  or (_06754_, _06753_, _06752_);
  and (_06755_, _06754_, _06730_);
  and (_06757_, _06729_, word_in[9]);
  or (_06758_, _06757_, _06738_);
  or (_06759_, _06758_, _06755_);
  and (_06760_, _06759_, _06749_);
  and (_06763_, _06760_, _06728_);
  and (_06764_, _06727_, word_in[25]);
  or (_26861_[1], _06764_, _06763_);
  or (_06765_, _06743_, _06514_);
  not (_06766_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_06767_, _06732_, _06766_);
  and (_06768_, _06732_, _06519_);
  or (_06769_, _06768_, _06767_);
  and (_06770_, _06769_, _06730_);
  and (_06772_, _06729_, word_in[10]);
  or (_06773_, _06772_, _06738_);
  or (_06774_, _06773_, _06770_);
  and (_06775_, _06774_, _06765_);
  and (_06776_, _06775_, _06728_);
  and (_06777_, _06727_, word_in[26]);
  or (_26861_[2], _06777_, _06776_);
  or (_06778_, _06743_, _06534_);
  not (_06779_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_06780_, _06732_, _06779_);
  and (_06781_, _06732_, _06538_);
  or (_06782_, _06781_, _06780_);
  and (_06783_, _06782_, _06730_);
  and (_06784_, _06729_, word_in[11]);
  or (_06786_, _06784_, _06738_);
  or (_06787_, _06786_, _06783_);
  and (_06788_, _06787_, _06778_);
  and (_06789_, _06788_, _06728_);
  and (_06790_, _06727_, word_in[27]);
  or (_26861_[3], _06790_, _06789_);
  or (_06791_, _06743_, _06549_);
  not (_06792_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_06793_, _06732_, _06792_);
  and (_06794_, _06732_, _06554_);
  or (_06795_, _06794_, _06793_);
  and (_06796_, _06795_, _06730_);
  and (_06797_, _06729_, word_in[12]);
  or (_06798_, _06797_, _06738_);
  or (_06799_, _06798_, _06796_);
  and (_06800_, _06799_, _06791_);
  and (_06801_, _06800_, _06728_);
  and (_06802_, _06727_, word_in[28]);
  or (_26861_[4], _06802_, _06801_);
  or (_06803_, _06743_, _06566_);
  not (_06804_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_06805_, _06732_, _06804_);
  and (_06806_, _06732_, _06570_);
  or (_06807_, _06806_, _06805_);
  and (_06809_, _06807_, _06730_);
  and (_06810_, _06729_, word_in[13]);
  or (_06811_, _06810_, _06738_);
  or (_06812_, _06811_, _06809_);
  and (_06813_, _06812_, _06803_);
  and (_06814_, _06813_, _06728_);
  and (_06815_, _06727_, word_in[29]);
  or (_26861_[5], _06815_, _06814_);
  or (_06816_, _06743_, _06580_);
  not (_06817_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_06818_, _06732_, _06817_);
  and (_06820_, _06732_, _06585_);
  or (_06821_, _06820_, _06818_);
  and (_06822_, _06821_, _06730_);
  and (_06823_, _06729_, word_in[14]);
  or (_06824_, _06823_, _06738_);
  or (_06826_, _06824_, _06822_);
  and (_06827_, _06826_, _06816_);
  and (_06828_, _06827_, _06728_);
  and (_06829_, _06727_, word_in[30]);
  or (_26861_[6], _06829_, _06828_);
  or (_06831_, _06743_, _05872_);
  nor (_06832_, _06732_, _05556_);
  and (_06833_, _06732_, _05862_);
  or (_06834_, _06833_, _06832_);
  and (_06835_, _06834_, _06730_);
  and (_06836_, _06729_, word_in[15]);
  or (_06837_, _06836_, _06738_);
  or (_06838_, _06837_, _06835_);
  and (_06839_, _06838_, _06831_);
  and (_06840_, _06839_, _06728_);
  and (_06841_, _06727_, word_in[31]);
  or (_26861_[7], _06841_, _06840_);
  and (_06842_, _05850_, _05760_);
  and (_06843_, _06842_, _05595_);
  and (_06844_, _05853_, _05895_);
  not (_06845_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_06846_, _05858_, _05913_);
  and (_06847_, _06846_, _06317_);
  nor (_06848_, _06847_, _06845_);
  and (_06849_, _06847_, _06482_);
  or (_06850_, _06849_, _06848_);
  or (_06851_, _06850_, _06844_);
  not (_06853_, _06844_);
  or (_06854_, _06853_, word_in[8]);
  and (_06855_, _06854_, _06851_);
  or (_06856_, _06855_, _06843_);
  and (_06857_, _05846_, _05921_);
  not (_06858_, _06857_);
  not (_06859_, _06843_);
  or (_06860_, _06859_, _06336_);
  and (_06861_, _06860_, _06858_);
  and (_06862_, _06861_, _06856_);
  and (_06863_, _06857_, word_in[24]);
  or (_26862_[0], _06863_, _06862_);
  and (_06864_, _06857_, word_in[25]);
  not (_06865_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_06866_, _06847_, _06865_);
  and (_06867_, _06847_, _06346_);
  or (_06868_, _06867_, _06866_);
  or (_06869_, _06868_, _06844_);
  or (_06870_, _06853_, word_in[9]);
  and (_06871_, _06870_, _06869_);
  or (_06872_, _06871_, _06843_);
  or (_06873_, _06859_, _06500_);
  and (_06874_, _06873_, _06858_);
  and (_06875_, _06874_, _06872_);
  or (_26862_[1], _06875_, _06864_);
  not (_06876_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_06877_, _06847_, _06876_);
  and (_06878_, _06847_, _06519_);
  or (_06879_, _06878_, _06877_);
  or (_06880_, _06879_, _06844_);
  or (_06881_, _06853_, word_in[10]);
  and (_06882_, _06881_, _06880_);
  or (_06883_, _06882_, _06843_);
  or (_06884_, _06859_, _06514_);
  and (_06885_, _06884_, _06858_);
  and (_06886_, _06885_, _06883_);
  and (_06887_, _06857_, word_in[26]);
  or (_26862_[2], _06887_, _06886_);
  not (_06889_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_06891_, _06847_, _06889_);
  and (_06893_, _06847_, _06538_);
  or (_06895_, _06893_, _06891_);
  or (_06896_, _06895_, _06844_);
  or (_06898_, _06853_, word_in[11]);
  and (_06899_, _06898_, _06896_);
  or (_06901_, _06899_, _06843_);
  or (_06902_, _06859_, _06534_);
  and (_06903_, _06902_, _06858_);
  and (_06905_, _06903_, _06901_);
  and (_06906_, _06857_, word_in[27]);
  or (_26862_[3], _06906_, _06905_);
  not (_06910_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_06912_, _06847_, _06910_);
  and (_06913_, _06847_, _06554_);
  or (_06915_, _06913_, _06912_);
  or (_06917_, _06915_, _06844_);
  or (_06919_, _06853_, word_in[12]);
  and (_06920_, _06919_, _06917_);
  or (_06921_, _06920_, _06843_);
  or (_06922_, _06859_, _06549_);
  and (_06924_, _06922_, _06858_);
  and (_06926_, _06924_, _06921_);
  and (_06927_, _06857_, word_in[28]);
  or (_26862_[4], _06927_, _06926_);
  not (_06929_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_06930_, _06847_, _06929_);
  and (_06931_, _06847_, _06570_);
  or (_06932_, _06931_, _06930_);
  or (_06933_, _06932_, _06844_);
  or (_06934_, _06853_, word_in[13]);
  and (_06936_, _06934_, _06933_);
  or (_06937_, _06936_, _06843_);
  or (_06938_, _06859_, _06566_);
  and (_06939_, _06938_, _06858_);
  and (_06940_, _06939_, _06937_);
  and (_06941_, _06857_, word_in[29]);
  or (_26862_[5], _06941_, _06940_);
  or (_06942_, _06859_, _06580_);
  not (_06943_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_06944_, _06847_, _06943_);
  and (_06945_, _06847_, _06585_);
  or (_06946_, _06945_, _06944_);
  and (_06947_, _06946_, _06853_);
  and (_06948_, _05853_, word_in[14]);
  and (_06949_, _06844_, _06948_);
  or (_06950_, _06949_, _06843_);
  or (_06951_, _06950_, _06947_);
  and (_06952_, _06951_, _06942_);
  and (_06953_, _06952_, _06858_);
  and (_06954_, _06857_, word_in[30]);
  or (_26862_[6], _06954_, _06953_);
  nor (_06957_, _06847_, _05677_);
  and (_06958_, _06847_, _05862_);
  or (_06959_, _06958_, _06957_);
  or (_06960_, _06959_, _06844_);
  or (_06961_, _06853_, word_in[15]);
  and (_06963_, _06961_, _06960_);
  or (_06964_, _06963_, _06843_);
  or (_06965_, _06859_, _05872_);
  and (_06967_, _06965_, _06858_);
  and (_06968_, _06967_, _06964_);
  and (_06969_, _06857_, word_in[31]);
  or (_26862_[7], _06969_, _06968_);
  and (_06971_, _25742_, _23589_);
  and (_06972_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_01998_, _06972_, _06971_);
  and (_06974_, _05846_, _05891_);
  not (_06976_, _06974_);
  and (_06977_, _06842_, _05597_);
  and (_06978_, _06475_, _05670_);
  not (_06979_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_06980_, _06846_, _06479_);
  nor (_06981_, _06980_, _06979_);
  and (_06983_, _06980_, _06482_);
  or (_06984_, _06983_, _06981_);
  or (_06985_, _06984_, _06978_);
  not (_06987_, _06978_);
  or (_06989_, _06987_, word_in[8]);
  and (_06990_, _06989_, _06985_);
  or (_06991_, _06990_, _06977_);
  not (_06992_, _06977_);
  or (_06993_, _06992_, _06336_);
  and (_06995_, _06993_, _06991_);
  and (_06996_, _06995_, _06976_);
  and (_06997_, _06974_, word_in[24]);
  or (_26863_[0], _06997_, _06996_);
  and (_06998_, _06977_, _06500_);
  not (_07000_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_07001_, _06980_, _07000_);
  and (_07002_, _06980_, _06346_);
  nor (_07005_, _07002_, _07001_);
  nor (_07006_, _07005_, _06978_);
  and (_07007_, _06978_, word_in[9]);
  nor (_07008_, _07007_, _07006_);
  nor (_07010_, _07008_, _06977_);
  or (_07011_, _07010_, _06998_);
  and (_07012_, _07011_, _06976_);
  and (_07014_, _06974_, word_in[25]);
  or (_26863_[1], _07014_, _07012_);
  and (_07015_, _06977_, _06514_);
  not (_07016_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_07018_, _06980_, _07016_);
  and (_07019_, _06980_, _06519_);
  nor (_07021_, _07019_, _07018_);
  nor (_07022_, _07021_, _06978_);
  and (_07024_, _06978_, word_in[10]);
  nor (_07025_, _07024_, _07022_);
  nor (_07026_, _07025_, _06977_);
  or (_07028_, _07026_, _07015_);
  and (_07029_, _07028_, _06976_);
  and (_07030_, _06974_, word_in[26]);
  or (_26863_[2], _07030_, _07029_);
  and (_07031_, _06977_, _06534_);
  and (_07032_, _06980_, _06538_);
  not (_07033_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_07034_, _06980_, _07033_);
  nor (_07035_, _07034_, _07032_);
  nor (_07036_, _07035_, _06978_);
  and (_07037_, _06978_, word_in[11]);
  nor (_07038_, _07037_, _07036_);
  nor (_07040_, _07038_, _06977_);
  or (_07041_, _07040_, _07031_);
  and (_07043_, _07041_, _06976_);
  and (_07044_, _06974_, word_in[27]);
  or (_26863_[3], _07044_, _07043_);
  and (_07045_, _06977_, _06549_);
  not (_07047_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_07048_, _06980_, _07047_);
  and (_07049_, _06980_, _06554_);
  nor (_07050_, _07049_, _07048_);
  nor (_07051_, _07050_, _06978_);
  and (_07052_, _06978_, word_in[12]);
  nor (_07053_, _07052_, _07051_);
  nor (_07054_, _07053_, _06977_);
  or (_07055_, _07054_, _07045_);
  and (_07056_, _07055_, _06976_);
  and (_07057_, _06974_, word_in[28]);
  or (_26863_[4], _07057_, _07056_);
  and (_07058_, _06977_, _06566_);
  and (_07059_, _06980_, _06570_);
  not (_07061_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_07062_, _06980_, _07061_);
  nor (_07063_, _07062_, _07059_);
  nor (_07064_, _07063_, _06978_);
  and (_07065_, _06978_, word_in[13]);
  nor (_07066_, _07065_, _07064_);
  nor (_07068_, _07066_, _06977_);
  or (_07069_, _07068_, _07058_);
  and (_07070_, _07069_, _06976_);
  and (_07071_, _06974_, word_in[29]);
  or (_26863_[5], _07071_, _07070_);
  and (_07072_, _06977_, _06580_);
  and (_07073_, _06980_, _06585_);
  not (_07074_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_07075_, _06980_, _07074_);
  nor (_07076_, _07075_, _07073_);
  nor (_07077_, _07076_, _06978_);
  and (_07079_, _06978_, word_in[14]);
  nor (_07081_, _07079_, _07077_);
  nor (_07083_, _07081_, _06977_);
  or (_07084_, _07083_, _07072_);
  and (_07085_, _07084_, _06976_);
  and (_07086_, _06974_, word_in[30]);
  or (_26863_[6], _07086_, _07085_);
  and (_07087_, _06977_, _05872_);
  nor (_07088_, _06980_, _05551_);
  and (_07090_, _06980_, _05862_);
  nor (_07091_, _07090_, _07088_);
  nor (_07092_, _07091_, _06978_);
  and (_07093_, _06978_, word_in[15]);
  nor (_07094_, _07093_, _07092_);
  nor (_07095_, _07094_, _06977_);
  or (_07096_, _07095_, _07087_);
  and (_07097_, _07096_, _06976_);
  and (_07099_, _06974_, word_in[31]);
  or (_26863_[7], _07099_, _07097_);
  and (_07101_, _24117_, _23599_);
  and (_07102_, _07101_, _23589_);
  not (_07103_, _07101_);
  and (_07104_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or (_02068_, _07104_, _07102_);
  and (_07107_, _07101_, _23755_);
  and (_07108_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or (_02085_, _07108_, _07107_);
  and (_07109_, _05846_, _05895_);
  not (_07110_, _07109_);
  and (_07111_, _06613_, _05670_);
  not (_07112_, _07111_);
  not (_07113_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_07115_, _06618_, _05913_);
  nor (_07116_, _07115_, _07113_);
  and (_07118_, _07115_, _06482_);
  or (_07119_, _07118_, _07116_);
  and (_07120_, _07119_, _07112_);
  and (_07122_, _06842_, _05613_);
  and (_07123_, _07111_, word_in[8]);
  or (_07124_, _07123_, _07122_);
  or (_07126_, _07124_, _07120_);
  not (_07127_, _07122_);
  or (_07128_, _07127_, _06336_);
  and (_07129_, _07128_, _07126_);
  and (_07130_, _07129_, _07110_);
  and (_07132_, _07109_, word_in[24]);
  or (_26864_[0], _07132_, _07130_);
  not (_07133_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_07134_, _07115_, _07133_);
  and (_07135_, _07115_, _06346_);
  or (_07136_, _07135_, _07134_);
  or (_07137_, _07136_, _07111_);
  or (_07138_, _07112_, word_in[9]);
  and (_07139_, _07138_, _07137_);
  or (_07140_, _07139_, _07122_);
  or (_07142_, _07127_, _06500_);
  and (_07143_, _07142_, _07110_);
  and (_07144_, _07143_, _07140_);
  and (_07145_, _07109_, word_in[25]);
  or (_26864_[1], _07145_, _07144_);
  not (_07146_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_07147_, _07115_, _07146_);
  and (_07149_, _07115_, _06519_);
  or (_07150_, _07149_, _07147_);
  or (_07151_, _07150_, _07111_);
  or (_07152_, _07112_, word_in[10]);
  and (_07153_, _07152_, _07151_);
  or (_07154_, _07153_, _07122_);
  or (_07155_, _07127_, _06514_);
  and (_07156_, _07155_, _07110_);
  and (_07157_, _07156_, _07154_);
  and (_07158_, _07109_, word_in[26]);
  or (_26864_[2], _07158_, _07157_);
  not (_07160_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_07161_, _07115_, _07160_);
  and (_07162_, _07115_, _06538_);
  or (_07163_, _07162_, _07161_);
  or (_07164_, _07163_, _07111_);
  or (_07165_, _07112_, word_in[11]);
  and (_07166_, _07165_, _07164_);
  or (_07167_, _07166_, _07122_);
  or (_07168_, _07127_, _06534_);
  and (_07170_, _07168_, _07110_);
  and (_07171_, _07170_, _07167_);
  and (_07172_, _07109_, word_in[27]);
  or (_26864_[3], _07172_, _07171_);
  not (_07174_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_07176_, _07115_, _07174_);
  and (_07177_, _07115_, _06554_);
  or (_07179_, _07177_, _07176_);
  and (_07180_, _07179_, _07112_);
  and (_07181_, _07111_, word_in[12]);
  or (_07182_, _07181_, _07180_);
  or (_07185_, _07182_, _07122_);
  or (_07186_, _07127_, _06549_);
  and (_07188_, _07186_, _07110_);
  and (_07190_, _07188_, _07185_);
  and (_07191_, _07109_, word_in[28]);
  or (_26864_[4], _07191_, _07190_);
  not (_07192_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_07193_, _07115_, _07192_);
  and (_07194_, _07115_, _06570_);
  or (_07196_, _07194_, _07193_);
  or (_07198_, _07196_, _07111_);
  or (_07199_, _07112_, word_in[13]);
  and (_07200_, _07199_, _07198_);
  or (_07201_, _07200_, _07122_);
  or (_07203_, _07127_, _06566_);
  and (_07204_, _07203_, _07110_);
  and (_07205_, _07204_, _07201_);
  and (_07207_, _07109_, word_in[29]);
  or (_26864_[5], _07207_, _07205_);
  not (_07209_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_07212_, _07115_, _07209_);
  and (_07214_, _07115_, _06585_);
  or (_07215_, _07214_, _07212_);
  or (_07216_, _07215_, _07111_);
  or (_07218_, _07112_, word_in[14]);
  and (_07220_, _07218_, _07216_);
  or (_07222_, _07220_, _07122_);
  or (_07223_, _07127_, _06580_);
  and (_07224_, _07223_, _07110_);
  and (_07225_, _07224_, _07222_);
  and (_07226_, _07109_, word_in[30]);
  or (_26864_[6], _07226_, _07225_);
  nor (_07227_, _07115_, _05671_);
  and (_07228_, _07115_, _05862_);
  or (_07229_, _07228_, _07227_);
  or (_07230_, _07229_, _07111_);
  or (_07231_, _07112_, word_in[15]);
  and (_07233_, _07231_, _07230_);
  or (_07234_, _07233_, _07122_);
  or (_07235_, _07127_, _05872_);
  and (_07236_, _07235_, _07110_);
  and (_07237_, _07236_, _07234_);
  and (_07238_, _07109_, word_in[31]);
  or (_26864_[7], _07238_, _07237_);
  and (_07240_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_07241_, _06040_, _23791_);
  or (_02136_, _07241_, _07240_);
  and (_07242_, _05846_, _05914_);
  not (_07243_, _07242_);
  and (_07244_, _06842_, _05622_);
  and (_07245_, _07244_, _06336_);
  and (_07246_, _05854_, _05670_);
  not (_07248_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_07250_, _06846_, _05857_);
  nor (_07251_, _07250_, _07248_);
  and (_07253_, _07250_, _06482_);
  nor (_07254_, _07253_, _07251_);
  nor (_07256_, _07254_, _07246_);
  and (_07257_, _07246_, word_in[8]);
  nor (_07258_, _07257_, _07256_);
  nor (_07259_, _07258_, _07244_);
  or (_07260_, _07259_, _07245_);
  and (_07261_, _07260_, _07243_);
  and (_07262_, _07242_, word_in[24]);
  or (_26865_[0], _07262_, _07261_);
  or (_07263_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_07264_, _07263_, _22761_);
  nand (_07265_, _23889_, _23832_);
  and (_02153_, _07265_, _07264_);
  and (_07266_, _07242_, word_in[25]);
  not (_07267_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_07268_, _07250_, _07267_);
  and (_07269_, _07250_, _06346_);
  or (_07270_, _07269_, _07268_);
  or (_07271_, _07270_, _07246_);
  not (_07272_, _07246_);
  or (_07274_, _07272_, word_in[9]);
  and (_07276_, _07274_, _07271_);
  or (_07278_, _07276_, _07244_);
  not (_07279_, _07244_);
  or (_07280_, _07279_, _06500_);
  and (_07281_, _07280_, _07243_);
  and (_07282_, _07281_, _07278_);
  or (_26865_[1], _07282_, _07266_);
  and (_07284_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and (_07285_, _06040_, _23676_);
  or (_27118_, _07285_, _07284_);
  and (_07286_, _07250_, _06519_);
  not (_07287_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_07288_, _07250_, _07287_);
  nor (_07289_, _07288_, _07286_);
  nor (_07290_, _07289_, _07246_);
  and (_07292_, _07246_, word_in[10]);
  nor (_07293_, _07292_, _07290_);
  nor (_07295_, _07293_, _07244_);
  and (_07296_, _07244_, _06514_);
  or (_07297_, _07296_, _07295_);
  and (_07299_, _07297_, _07243_);
  and (_07301_, _07242_, word_in[26]);
  or (_26865_[2], _07301_, _07299_);
  and (_07302_, _07242_, word_in[27]);
  not (_07303_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_07305_, _07250_, _07303_);
  and (_07306_, _07250_, _06538_);
  or (_07307_, _07306_, _07305_);
  or (_07308_, _07307_, _07246_);
  or (_07309_, _07272_, word_in[11]);
  and (_07310_, _07309_, _07308_);
  or (_07312_, _07310_, _07244_);
  or (_07313_, _07279_, _06534_);
  and (_07315_, _07313_, _07243_);
  and (_07317_, _07315_, _07312_);
  or (_26865_[3], _07317_, _07302_);
  and (_07319_, _07244_, _06549_);
  not (_07321_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_07322_, _07250_, _07321_);
  and (_07324_, _07250_, _06554_);
  nor (_07326_, _07324_, _07322_);
  nor (_07328_, _07326_, _07246_);
  and (_07329_, _07246_, word_in[12]);
  nor (_07331_, _07329_, _07328_);
  nor (_07332_, _07331_, _07244_);
  or (_07334_, _07332_, _07319_);
  and (_07336_, _07334_, _07243_);
  and (_07337_, _07242_, word_in[28]);
  or (_26865_[4], _07337_, _07336_);
  and (_07340_, _07250_, _06570_);
  not (_07341_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_07343_, _07250_, _07341_);
  nor (_07344_, _07343_, _07340_);
  nor (_07346_, _07344_, _07246_);
  and (_07348_, _07246_, word_in[13]);
  nor (_07349_, _07348_, _07346_);
  nor (_07351_, _07349_, _07244_);
  and (_07353_, _07244_, _06566_);
  or (_07354_, _07353_, _07351_);
  and (_07356_, _07354_, _07243_);
  and (_07357_, _07242_, word_in[29]);
  or (_26865_[5], _07357_, _07356_);
  or (_07359_, _07279_, _06580_);
  not (_07361_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_07363_, _07250_, _07361_);
  and (_07365_, _07250_, _06585_);
  or (_07366_, _07365_, _07363_);
  or (_07368_, _07366_, _07246_);
  or (_07369_, _07272_, word_in[14]);
  and (_07370_, _07369_, _07368_);
  or (_07371_, _07370_, _07244_);
  and (_07372_, _07371_, _07359_);
  and (_07373_, _07372_, _07243_);
  and (_07374_, _07242_, word_in[30]);
  or (_26865_[6], _07374_, _07373_);
  or (_07375_, _07279_, _05872_);
  nor (_07376_, _07250_, _05546_);
  and (_07377_, _07250_, _05862_);
  or (_07378_, _07377_, _07376_);
  or (_07379_, _07378_, _07246_);
  or (_07380_, _07272_, word_in[15]);
  and (_07381_, _07380_, _07379_);
  or (_07382_, _07381_, _07244_);
  and (_07383_, _07382_, _07375_);
  and (_07384_, _07383_, _07243_);
  and (_07385_, _07242_, word_in[31]);
  or (_26865_[7], _07385_, _07384_);
  and (_07386_, _06009_, _23838_);
  and (_07387_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_02219_, _07387_, _07386_);
  and (_07388_, _05846_, _05938_);
  not (_07389_, _07388_);
  and (_07390_, _05849_, _05955_);
  and (_07391_, _07390_, word_in[16]);
  and (_07392_, _05853_, _05604_);
  not (_07393_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_07394_, _05471_, _05511_);
  and (_07396_, _05858_, _07394_);
  and (_07397_, _07396_, _06317_);
  nor (_07398_, _07397_, _07393_);
  and (_07399_, _07397_, word_in[0]);
  or (_07400_, _07399_, _07398_);
  or (_07402_, _07400_, _07392_);
  not (_07405_, _07390_);
  not (_07406_, _07392_);
  or (_07407_, _07406_, word_in[8]);
  and (_07408_, _07407_, _07405_);
  and (_07410_, _07408_, _07402_);
  or (_07412_, _07410_, _07391_);
  and (_07413_, _07412_, _07389_);
  and (_07415_, _07388_, word_in[24]);
  or (_26866_[0], _07415_, _07413_);
  and (_07417_, _07388_, word_in[25]);
  not (_07419_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_07421_, _07397_, _07419_);
  and (_07422_, _07397_, _06346_);
  or (_07424_, _07422_, _07421_);
  and (_07425_, _07424_, _07406_);
  and (_07426_, _07392_, word_in[9]);
  or (_07427_, _07426_, _07425_);
  or (_07428_, _07427_, _07390_);
  or (_07429_, _07405_, word_in[17]);
  and (_07431_, _07429_, _07389_);
  and (_07433_, _07431_, _07428_);
  or (_26866_[1], _07433_, _07417_);
  and (_07435_, _07388_, word_in[26]);
  not (_07436_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_07438_, _07397_, _07436_);
  and (_07439_, _07397_, _06519_);
  or (_07440_, _07439_, _07438_);
  or (_07441_, _07440_, _07392_);
  or (_07443_, _07406_, word_in[10]);
  and (_07444_, _07443_, _07441_);
  or (_07446_, _07444_, _07390_);
  or (_07447_, _07405_, word_in[18]);
  and (_07449_, _07447_, _07389_);
  and (_07450_, _07449_, _07446_);
  or (_26866_[2], _07450_, _07435_);
  and (_07453_, _07388_, word_in[27]);
  not (_07455_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_07456_, _07397_, _07455_);
  and (_07457_, _07397_, word_in[3]);
  or (_07458_, _07457_, _07456_);
  and (_07459_, _07458_, _07406_);
  and (_07461_, _07392_, word_in[11]);
  or (_07462_, _07461_, _07459_);
  or (_07464_, _07462_, _07390_);
  or (_07466_, _07405_, word_in[19]);
  and (_07468_, _07466_, _07389_);
  and (_07469_, _07468_, _07464_);
  or (_26866_[3], _07469_, _07453_);
  and (_07472_, _07388_, word_in[28]);
  not (_07473_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_07474_, _07397_, _07473_);
  and (_07475_, _07397_, word_in[4]);
  or (_07476_, _07475_, _07474_);
  and (_07477_, _07476_, _07406_);
  and (_07478_, _07392_, word_in[12]);
  or (_07479_, _07478_, _07477_);
  or (_07480_, _07479_, _07390_);
  or (_07481_, _07405_, word_in[20]);
  and (_07482_, _07481_, _07389_);
  and (_07483_, _07482_, _07480_);
  or (_26866_[4], _07483_, _07472_);
  not (_07485_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_07486_, _07397_, _07485_);
  and (_07487_, _07397_, _06570_);
  or (_07488_, _07487_, _07486_);
  or (_07490_, _07488_, _07392_);
  or (_07491_, _07406_, word_in[13]);
  and (_07492_, _07491_, _07490_);
  or (_07493_, _07492_, _07390_);
  or (_07494_, _07405_, word_in[21]);
  and (_07496_, _07494_, _07493_);
  or (_07497_, _07496_, _07388_);
  or (_07498_, _07389_, word_in[29]);
  and (_26866_[5], _07498_, _07497_);
  not (_07500_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_07501_, _07397_, _07500_);
  and (_07502_, _07397_, word_in[6]);
  or (_07503_, _07502_, _07501_);
  and (_07504_, _07503_, _07406_);
  and (_07505_, _07392_, word_in[14]);
  or (_07506_, _07505_, _07504_);
  and (_07507_, _07506_, _07405_);
  and (_07508_, _07390_, word_in[22]);
  or (_07509_, _07508_, _07507_);
  and (_07510_, _07509_, _07389_);
  and (_07511_, _07388_, word_in[30]);
  or (_26866_[6], _07511_, _07510_);
  nor (_07512_, _07397_, _05647_);
  and (_07513_, _07397_, _05862_);
  or (_07515_, _07513_, _07512_);
  or (_07517_, _07515_, _07392_);
  or (_07518_, _07406_, word_in[15]);
  and (_07519_, _07518_, _07517_);
  or (_07520_, _07519_, _07390_);
  or (_07521_, _07405_, word_in[23]);
  and (_07522_, _07521_, _07389_);
  and (_07523_, _07522_, _07520_);
  and (_07524_, _07388_, word_in[31]);
  or (_26866_[7], _07524_, _07523_);
  and (_07525_, _06044_, _23718_);
  and (_07527_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_02258_, _07527_, _07525_);
  and (_07528_, _06009_, _23718_);
  and (_07529_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_02270_, _07529_, _07528_);
  and (_07530_, _05846_, _05955_);
  and (_07531_, _06475_, _05608_);
  not (_07532_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_07533_, _07396_, _06479_);
  nor (_07534_, _07533_, _07532_);
  and (_07535_, _07533_, _06482_);
  nor (_07536_, _07535_, _07534_);
  nor (_07537_, _07536_, _07531_);
  and (_07538_, _06487_, _05710_);
  and (_07539_, _07531_, word_in[8]);
  or (_07540_, _07539_, _07538_);
  or (_07541_, _07540_, _07537_);
  not (_07542_, _07538_);
  or (_07543_, _07542_, _06336_);
  and (_07545_, _07543_, _07541_);
  or (_07546_, _07545_, _07530_);
  not (_07548_, _07530_);
  or (_07549_, _07548_, word_in[24]);
  and (_26867_[0], _07549_, _07546_);
  or (_07550_, _07542_, _06500_);
  not (_07551_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_07553_, _07533_, _07551_);
  and (_07554_, _07533_, _06346_);
  nor (_07555_, _07554_, _07553_);
  nor (_07556_, _07555_, _07531_);
  and (_07557_, _07531_, word_in[9]);
  or (_07558_, _07557_, _07538_);
  or (_07559_, _07558_, _07556_);
  and (_07560_, _07559_, _07550_);
  or (_07561_, _07560_, _07530_);
  or (_07562_, _07548_, word_in[25]);
  and (_26867_[1], _07562_, _07561_);
  or (_07563_, _07542_, _06514_);
  not (_07564_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_07565_, _07533_, _07564_);
  and (_07566_, _07533_, _06519_);
  nor (_07567_, _07566_, _07565_);
  nor (_07568_, _07567_, _07531_);
  and (_07569_, _07531_, word_in[10]);
  or (_07570_, _07569_, _07538_);
  or (_07571_, _07570_, _07568_);
  and (_07572_, _07571_, _07563_);
  or (_07573_, _07572_, _07530_);
  or (_07574_, _07548_, word_in[26]);
  and (_26867_[2], _07574_, _07573_);
  or (_07575_, _07542_, _06534_);
  not (_07576_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_07577_, _07533_, _07576_);
  and (_07578_, _07533_, _06538_);
  nor (_07579_, _07578_, _07577_);
  nor (_07580_, _07579_, _07531_);
  and (_07581_, _07531_, word_in[11]);
  or (_07582_, _07581_, _07538_);
  or (_07583_, _07582_, _07580_);
  and (_07584_, _07583_, _07575_);
  or (_07586_, _07584_, _07530_);
  or (_07587_, _07548_, word_in[27]);
  and (_26867_[3], _07587_, _07586_);
  or (_07588_, _07542_, _06549_);
  not (_07589_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_07590_, _07533_, _07589_);
  and (_07591_, _07533_, _06554_);
  nor (_07592_, _07591_, _07590_);
  nor (_07593_, _07592_, _07531_);
  and (_07594_, _07531_, word_in[12]);
  or (_07595_, _07594_, _07538_);
  or (_07596_, _07595_, _07593_);
  and (_07597_, _07596_, _07588_);
  or (_07598_, _07597_, _07530_);
  or (_07599_, _07548_, word_in[28]);
  and (_26867_[4], _07599_, _07598_);
  or (_07600_, _07542_, _06566_);
  not (_07601_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_07602_, _07533_, _07601_);
  and (_07603_, _07533_, _06570_);
  nor (_07605_, _07603_, _07602_);
  nor (_07606_, _07605_, _07531_);
  and (_07607_, _07531_, word_in[13]);
  or (_07608_, _07607_, _07538_);
  or (_07609_, _07608_, _07606_);
  and (_07610_, _07609_, _07600_);
  or (_07611_, _07610_, _07530_);
  or (_07612_, _07548_, word_in[29]);
  and (_26867_[5], _07612_, _07611_);
  or (_07613_, _07542_, _06580_);
  not (_07614_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_07615_, _07533_, _07614_);
  and (_07616_, _07533_, _06585_);
  nor (_07617_, _07616_, _07615_);
  nor (_07618_, _07617_, _07531_);
  and (_07619_, _07531_, word_in[14]);
  or (_07620_, _07619_, _07538_);
  or (_07621_, _07620_, _07618_);
  and (_07622_, _07621_, _07613_);
  or (_07623_, _07622_, _07530_);
  or (_07625_, _07548_, word_in[30]);
  and (_26867_[6], _07625_, _07623_);
  or (_07626_, _07542_, _05872_);
  nor (_07627_, _07533_, _05564_);
  and (_07628_, _07533_, _05862_);
  nor (_07629_, _07628_, _07627_);
  nor (_07630_, _07629_, _07531_);
  and (_07631_, _07531_, word_in[15]);
  or (_07632_, _07631_, _07538_);
  or (_07633_, _07632_, _07630_);
  and (_07634_, _07633_, _07626_);
  or (_07635_, _07634_, _07530_);
  or (_07636_, _07548_, word_in[31]);
  and (_26867_[7], _07636_, _07635_);
  and (_07637_, _06607_, _05782_);
  and (_07638_, _06609_, _05710_);
  not (_07639_, _07638_);
  or (_07640_, _07639_, _06336_);
  and (_07641_, _06613_, _05608_);
  not (_07642_, _07641_);
  not (_07643_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_07644_, _07396_, _06618_);
  nor (_07645_, _07644_, _07643_);
  and (_07646_, _07644_, _06482_);
  or (_07647_, _07646_, _07645_);
  and (_07648_, _07647_, _07642_);
  and (_07649_, _07641_, word_in[8]);
  or (_07650_, _07649_, _07638_);
  or (_07651_, _07650_, _07648_);
  and (_07652_, _07651_, _07640_);
  or (_07653_, _07652_, _07637_);
  not (_07654_, _07637_);
  or (_07655_, _07654_, word_in[24]);
  and (_26853_[0], _07655_, _07653_);
  or (_07656_, _07639_, _06500_);
  not (_07657_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_07658_, _07644_, _07657_);
  and (_07659_, _07644_, _06346_);
  or (_07660_, _07659_, _07658_);
  and (_07661_, _07660_, _07642_);
  and (_07662_, _07641_, word_in[9]);
  or (_07663_, _07662_, _07638_);
  or (_07664_, _07663_, _07661_);
  and (_07665_, _07664_, _07656_);
  or (_07666_, _07665_, _07637_);
  or (_07667_, _07654_, word_in[25]);
  and (_26853_[1], _07667_, _07666_);
  not (_07668_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_07669_, _07644_, _07668_);
  and (_07670_, _07644_, _06519_);
  or (_07671_, _07670_, _07669_);
  and (_07672_, _07671_, _07642_);
  and (_07673_, _07641_, word_in[10]);
  or (_07674_, _07673_, _07638_);
  or (_07675_, _07674_, _07672_);
  or (_07676_, _07639_, _06514_);
  and (_07677_, _07676_, _07675_);
  or (_07678_, _07677_, _07637_);
  or (_07679_, _07654_, word_in[26]);
  and (_26853_[2], _07679_, _07678_);
  not (_07680_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_07681_, _07644_, _07680_);
  and (_07682_, _07644_, _06538_);
  or (_07683_, _07682_, _07681_);
  and (_07684_, _07683_, _07642_);
  and (_07685_, _07641_, word_in[11]);
  or (_07686_, _07685_, _07638_);
  or (_07687_, _07686_, _07684_);
  or (_07688_, _07639_, _06534_);
  and (_07689_, _07688_, _07687_);
  or (_07691_, _07689_, _07637_);
  or (_07692_, _07654_, word_in[27]);
  and (_26853_[3], _07692_, _07691_);
  or (_07693_, _07639_, _06549_);
  not (_07694_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_07695_, _07644_, _07694_);
  and (_07696_, _07644_, _06554_);
  or (_07697_, _07696_, _07695_);
  and (_07698_, _07697_, _07642_);
  and (_07699_, _07641_, word_in[12]);
  or (_07700_, _07699_, _07638_);
  or (_07701_, _07700_, _07698_);
  and (_07702_, _07701_, _07693_);
  or (_07703_, _07702_, _07637_);
  or (_07704_, _07654_, word_in[28]);
  and (_26853_[4], _07704_, _07703_);
  not (_07705_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_07706_, _07644_, _07705_);
  and (_07707_, _07644_, _06570_);
  or (_07708_, _07707_, _07706_);
  and (_07710_, _07708_, _07642_);
  and (_07711_, _07641_, word_in[13]);
  or (_07712_, _07711_, _07638_);
  or (_07713_, _07712_, _07710_);
  or (_07714_, _07639_, _06566_);
  and (_07715_, _07714_, _07713_);
  or (_07716_, _07715_, _07637_);
  or (_07717_, _07654_, word_in[29]);
  and (_26853_[5], _07717_, _07716_);
  not (_07718_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_07719_, _07644_, _07718_);
  and (_07720_, _07644_, _06585_);
  or (_07721_, _07720_, _07719_);
  and (_07722_, _07721_, _07642_);
  and (_07723_, _07641_, word_in[14]);
  or (_07724_, _07723_, _07638_);
  or (_07725_, _07724_, _07722_);
  or (_07726_, _07639_, _06580_);
  and (_07727_, _07726_, _07725_);
  and (_07728_, _07727_, _07654_);
  and (_07730_, _07637_, word_in[30]);
  or (_26853_[6], _07730_, _07728_);
  or (_07731_, _07639_, _05872_);
  nor (_07732_, _07644_, _05642_);
  and (_07733_, _07644_, _05862_);
  or (_07734_, _07733_, _07732_);
  and (_07735_, _07734_, _07642_);
  and (_07736_, _07641_, word_in[15]);
  or (_07737_, _07736_, _07638_);
  or (_07738_, _07737_, _07735_);
  and (_07739_, _07738_, _07731_);
  or (_07740_, _07739_, _07637_);
  or (_07741_, _07654_, word_in[31]);
  and (_26853_[7], _07741_, _07740_);
  and (_07742_, _05854_, _05608_);
  not (_07743_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_07744_, _07396_, _05857_);
  nor (_07745_, _07744_, _07743_);
  and (_07746_, _07744_, _06482_);
  nor (_07747_, _07746_, _07745_);
  nor (_07748_, _07747_, _07742_);
  and (_07749_, _06737_, _05710_);
  and (_07750_, _07742_, word_in[8]);
  or (_07751_, _07750_, _07749_);
  or (_07752_, _07751_, _07748_);
  and (_07753_, _05846_, _05999_);
  not (_07754_, _07753_);
  not (_07755_, _07749_);
  or (_07756_, _07755_, _06336_);
  and (_07757_, _07756_, _07754_);
  and (_07758_, _07757_, _07752_);
  and (_07759_, _07753_, word_in[24]);
  or (_26854_[0], _07759_, _07758_);
  and (_07760_, _07753_, word_in[25]);
  not (_07761_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_07762_, _07744_, _07761_);
  and (_07763_, _07744_, _06346_);
  nor (_07764_, _07763_, _07762_);
  nor (_07765_, _07764_, _07742_);
  and (_07766_, _07742_, word_in[9]);
  or (_07767_, _07766_, _07749_);
  or (_07768_, _07767_, _07765_);
  or (_07769_, _07755_, _06500_);
  and (_07770_, _07769_, _07754_);
  and (_07771_, _07770_, _07768_);
  or (_26854_[1], _07771_, _07760_);
  not (_07772_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_07773_, _07744_, _07772_);
  and (_07774_, _07744_, _06519_);
  nor (_07775_, _07774_, _07773_);
  nor (_07776_, _07775_, _07742_);
  and (_07777_, _07742_, word_in[10]);
  or (_07778_, _07777_, _07749_);
  or (_07779_, _07778_, _07776_);
  or (_07780_, _07755_, _06514_);
  and (_07781_, _07780_, _07754_);
  and (_07782_, _07781_, _07779_);
  and (_07784_, _07753_, word_in[26]);
  or (_26854_[2], _07784_, _07782_);
  and (_07785_, _07753_, word_in[27]);
  not (_07786_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_07788_, _07744_, _07786_);
  and (_07790_, _07744_, _06538_);
  nor (_07792_, _07790_, _07788_);
  nor (_07793_, _07792_, _07742_);
  and (_07794_, _07742_, word_in[11]);
  or (_07795_, _07794_, _07749_);
  or (_07796_, _07795_, _07793_);
  or (_07797_, _07755_, _06534_);
  and (_07798_, _07797_, _07754_);
  and (_07799_, _07798_, _07796_);
  or (_26854_[3], _07799_, _07785_);
  not (_07800_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_07801_, _07744_, _07800_);
  and (_07802_, _07744_, _06554_);
  nor (_07803_, _07802_, _07801_);
  nor (_07804_, _07803_, _07742_);
  and (_07806_, _07742_, word_in[12]);
  or (_07807_, _07806_, _07749_);
  or (_07808_, _07807_, _07804_);
  or (_07810_, _07755_, _06549_);
  and (_07811_, _07810_, _07754_);
  and (_07812_, _07811_, _07808_);
  and (_07813_, _07753_, word_in[28]);
  or (_26854_[4], _07813_, _07812_);
  not (_07814_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_07815_, _07744_, _07814_);
  and (_07817_, _07744_, _06570_);
  nor (_07818_, _07817_, _07815_);
  nor (_07820_, _07818_, _07742_);
  and (_07821_, _07742_, word_in[13]);
  or (_07822_, _07821_, _07749_);
  or (_07824_, _07822_, _07820_);
  or (_07825_, _07755_, _06566_);
  and (_07826_, _07825_, _07754_);
  and (_07827_, _07826_, _07824_);
  and (_07828_, _07753_, word_in[29]);
  or (_26854_[5], _07828_, _07827_);
  not (_07829_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_07830_, _07744_, _07829_);
  and (_07832_, _07744_, _06585_);
  nor (_07833_, _07832_, _07830_);
  nor (_07834_, _07833_, _07742_);
  and (_07835_, _07742_, word_in[14]);
  or (_07836_, _07835_, _07749_);
  or (_07837_, _07836_, _07834_);
  or (_07838_, _07755_, _06580_);
  and (_07839_, _07838_, _07754_);
  and (_07840_, _07839_, _07837_);
  and (_07841_, _07753_, word_in[30]);
  or (_26854_[6], _07841_, _07840_);
  nor (_07842_, _07744_, _05584_);
  and (_07843_, _07744_, _05862_);
  nor (_07844_, _07843_, _07842_);
  nor (_07845_, _07844_, _07742_);
  and (_07846_, _07742_, word_in[15]);
  or (_07847_, _07846_, _07749_);
  or (_07848_, _07847_, _07845_);
  or (_07849_, _07755_, _05872_);
  and (_07850_, _07849_, _07754_);
  and (_07851_, _07850_, _07848_);
  and (_07852_, _07753_, word_in[31]);
  or (_26854_[7], _07852_, _07851_);
  and (_07853_, _03015_, _23838_);
  and (_07854_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_02406_, _07854_, _07853_);
  and (_07855_, _24573_, _23982_);
  and (_07856_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or (_02417_, _07856_, _07855_);
  and (_07857_, _06255_, _23838_);
  and (_07858_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or (_02433_, _07858_, _07857_);
  and (_07859_, _06255_, _23791_);
  and (_07860_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or (_02435_, _07860_, _07859_);
  and (_07861_, _03233_, _23594_);
  and (_07863_, _07861_, _23635_);
  not (_07865_, _07861_);
  and (_07866_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_26995_, _07866_, _07863_);
  and (_07869_, _02342_, _23982_);
  and (_07870_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_02445_, _07870_, _07869_);
  and (_07871_, _02342_, _23718_);
  and (_07872_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_02448_, _07872_, _07871_);
  and (_07873_, _02237_, _23982_);
  and (_07875_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_27157_, _07875_, _07873_);
  and (_07876_, _02237_, _23718_);
  and (_07878_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_02455_, _07878_, _07876_);
  and (_07879_, _05851_, _05595_);
  not (_07880_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_07881_, _06317_, _05860_);
  nor (_07883_, _07881_, _07880_);
  and (_07884_, _07881_, _06482_);
  or (_07885_, _07884_, _07883_);
  and (_07886_, _05853_, _06114_);
  or (_07888_, _07886_, _07885_);
  not (_07889_, _07886_);
  or (_07891_, _07889_, word_in[8]);
  and (_07893_, _07891_, _07888_);
  or (_07894_, _07893_, _07879_);
  and (_07895_, _05846_, _05827_);
  and (_07897_, _07895_, _05622_);
  not (_07898_, _07897_);
  not (_07900_, _07879_);
  or (_07901_, _07900_, _06336_);
  and (_07903_, _07901_, _07898_);
  and (_07904_, _07903_, _07894_);
  and (_07905_, _05846_, word_in[24]);
  and (_07906_, _07897_, _07905_);
  or (_26855_[0], _07906_, _07904_);
  and (_07908_, _07861_, _23982_);
  and (_07910_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_02461_, _07910_, _07908_);
  not (_07911_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_07912_, _07881_, _07911_);
  and (_07913_, _07881_, _06346_);
  or (_07915_, _07913_, _07912_);
  or (_07917_, _07915_, _07886_);
  or (_07918_, _07889_, word_in[9]);
  and (_07919_, _07918_, _07917_);
  and (_07921_, _07919_, _07900_);
  and (_07922_, _07879_, _06500_);
  or (_07924_, _07922_, _07897_);
  or (_07926_, _07924_, _07921_);
  and (_07927_, _05846_, word_in[25]);
  or (_07928_, _07898_, _07927_);
  and (_26855_[1], _07928_, _07926_);
  and (_07929_, _03354_, _23589_);
  and (_07930_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_02464_, _07930_, _07929_);
  not (_07931_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_07932_, _07881_, _07931_);
  and (_07933_, _07881_, word_in[2]);
  or (_07935_, _07933_, _07932_);
  and (_07937_, _07935_, _07889_);
  and (_07938_, _07886_, word_in[10]);
  or (_07939_, _07938_, _07937_);
  or (_07940_, _07939_, _07879_);
  or (_07941_, _07900_, _06514_);
  and (_07942_, _07941_, _07898_);
  and (_07943_, _07942_, _07940_);
  and (_07944_, _05846_, word_in[26]);
  and (_07945_, _07897_, _07944_);
  or (_26855_[2], _07945_, _07943_);
  and (_07946_, _02289_, _23635_);
  and (_07947_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or (_02467_, _07947_, _07946_);
  not (_07948_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_07949_, _07881_, _07948_);
  and (_07950_, _07881_, word_in[3]);
  or (_07951_, _07950_, _07949_);
  and (_07952_, _07951_, _07889_);
  and (_07953_, _07886_, word_in[11]);
  or (_07954_, _07953_, _07952_);
  or (_07955_, _07954_, _07879_);
  or (_07956_, _07900_, _06534_);
  and (_07958_, _07956_, _07898_);
  and (_07959_, _07958_, _07955_);
  and (_07960_, _05846_, word_in[27]);
  and (_07961_, _07897_, _07960_);
  or (_26855_[3], _07961_, _07959_);
  and (_07962_, _02289_, _23838_);
  and (_07963_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or (_02470_, _07963_, _07962_);
  not (_07964_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_07965_, _07881_, _07964_);
  and (_07966_, _07881_, word_in[4]);
  or (_07967_, _07966_, _07965_);
  and (_07968_, _07967_, _07889_);
  and (_07969_, _07886_, word_in[12]);
  or (_07970_, _07969_, _07968_);
  or (_07971_, _07970_, _07879_);
  or (_07972_, _07900_, _06549_);
  and (_07973_, _07972_, _07898_);
  and (_07974_, _07973_, _07971_);
  and (_07975_, _05846_, word_in[28]);
  and (_07977_, _07897_, _07975_);
  or (_26855_[4], _07977_, _07974_);
  not (_07978_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_07979_, _07881_, _07978_);
  and (_07980_, _07881_, word_in[5]);
  or (_07981_, _07980_, _07979_);
  and (_07982_, _07981_, _07889_);
  and (_07983_, _07886_, word_in[13]);
  or (_07984_, _07983_, _07982_);
  and (_07985_, _07984_, _07900_);
  and (_07986_, _07879_, _06566_);
  or (_07987_, _07986_, _07985_);
  and (_07988_, _07987_, _07898_);
  and (_07989_, _07897_, _06412_);
  or (_26855_[5], _07989_, _07988_);
  and (_07990_, _02318_, _23589_);
  and (_07991_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_02476_, _07991_, _07990_);
  not (_07992_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_07993_, _07881_, _07992_);
  and (_07994_, _07881_, _06585_);
  or (_07995_, _07994_, _07993_);
  or (_07996_, _07995_, _07886_);
  or (_07997_, _07889_, word_in[14]);
  and (_07998_, _07997_, _07996_);
  or (_07999_, _07998_, _07879_);
  or (_08000_, _07900_, _06580_);
  and (_08001_, _08000_, _07999_);
  or (_08002_, _08001_, _07897_);
  and (_08003_, _05846_, word_in[30]);
  or (_08004_, _07898_, _08003_);
  and (_26855_[6], _08004_, _08002_);
  nor (_08005_, _07881_, _05690_);
  and (_08006_, _07881_, word_in[7]);
  or (_08007_, _08006_, _08005_);
  and (_08008_, _08007_, _07889_);
  and (_08009_, _07886_, word_in[15]);
  or (_08010_, _08009_, _08008_);
  or (_08011_, _08010_, _07879_);
  or (_08012_, _07900_, _05872_);
  and (_08013_, _08012_, _07898_);
  and (_08014_, _08013_, _08011_);
  and (_08015_, _05846_, word_in[31]);
  and (_08016_, _07897_, _08015_);
  or (_26855_[7], _08016_, _08014_);
  and (_08017_, _02318_, _23718_);
  and (_08018_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_02489_, _08018_, _08017_);
  and (_08019_, _02383_, _23838_);
  and (_08020_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or (_02507_, _08020_, _08019_);
  and (_08022_, _02779_, _23791_);
  and (_08023_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_02511_, _08023_, _08022_);
  and (_08024_, _02914_, _23755_);
  and (_08025_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_02515_, _08025_, _08024_);
  and (_08026_, _02914_, _23718_);
  and (_08027_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_02523_, _08027_, _08026_);
  and (_08028_, _02914_, _23676_);
  and (_08029_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_02529_, _08029_, _08028_);
  and (_08030_, _04704_, _23589_);
  and (_08031_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or (_27146_, _08031_, _08030_);
  and (_08032_, _04704_, _23982_);
  and (_08033_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or (_02534_, _08033_, _08032_);
  and (_08034_, _05329_, _23635_);
  and (_08035_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or (_02541_, _08035_, _08034_);
  and (_08036_, _07895_, _05595_);
  not (_08037_, _08036_);
  and (_08038_, _05851_, _05597_);
  and (_08039_, _08038_, _06336_);
  and (_08040_, _06475_, _05684_);
  and (_08041_, _06479_, _05860_);
  and (_08042_, _08041_, _06482_);
  not (_08043_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_08044_, _08041_, _08043_);
  nor (_08045_, _08044_, _08042_);
  nor (_08046_, _08045_, _08040_);
  and (_08047_, _08040_, word_in[8]);
  nor (_08048_, _08047_, _08046_);
  nor (_08049_, _08048_, _08038_);
  or (_08050_, _08049_, _08039_);
  and (_08051_, _08050_, _08037_);
  and (_08052_, _08036_, _07905_);
  or (_26856_[0], _08052_, _08051_);
  not (_08053_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_08054_, _08041_, _08053_);
  and (_08055_, _08041_, _06346_);
  or (_08056_, _08055_, _08054_);
  or (_08057_, _08056_, _08040_);
  not (_08058_, _08040_);
  or (_08059_, _08058_, word_in[9]);
  and (_08060_, _08059_, _08057_);
  or (_08061_, _08060_, _08038_);
  not (_08062_, _08038_);
  or (_08064_, _08062_, _06500_);
  and (_08065_, _08064_, _08061_);
  or (_08066_, _08065_, _08036_);
  or (_08067_, _08037_, _07927_);
  and (_26856_[1], _08067_, _08066_);
  and (_08068_, _03354_, _23755_);
  and (_08069_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_02551_, _08069_, _08068_);
  and (_08070_, _08038_, _06514_);
  and (_08071_, _08041_, _06519_);
  not (_08072_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_08073_, _08041_, _08072_);
  nor (_08074_, _08073_, _08071_);
  nor (_08075_, _08074_, _08040_);
  and (_08076_, _08040_, word_in[10]);
  nor (_08077_, _08076_, _08075_);
  nor (_08078_, _08077_, _08038_);
  or (_08079_, _08078_, _08070_);
  and (_08080_, _08079_, _08037_);
  and (_08081_, _08036_, _07944_);
  or (_26856_[2], _08081_, _08080_);
  and (_08083_, _05329_, _23676_);
  and (_08084_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or (_02555_, _08084_, _08083_);
  not (_08085_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_08086_, _08041_, _08085_);
  and (_08087_, _08041_, _06538_);
  or (_08088_, _08087_, _08086_);
  or (_08089_, _08088_, _08040_);
  or (_08090_, _08058_, word_in[11]);
  and (_08091_, _08090_, _08089_);
  or (_08092_, _08091_, _08038_);
  or (_08093_, _08062_, _06534_);
  and (_08094_, _08093_, _08092_);
  or (_08095_, _08094_, _08036_);
  or (_08096_, _08037_, _07960_);
  and (_26856_[3], _08096_, _08095_);
  and (_08097_, _08041_, _06554_);
  not (_08098_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_08099_, _08041_, _08098_);
  nor (_08100_, _08099_, _08097_);
  nor (_08101_, _08100_, _08040_);
  and (_08102_, _08040_, word_in[12]);
  nor (_08103_, _08102_, _08101_);
  nor (_08104_, _08103_, _08038_);
  and (_08105_, _08038_, _06549_);
  or (_08106_, _08105_, _08036_);
  or (_08107_, _08106_, _08104_);
  or (_08108_, _08037_, _07975_);
  and (_26856_[4], _08108_, _08107_);
  and (_08109_, _08041_, _06570_);
  not (_08110_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_08111_, _08041_, _08110_);
  nor (_08112_, _08111_, _08109_);
  nor (_08113_, _08112_, _08040_);
  and (_08114_, _08040_, word_in[13]);
  nor (_08115_, _08114_, _08113_);
  nor (_08116_, _08115_, _08038_);
  and (_08117_, _08038_, _06566_);
  or (_08118_, _08117_, _08036_);
  or (_08119_, _08118_, _08116_);
  or (_08120_, _08037_, _06412_);
  and (_26856_[5], _08120_, _08119_);
  not (_08121_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_08122_, _08041_, _08121_);
  and (_08123_, _08041_, _06585_);
  or (_08124_, _08123_, _08122_);
  or (_08125_, _08124_, _08040_);
  or (_08126_, _08058_, word_in[14]);
  and (_08127_, _08126_, _08125_);
  or (_08128_, _08127_, _08038_);
  or (_08129_, _08062_, _06580_);
  and (_08130_, _08129_, _08128_);
  or (_08131_, _08130_, _08036_);
  or (_08132_, _08037_, _08003_);
  and (_26856_[6], _08132_, _08131_);
  and (_08133_, _25517_, _23982_);
  and (_08134_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_27267_, _08134_, _08133_);
  nor (_08135_, _08041_, _05570_);
  and (_08136_, _08041_, _05862_);
  or (_08137_, _08136_, _08135_);
  or (_08138_, _08137_, _08040_);
  or (_08139_, _08058_, word_in[15]);
  and (_08140_, _08139_, _08138_);
  and (_08141_, _08140_, _08062_);
  and (_08142_, _08038_, _05872_);
  or (_08143_, _08142_, _08036_);
  or (_08144_, _08143_, _08141_);
  or (_08145_, _08037_, _08015_);
  and (_26856_[7], _08145_, _08144_);
  and (_08146_, _02937_, _23838_);
  and (_08147_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or (_02569_, _08147_, _08146_);
  and (_08148_, _02779_, _23755_);
  and (_08149_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_02574_, _08149_, _08148_);
  and (_08150_, _02937_, _23791_);
  and (_08151_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or (_02577_, _08151_, _08150_);
  and (_08152_, _03015_, _23676_);
  and (_08153_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_02584_, _08153_, _08152_);
  and (_08154_, _24573_, _23791_);
  and (_08155_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or (_27163_, _08155_, _08154_);
  and (_08156_, _06255_, _23635_);
  and (_08157_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or (_02597_, _08157_, _08156_);
  and (_08158_, _02342_, _23755_);
  and (_08159_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_02600_, _08159_, _08158_);
  and (_08162_, _02237_, _23755_);
  and (_08164_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_02605_, _08164_, _08162_);
  and (_08165_, _02289_, _23589_);
  and (_08166_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or (_02612_, _08166_, _08165_);
  and (_08168_, _02318_, _23982_);
  and (_08169_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_02617_, _08169_, _08168_);
  and (_08171_, _02318_, _23676_);
  and (_08173_, _02320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_02620_, _08173_, _08171_);
  and (_08174_, _02383_, _23635_);
  and (_08176_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or (_27154_, _08176_, _08174_);
  and (_08178_, _05851_, _05613_);
  and (_08179_, _06613_, _05684_);
  not (_08180_, _08179_);
  not (_08182_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_08183_, _06618_, _05839_);
  nor (_08185_, _08183_, _08182_);
  and (_08186_, _08183_, _06482_);
  or (_08187_, _08186_, _08185_);
  and (_08188_, _08187_, _08180_);
  and (_08190_, _08179_, word_in[8]);
  or (_08191_, _08190_, _08188_);
  or (_08192_, _08191_, _08178_);
  and (_08193_, _07895_, _05597_);
  not (_08194_, _08193_);
  not (_08195_, _08178_);
  or (_08197_, _08195_, _06336_);
  and (_08198_, _08197_, _08194_);
  and (_08199_, _08198_, _08192_);
  and (_08200_, _08193_, _07905_);
  or (_26857_[0], _08200_, _08199_);
  and (_08202_, _02779_, _23838_);
  and (_08204_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_02627_, _08204_, _08202_);
  not (_08205_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_08206_, _08183_, _08205_);
  and (_08207_, _08183_, _06346_);
  or (_08208_, _08207_, _08206_);
  and (_08209_, _08208_, _08180_);
  and (_08210_, _08179_, word_in[9]);
  or (_08211_, _08210_, _08209_);
  or (_08212_, _08211_, _08178_);
  or (_08213_, _08195_, _06500_);
  and (_08214_, _08213_, _08194_);
  and (_08215_, _08214_, _08212_);
  and (_08216_, _08193_, _07927_);
  or (_26857_[1], _08216_, _08215_);
  not (_08217_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_08218_, _08183_, _08217_);
  and (_08219_, _08183_, _06519_);
  or (_08220_, _08219_, _08218_);
  and (_08221_, _08220_, _08180_);
  and (_08222_, _08179_, word_in[10]);
  or (_08223_, _08222_, _08221_);
  or (_08225_, _08223_, _08178_);
  or (_08226_, _08195_, _06514_);
  and (_08227_, _08226_, _08194_);
  and (_08228_, _08227_, _08225_);
  and (_08229_, _08193_, _07944_);
  or (_26857_[2], _08229_, _08228_);
  and (_08230_, _02914_, _23982_);
  and (_08231_, _02916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_02631_, _08231_, _08230_);
  not (_08232_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_08233_, _08183_, _08232_);
  and (_08234_, _08183_, _06538_);
  or (_08235_, _08234_, _08233_);
  or (_08236_, _08235_, _08179_);
  or (_08237_, _08180_, word_in[11]);
  and (_08238_, _08237_, _08236_);
  or (_08239_, _08238_, _08178_);
  or (_08240_, _08195_, _06534_);
  and (_08241_, _08240_, _08194_);
  and (_08242_, _08241_, _08239_);
  and (_08243_, _08193_, _07960_);
  or (_26857_[3], _08243_, _08242_);
  not (_08244_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_08245_, _08183_, _08244_);
  and (_08246_, _08183_, _06554_);
  or (_08247_, _08246_, _08245_);
  and (_08248_, _08247_, _08180_);
  and (_08249_, _08179_, word_in[12]);
  or (_08250_, _08249_, _08248_);
  or (_08251_, _08250_, _08178_);
  or (_08252_, _08195_, _06549_);
  and (_08253_, _08252_, _08194_);
  and (_08254_, _08253_, _08251_);
  and (_08255_, _08193_, _07975_);
  or (_26857_[4], _08255_, _08254_);
  not (_08257_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_08258_, _08183_, _08257_);
  and (_08259_, _08183_, _06570_);
  or (_08260_, _08259_, _08258_);
  and (_08261_, _08260_, _08180_);
  and (_08262_, _08179_, word_in[13]);
  or (_08263_, _08262_, _08261_);
  or (_08264_, _08263_, _08178_);
  or (_08265_, _08195_, _06566_);
  and (_08266_, _08265_, _08194_);
  and (_08267_, _08266_, _08264_);
  and (_08268_, _08193_, _06412_);
  or (_26857_[5], _08268_, _08267_);
  and (_08269_, _04704_, _23791_);
  and (_08270_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or (_02637_, _08270_, _08269_);
  not (_08271_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_08272_, _08183_, _08271_);
  and (_08273_, _08183_, _06585_);
  or (_08274_, _08273_, _08272_);
  and (_08275_, _08274_, _08180_);
  and (_08276_, _08179_, word_in[14]);
  or (_08277_, _08276_, _08275_);
  or (_08278_, _08277_, _08178_);
  or (_08279_, _08195_, _06580_);
  and (_08280_, _08279_, _08194_);
  and (_08281_, _08280_, _08278_);
  and (_08282_, _08193_, _08003_);
  or (_26857_[6], _08282_, _08281_);
  and (_08283_, _06081_, _23982_);
  and (_08284_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or (_02641_, _08284_, _08283_);
  nor (_08285_, _08183_, _05685_);
  and (_08286_, _08183_, _05862_);
  or (_08287_, _08286_, _08285_);
  or (_08288_, _08287_, _08179_);
  or (_08289_, _08180_, word_in[15]);
  and (_08290_, _08289_, _08288_);
  or (_08291_, _08290_, _08178_);
  or (_08292_, _08195_, _05872_);
  and (_08293_, _08292_, _08291_);
  or (_08294_, _08293_, _08193_);
  or (_08296_, _08194_, _08015_);
  and (_26857_[7], _08296_, _08294_);
  and (_08297_, _07861_, _23589_);
  and (_08298_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_02648_, _08298_, _08297_);
  and (_08299_, _05329_, _23718_);
  and (_08300_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or (_02653_, _08300_, _08299_);
  and (_08302_, _02383_, _23676_);
  and (_08303_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or (_02657_, _08303_, _08302_);
  and (_08304_, _02937_, _23635_);
  and (_08305_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or (_02661_, _08305_, _08304_);
  and (_08306_, _03015_, _23982_);
  and (_08307_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_27165_, _08307_, _08306_);
  and (_08308_, _24573_, _23635_);
  and (_08309_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or (_27164_, _08309_, _08308_);
  and (_08310_, _07861_, _23755_);
  and (_08311_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_26996_, _08311_, _08310_);
  and (_08312_, _04704_, _23635_);
  and (_08313_, _04706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or (_27145_, _08313_, _08312_);
  and (_08314_, _05329_, _23755_);
  and (_08315_, _05331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or (_27144_, _08315_, _08314_);
  and (_08316_, _06264_, _23676_);
  and (_08317_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_26975_, _08317_, _08316_);
  and (_08318_, _07905_, _05847_);
  and (_08319_, _06482_, _05861_);
  not (_08320_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_08321_, _05861_, _08320_);
  nor (_08322_, _08321_, _08319_);
  nor (_08323_, _08322_, _05855_);
  and (_08324_, _05855_, word_in[8]);
  nor (_08325_, _08324_, _08323_);
  nor (_08326_, _08325_, _05852_);
  and (_08327_, _06336_, _05852_);
  or (_08328_, _08327_, _08326_);
  and (_08329_, _08328_, _05848_);
  or (_26858_[0], _08329_, _08318_);
  and (_08330_, _06255_, _23755_);
  and (_08331_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or (_27160_, _08331_, _08330_);
  and (_08332_, _07927_, _05847_);
  and (_08333_, _06346_, _05861_);
  not (_08334_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_08335_, _05861_, _08334_);
  nor (_08336_, _08335_, _08333_);
  nor (_08338_, _08336_, _05855_);
  and (_08339_, _05855_, word_in[9]);
  nor (_08340_, _08339_, _08338_);
  nor (_08341_, _08340_, _05852_);
  and (_08342_, _06500_, _05852_);
  or (_08343_, _08342_, _08341_);
  and (_08344_, _08343_, _05848_);
  or (_26858_[1], _08344_, _08332_);
  and (_08345_, _02237_, _23589_);
  and (_08346_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_27158_, _08346_, _08345_);
  and (_08347_, _07944_, _05847_);
  and (_08348_, _06519_, _05861_);
  not (_08349_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_08350_, _05861_, _08349_);
  nor (_08351_, _08350_, _08348_);
  nor (_08352_, _08351_, _05855_);
  and (_08353_, _05855_, word_in[10]);
  nor (_08354_, _08353_, _08352_);
  nor (_08355_, _08354_, _05852_);
  and (_08356_, _06514_, _05852_);
  or (_08357_, _08356_, _08355_);
  and (_08358_, _08357_, _05848_);
  or (_26858_[2], _08358_, _08347_);
  and (_08359_, _02289_, _23676_);
  and (_08360_, _02291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or (_27155_, _08360_, _08359_);
  and (_08361_, _07960_, _05847_);
  and (_08362_, _06538_, _05861_);
  not (_08363_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_08364_, _05861_, _08363_);
  nor (_08365_, _08364_, _08362_);
  nor (_08366_, _08365_, _05855_);
  and (_08367_, _05855_, word_in[11]);
  or (_08368_, _08367_, _08366_);
  or (_08369_, _08368_, _05852_);
  not (_08370_, _05852_);
  or (_08371_, _06534_, _08370_);
  and (_08372_, _08371_, _05848_);
  and (_08373_, _08372_, _08369_);
  or (_26858_[3], _08373_, _08361_);
  and (_08375_, _02779_, _23982_);
  and (_08376_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_27148_, _08376_, _08375_);
  and (_08377_, _07975_, _05847_);
  and (_08378_, _06554_, _05861_);
  not (_08379_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_08380_, _05861_, _08379_);
  nor (_08381_, _08380_, _08378_);
  nor (_08382_, _08381_, _05855_);
  and (_08383_, _05855_, word_in[12]);
  nor (_08384_, _08383_, _08382_);
  nor (_08385_, _08384_, _05852_);
  and (_08386_, _06549_, _05852_);
  or (_08387_, _08386_, _08385_);
  and (_08388_, _08387_, _05848_);
  or (_26858_[4], _08388_, _08377_);
  and (_08389_, _06412_, _05847_);
  and (_08390_, _06570_, _05861_);
  not (_08391_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_08393_, _05861_, _08391_);
  nor (_08394_, _08393_, _08390_);
  nor (_08395_, _08394_, _05855_);
  and (_08396_, _05855_, word_in[13]);
  or (_08397_, _08396_, _08395_);
  or (_08398_, _08397_, _05852_);
  or (_08399_, _06566_, _08370_);
  and (_08400_, _08399_, _05848_);
  and (_08401_, _08400_, _08398_);
  or (_26858_[5], _08401_, _08389_);
  and (_08402_, _02383_, _23791_);
  and (_08403_, _02385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or (_27153_, _08403_, _08402_);
  and (_08404_, _08003_, _05847_);
  and (_08405_, _06585_, _05861_);
  not (_08406_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_08407_, _05861_, _08406_);
  nor (_08408_, _08407_, _08405_);
  nor (_08409_, _08408_, _05855_);
  and (_08410_, _05855_, word_in[14]);
  nor (_08412_, _08410_, _08409_);
  nor (_08413_, _08412_, _05852_);
  and (_08414_, _06580_, _05852_);
  or (_08415_, _08414_, _08413_);
  and (_08416_, _08415_, _05848_);
  or (_26858_[6], _08416_, _08404_);
  and (_08417_, _03015_, _23635_);
  and (_08418_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_27166_, _08418_, _08417_);
  and (_08419_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and (_08420_, _06296_, _23718_);
  or (_27043_, _08420_, _08419_);
  and (_08421_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  and (_08422_, _06296_, _23635_);
  or (_27045_, _08422_, _08421_);
  and (_08423_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and (_08424_, _06296_, _23755_);
  or (_27046_, _08424_, _08423_);
  and (_08425_, _24567_, _23791_);
  and (_08426_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or (_27085_, _08426_, _08425_);
  and (_08427_, _24558_, _23863_);
  not (_08428_, _08427_);
  and (_08429_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_08430_, _08427_, _23676_);
  or (_27048_, _08430_, _08429_);
  and (_08431_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  and (_08432_, _03641_, _23838_);
  or (_27120_, _08432_, _08431_);
  and (_08433_, _06081_, _23838_);
  and (_08434_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or (_27265_, _08434_, _08433_);
  and (_08435_, _05537_, word_in[0]);
  nand (_08436_, _05455_, _06478_);
  or (_08437_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_08438_, _08437_, _08436_);
  and (_08439_, _08438_, _05497_);
  or (_08440_, _08439_, _05459_);
  nand (_08441_, _05455_, _06979_);
  or (_08442_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_08443_, _08442_, _08441_);
  and (_08444_, _08443_, _05473_);
  nand (_08445_, _05455_, _07248_);
  or (_08446_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_08447_, _08446_, _08445_);
  and (_08448_, _08447_, _05484_);
  nand (_08449_, _05455_, _06731_);
  or (_08450_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_08451_, _08450_, _08449_);
  and (_08452_, _08451_, _05477_);
  or (_08454_, _08452_, _08448_);
  or (_08455_, _08454_, _08444_);
  or (_08456_, _08455_, _08440_);
  nand (_08457_, _05455_, _07532_);
  or (_08458_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_08459_, _08458_, _08457_);
  and (_08460_, _08459_, _05497_);
  or (_08461_, _08460_, _05511_);
  nand (_08462_, _05455_, _08043_);
  or (_08463_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_08465_, _08463_, _08462_);
  and (_08466_, _08465_, _05473_);
  nand (_08467_, _05455_, _08320_);
  or (_08468_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_08469_, _08468_, _08467_);
  and (_08470_, _08469_, _05484_);
  nand (_08471_, _05455_, _07743_);
  or (_08472_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_08473_, _08472_, _08471_);
  and (_08474_, _08473_, _05477_);
  or (_08476_, _08474_, _08470_);
  or (_08477_, _08476_, _08466_);
  or (_08478_, _08477_, _08461_);
  and (_08479_, _08478_, _08456_);
  and (_08480_, _08479_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _08480_, _08435_);
  and (_08481_, _05537_, word_in[1]);
  nand (_08482_, _05455_, _06502_);
  or (_08483_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_08484_, _08483_, _08482_);
  and (_08485_, _08484_, _05497_);
  or (_08486_, _08485_, _05459_);
  nand (_08487_, _05455_, _07000_);
  or (_08488_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_08489_, _08488_, _08487_);
  and (_08490_, _08489_, _05473_);
  nand (_08491_, _05455_, _07267_);
  or (_08492_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_08493_, _08492_, _08491_);
  and (_08494_, _08493_, _05484_);
  nand (_08495_, _05455_, _06751_);
  or (_08496_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_08497_, _08496_, _08495_);
  and (_08498_, _08497_, _05477_);
  or (_08499_, _08498_, _08494_);
  or (_08501_, _08499_, _08490_);
  or (_08502_, _08501_, _08486_);
  nand (_08503_, _05455_, _07551_);
  or (_08504_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_08505_, _08504_, _08503_);
  and (_08506_, _08505_, _05497_);
  or (_08508_, _08506_, _05511_);
  nand (_08509_, _05455_, _08334_);
  or (_08511_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_08512_, _08511_, _08509_);
  and (_08513_, _08512_, _05484_);
  nand (_08514_, _05455_, _08053_);
  or (_08515_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_08516_, _08515_, _08514_);
  and (_08518_, _08516_, _05473_);
  or (_08519_, _08518_, _08513_);
  nand (_08520_, _05455_, _07761_);
  or (_08521_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_08522_, _08521_, _08520_);
  and (_08523_, _08522_, _05477_);
  or (_08524_, _08523_, _08519_);
  or (_08525_, _08524_, _08508_);
  and (_08526_, _08525_, _08502_);
  and (_08527_, _08526_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _08527_, _08481_);
  and (_08528_, _05537_, word_in[2]);
  nand (_08530_, _05455_, _06516_);
  or (_08531_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_08532_, _08531_, _08530_);
  and (_08533_, _08532_, _05497_);
  or (_08534_, _08533_, _05459_);
  nand (_08535_, _05455_, _07016_);
  or (_08536_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_08537_, _08536_, _08535_);
  and (_08538_, _08537_, _05473_);
  nand (_08540_, _05455_, _07287_);
  or (_08541_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_08542_, _08541_, _08540_);
  and (_08544_, _08542_, _05484_);
  nand (_08545_, _05455_, _06766_);
  or (_08546_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_08547_, _08546_, _08545_);
  and (_08548_, _08547_, _05477_);
  or (_08549_, _08548_, _08544_);
  or (_08550_, _08549_, _08538_);
  or (_08551_, _08550_, _08534_);
  nand (_08553_, _05455_, _07564_);
  or (_08554_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_08555_, _08554_, _08553_);
  and (_08556_, _08555_, _05497_);
  or (_08557_, _08556_, _05511_);
  nand (_08558_, _05455_, _08349_);
  or (_08559_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_08560_, _08559_, _08558_);
  and (_08561_, _08560_, _05484_);
  nand (_08563_, _05455_, _08072_);
  or (_08564_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_08565_, _08564_, _08563_);
  and (_08566_, _08565_, _05473_);
  or (_08567_, _08566_, _08561_);
  nand (_08568_, _05455_, _07772_);
  or (_08569_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_08571_, _08569_, _08568_);
  and (_08572_, _08571_, _05477_);
  or (_08573_, _08572_, _08567_);
  or (_08575_, _08573_, _08557_);
  and (_08576_, _08575_, _08551_);
  and (_08577_, _08576_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _08577_, _08528_);
  and (_08578_, _05537_, word_in[3]);
  nand (_08579_, _05455_, _06536_);
  or (_08580_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_08581_, _08580_, _08579_);
  and (_08582_, _08581_, _05497_);
  or (_08583_, _08582_, _05459_);
  nand (_08584_, _05455_, _07033_);
  or (_08585_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_08586_, _08585_, _08584_);
  and (_08587_, _08586_, _05473_);
  nand (_08588_, _05455_, _07303_);
  or (_08589_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_08590_, _08589_, _08588_);
  and (_08591_, _08590_, _05484_);
  nand (_08592_, _05455_, _06779_);
  or (_08594_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_08596_, _08594_, _08592_);
  and (_08597_, _08596_, _05477_);
  or (_08598_, _08597_, _08591_);
  or (_08599_, _08598_, _08587_);
  or (_08600_, _08599_, _08583_);
  nand (_08601_, _05455_, _07576_);
  or (_08602_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_08603_, _08602_, _08601_);
  and (_08604_, _08603_, _05497_);
  or (_08605_, _08604_, _05511_);
  nand (_08606_, _05455_, _08085_);
  or (_08608_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_08610_, _08608_, _08606_);
  and (_08611_, _08610_, _05473_);
  nand (_08612_, _05455_, _08363_);
  or (_08613_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_08614_, _08613_, _08612_);
  and (_08615_, _08614_, _05484_);
  nand (_08616_, _05455_, _07786_);
  or (_08617_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_08618_, _08617_, _08616_);
  and (_08619_, _08618_, _05477_);
  or (_08620_, _08619_, _08615_);
  or (_08621_, _08620_, _08611_);
  or (_08622_, _08621_, _08605_);
  and (_08623_, _08622_, _08600_);
  and (_08624_, _08623_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _08624_, _08578_);
  and (_08625_, _05537_, word_in[4]);
  nand (_08626_, _05455_, _06792_);
  or (_08628_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_08629_, _08628_, _08626_);
  and (_08630_, _08629_, _05477_);
  or (_08631_, _08630_, _05459_);
  nand (_08632_, _05455_, _07047_);
  or (_08633_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_08634_, _08633_, _08632_);
  and (_08635_, _08634_, _05473_);
  nand (_08636_, _05455_, _07321_);
  or (_08637_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_08638_, _08637_, _08636_);
  and (_08639_, _08638_, _05484_);
  nand (_08640_, _05455_, _06551_);
  or (_08641_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_08642_, _08641_, _08640_);
  and (_08643_, _08642_, _05497_);
  or (_08644_, _08643_, _08639_);
  or (_08645_, _08644_, _08635_);
  or (_08646_, _08645_, _08631_);
  nand (_08647_, _05455_, _07800_);
  or (_08648_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_08649_, _08648_, _08647_);
  and (_08650_, _08649_, _05477_);
  or (_08651_, _08650_, _05511_);
  nand (_08652_, _05455_, _08379_);
  or (_08653_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_08654_, _08653_, _08652_);
  and (_08655_, _08654_, _05484_);
  nand (_08656_, _05455_, _08098_);
  or (_08657_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_08659_, _08657_, _08656_);
  and (_08660_, _08659_, _05473_);
  or (_08661_, _08660_, _08655_);
  nand (_08662_, _05455_, _07589_);
  or (_08663_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_08664_, _08663_, _08662_);
  and (_08665_, _08664_, _05497_);
  or (_08666_, _08665_, _08661_);
  or (_08667_, _08666_, _08651_);
  and (_08668_, _08667_, _08646_);
  and (_08669_, _08668_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _08669_, _08625_);
  and (_08670_, _05537_, word_in[5]);
  nand (_08671_, _05455_, _06804_);
  or (_08672_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_08673_, _08672_, _08671_);
  and (_08674_, _08673_, _05477_);
  or (_08675_, _08674_, _05459_);
  nand (_08676_, _05455_, _07061_);
  or (_08677_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_08678_, _08677_, _08676_);
  and (_08679_, _08678_, _05473_);
  nand (_08680_, _05455_, _07341_);
  or (_08681_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_08683_, _08681_, _08680_);
  and (_08684_, _08683_, _05484_);
  nand (_08685_, _05455_, _06568_);
  or (_08686_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_08687_, _08686_, _08685_);
  and (_08688_, _08687_, _05497_);
  or (_08689_, _08688_, _08684_);
  or (_08690_, _08689_, _08679_);
  or (_08691_, _08690_, _08675_);
  nand (_08692_, _05455_, _07814_);
  or (_08693_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_08694_, _08693_, _08692_);
  and (_08695_, _08694_, _05477_);
  or (_08697_, _08695_, _05511_);
  nand (_08698_, _05455_, _08391_);
  or (_08699_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_08700_, _08699_, _08698_);
  and (_08702_, _08700_, _05484_);
  nand (_08703_, _05455_, _08110_);
  or (_08704_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_08706_, _08704_, _08703_);
  and (_08707_, _08706_, _05473_);
  or (_08708_, _08707_, _08702_);
  nand (_08709_, _05455_, _07601_);
  or (_08710_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_08711_, _08710_, _08709_);
  and (_08712_, _08711_, _05497_);
  or (_08713_, _08712_, _08708_);
  or (_08714_, _08713_, _08697_);
  and (_08715_, _08714_, _08691_);
  and (_08716_, _08715_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _08716_, _08670_);
  and (_08719_, _05537_, word_in[6]);
  nand (_08720_, _05455_, _06582_);
  or (_08722_, _05455_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_08724_, _08722_, _08720_);
  and (_08725_, _08724_, _05497_);
  or (_08727_, _08725_, _05459_);
  nand (_08728_, _05455_, _07074_);
  or (_08729_, _05455_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_08731_, _08729_, _08728_);
  and (_08732_, _08731_, _05473_);
  nand (_08734_, _05455_, _07361_);
  or (_08735_, _05455_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_08736_, _08735_, _08734_);
  and (_08737_, _08736_, _05484_);
  nand (_08738_, _05455_, _06817_);
  or (_08739_, _05455_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_08740_, _08739_, _08738_);
  and (_08742_, _08740_, _05477_);
  or (_08743_, _08742_, _08737_);
  or (_08744_, _08743_, _08732_);
  or (_08745_, _08744_, _08727_);
  nand (_08746_, _05455_, _07614_);
  or (_08747_, _05455_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_08748_, _08747_, _08746_);
  and (_08749_, _08748_, _05497_);
  or (_08750_, _08749_, _05511_);
  nand (_08751_, _05455_, _08121_);
  or (_08752_, _05455_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_08753_, _08752_, _08751_);
  and (_08754_, _08753_, _05473_);
  nand (_08755_, _05455_, _08406_);
  or (_08756_, _05455_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_08757_, _08756_, _08755_);
  and (_08758_, _08757_, _05484_);
  nand (_08760_, _05455_, _07829_);
  or (_08762_, _05455_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_08763_, _08762_, _08760_);
  and (_08764_, _08763_, _05477_);
  or (_08765_, _08764_, _08758_);
  or (_08766_, _08765_, _08754_);
  or (_08767_, _08766_, _08750_);
  and (_08768_, _08767_, _08745_);
  and (_08769_, _08768_, _05536_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _08769_, _08719_);
  and (_08770_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_08771_, _08427_, _23791_);
  or (_27049_, _08771_, _08770_);
  and (_08773_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_08774_, _08427_, _23982_);
  or (_27051_, _08774_, _08773_);
  and (_08775_, _05639_, word_in[8]);
  nand (_08776_, _05455_, _06616_);
  or (_08778_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_08779_, _08778_, _08776_);
  and (_08781_, _08779_, _05641_);
  nand (_08782_, _05455_, _06326_);
  or (_08783_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_08784_, _08783_, _08782_);
  and (_08785_, _08784_, _05640_);
  or (_08786_, _08785_, _08781_);
  and (_08788_, _08786_, _05606_);
  nand (_08789_, _05455_, _07643_);
  or (_08791_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_08792_, _08791_, _08789_);
  and (_08793_, _08792_, _05641_);
  nand (_08794_, _05455_, _07393_);
  or (_08795_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_08796_, _08795_, _08794_);
  and (_08797_, _08796_, _05640_);
  or (_08798_, _08797_, _08793_);
  and (_08799_, _08798_, _05608_);
  nand (_08801_, _05455_, _07113_);
  or (_08802_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_08803_, _08802_, _08801_);
  and (_08804_, _08803_, _05641_);
  nand (_08805_, _05455_, _06845_);
  or (_08807_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_08808_, _08807_, _08805_);
  and (_08809_, _08808_, _05640_);
  or (_08810_, _08809_, _08804_);
  and (_08811_, _08810_, _05670_);
  nand (_08813_, _05455_, _08182_);
  or (_08814_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_08816_, _08814_, _08813_);
  and (_08817_, _08816_, _05641_);
  nand (_08818_, _05455_, _07880_);
  or (_08820_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_08822_, _08820_, _08818_);
  and (_08823_, _08822_, _05640_);
  or (_08824_, _08823_, _08817_);
  and (_08825_, _08824_, _05684_);
  or (_08826_, _08825_, _08811_);
  or (_08827_, _08826_, _08799_);
  nor (_08828_, _08827_, _08788_);
  nor (_08830_, _08828_, _05639_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _08830_, _08775_);
  and (_08831_, _05639_, word_in[9]);
  nand (_08832_, _05455_, _06633_);
  or (_08833_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_08834_, _08833_, _08832_);
  and (_08835_, _08834_, _05641_);
  nand (_08836_, _05455_, _06344_);
  or (_08837_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_08838_, _08837_, _08836_);
  and (_08839_, _08838_, _05640_);
  or (_08840_, _08839_, _08835_);
  and (_08841_, _08840_, _05606_);
  nand (_08843_, _05455_, _07657_);
  or (_08845_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_08846_, _08845_, _08843_);
  and (_08847_, _08846_, _05641_);
  nand (_08848_, _05455_, _07419_);
  or (_08850_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_08851_, _08850_, _08848_);
  and (_08853_, _08851_, _05640_);
  or (_08854_, _08853_, _08847_);
  and (_08855_, _08854_, _05608_);
  nand (_08856_, _05455_, _07133_);
  or (_08857_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_08858_, _08857_, _08856_);
  and (_08859_, _08858_, _05641_);
  nand (_08860_, _05455_, _06865_);
  or (_08861_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_08862_, _08861_, _08860_);
  and (_08863_, _08862_, _05640_);
  or (_08864_, _08863_, _08859_);
  and (_08865_, _08864_, _05670_);
  nand (_08866_, _05455_, _08205_);
  or (_08867_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_08868_, _08867_, _08866_);
  and (_08869_, _08868_, _05641_);
  nand (_08870_, _05455_, _07911_);
  or (_08871_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_08872_, _08871_, _08870_);
  and (_08873_, _08872_, _05640_);
  or (_08874_, _08873_, _08869_);
  and (_08875_, _08874_, _05684_);
  or (_08876_, _08875_, _08865_);
  or (_08877_, _08876_, _08855_);
  nor (_08879_, _08877_, _08841_);
  nor (_08880_, _08879_, _05639_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _08880_, _08831_);
  and (_08881_, _05639_, word_in[10]);
  nand (_08882_, _05455_, _06647_);
  or (_08883_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_08885_, _08883_, _08882_);
  and (_08886_, _08885_, _05641_);
  nand (_08887_, _05455_, _06361_);
  or (_08889_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_08890_, _08889_, _08887_);
  and (_08891_, _08890_, _05640_);
  or (_08892_, _08891_, _08886_);
  and (_08893_, _08892_, _05606_);
  nand (_08894_, _05455_, _07668_);
  or (_08895_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_08896_, _08895_, _08894_);
  and (_08897_, _08896_, _05641_);
  nand (_08898_, _05455_, _07436_);
  or (_08899_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_08900_, _08899_, _08898_);
  and (_08901_, _08900_, _05640_);
  or (_08902_, _08901_, _08897_);
  and (_08903_, _08902_, _05608_);
  nand (_08905_, _05455_, _07146_);
  or (_08906_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_08908_, _08906_, _08905_);
  and (_08909_, _08908_, _05641_);
  nand (_08910_, _05455_, _06876_);
  or (_08911_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_08912_, _08911_, _08910_);
  and (_08913_, _08912_, _05640_);
  or (_08915_, _08913_, _08909_);
  and (_08916_, _08915_, _05670_);
  nand (_08918_, _05455_, _08217_);
  or (_08919_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_08920_, _08919_, _08918_);
  and (_08922_, _08920_, _05641_);
  nand (_08924_, _05455_, _07931_);
  or (_08925_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_08926_, _08925_, _08924_);
  and (_08928_, _08926_, _05640_);
  or (_08929_, _08928_, _08922_);
  and (_08930_, _08929_, _05684_);
  or (_08931_, _08930_, _08916_);
  or (_08932_, _08931_, _08903_);
  nor (_08933_, _08932_, _08893_);
  nor (_08934_, _08933_, _05639_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _08934_, _08881_);
  and (_08936_, _05639_, word_in[11]);
  nand (_08938_, _05455_, _06661_);
  or (_08940_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_08942_, _08940_, _08938_);
  and (_08943_, _08942_, _05641_);
  nand (_08944_, _05455_, _06383_);
  or (_08945_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_08946_, _08945_, _08944_);
  and (_08947_, _08946_, _05640_);
  or (_08948_, _08947_, _08943_);
  and (_08949_, _08948_, _05606_);
  nand (_08950_, _05455_, _07680_);
  or (_08952_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_08953_, _08952_, _08950_);
  and (_08955_, _08953_, _05641_);
  nand (_08957_, _05455_, _07455_);
  or (_08958_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_08960_, _08958_, _08957_);
  and (_08962_, _08960_, _05640_);
  or (_08963_, _08962_, _08955_);
  and (_08964_, _08963_, _05608_);
  nand (_08966_, _05455_, _07160_);
  or (_08967_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_08969_, _08967_, _08966_);
  and (_08970_, _08969_, _05641_);
  nand (_08971_, _05455_, _06889_);
  or (_08974_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_08975_, _08974_, _08971_);
  and (_08977_, _08975_, _05640_);
  or (_08978_, _08977_, _08970_);
  and (_08979_, _08978_, _05670_);
  nand (_08980_, _05455_, _08232_);
  or (_08981_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_08982_, _08981_, _08980_);
  and (_08983_, _08982_, _05641_);
  nand (_08984_, _05455_, _07948_);
  or (_08986_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_08987_, _08986_, _08984_);
  and (_08988_, _08987_, _05640_);
  or (_08990_, _08988_, _08983_);
  and (_08991_, _08990_, _05684_);
  or (_08992_, _08991_, _08979_);
  or (_08993_, _08992_, _08964_);
  nor (_08994_, _08993_, _08949_);
  nor (_08995_, _08994_, _05639_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _08995_, _08936_);
  and (_08997_, _05639_, word_in[12]);
  nand (_08998_, _05455_, _06672_);
  or (_08999_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_09000_, _08999_, _08998_);
  and (_09001_, _09000_, _05641_);
  nand (_09002_, _05455_, _06399_);
  or (_09003_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_09004_, _09003_, _09002_);
  and (_09005_, _09004_, _05640_);
  or (_09006_, _09005_, _09001_);
  and (_09007_, _09006_, _05606_);
  nand (_09008_, _05455_, _07694_);
  or (_09009_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_09010_, _09009_, _09008_);
  and (_09011_, _09010_, _05641_);
  nand (_09012_, _05455_, _07473_);
  or (_09013_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_09014_, _09013_, _09012_);
  and (_09015_, _09014_, _05640_);
  or (_09016_, _09015_, _09011_);
  and (_09017_, _09016_, _05608_);
  nand (_09019_, _05455_, _07174_);
  or (_09020_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_09021_, _09020_, _09019_);
  and (_09022_, _09021_, _05641_);
  nand (_09023_, _05455_, _06910_);
  or (_09024_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_09025_, _09024_, _09023_);
  and (_09026_, _09025_, _05640_);
  or (_09028_, _09026_, _09022_);
  and (_09030_, _09028_, _05670_);
  nand (_09031_, _05455_, _08244_);
  or (_09032_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_09033_, _09032_, _09031_);
  and (_09034_, _09033_, _05641_);
  nand (_09035_, _05455_, _07964_);
  or (_09036_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_09037_, _09036_, _09035_);
  and (_09038_, _09037_, _05640_);
  or (_09039_, _09038_, _09034_);
  and (_09040_, _09039_, _05684_);
  or (_09041_, _09040_, _09030_);
  or (_09042_, _09041_, _09017_);
  nor (_09043_, _09042_, _09007_);
  nor (_09044_, _09043_, _05639_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _09044_, _08997_);
  and (_09045_, _05639_, word_in[13]);
  nand (_09046_, _05455_, _06685_);
  or (_09047_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_09048_, _09047_, _09046_);
  and (_09050_, _09048_, _05641_);
  nand (_09052_, _05455_, _06417_);
  or (_09054_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_09055_, _09054_, _09052_);
  and (_09057_, _09055_, _05640_);
  or (_09058_, _09057_, _09050_);
  and (_09059_, _09058_, _05606_);
  nand (_09060_, _05455_, _07705_);
  or (_09061_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_09063_, _09061_, _09060_);
  and (_09064_, _09063_, _05641_);
  nand (_09065_, _05455_, _07485_);
  or (_09066_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_09068_, _09066_, _09065_);
  and (_09070_, _09068_, _05640_);
  or (_09072_, _09070_, _09064_);
  and (_09073_, _09072_, _05608_);
  nand (_09074_, _05455_, _07192_);
  or (_09075_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_09077_, _09075_, _09074_);
  and (_09079_, _09077_, _05641_);
  nand (_09080_, _05455_, _06929_);
  or (_09081_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_09082_, _09081_, _09080_);
  and (_09084_, _09082_, _05640_);
  or (_09085_, _09084_, _09079_);
  and (_09086_, _09085_, _05670_);
  nand (_09087_, _05455_, _08257_);
  or (_09088_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_09089_, _09088_, _09087_);
  and (_09090_, _09089_, _05641_);
  nand (_09092_, _05455_, _07978_);
  or (_09093_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_09095_, _09093_, _09092_);
  and (_09096_, _09095_, _05640_);
  or (_09098_, _09096_, _09090_);
  and (_09099_, _09098_, _05684_);
  or (_09100_, _09099_, _09086_);
  or (_09102_, _09100_, _09073_);
  nor (_09103_, _09102_, _09059_);
  nor (_09105_, _09103_, _05639_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _09105_, _09045_);
  and (_09107_, _05639_, word_in[14]);
  nand (_09108_, _05455_, _06702_);
  or (_09110_, _05455_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_09111_, _09110_, _09108_);
  and (_09113_, _09111_, _05641_);
  nand (_09114_, _05455_, _06427_);
  or (_09116_, _05455_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_09117_, _09116_, _09114_);
  and (_09119_, _09117_, _05640_);
  or (_09120_, _09119_, _09113_);
  and (_09121_, _09120_, _05606_);
  nand (_09123_, _05455_, _07718_);
  or (_09124_, _05455_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_09125_, _09124_, _09123_);
  and (_09127_, _09125_, _05641_);
  nand (_09128_, _05455_, _07500_);
  or (_09129_, _05455_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_09131_, _09129_, _09128_);
  and (_09133_, _09131_, _05640_);
  or (_09134_, _09133_, _09127_);
  and (_09135_, _09134_, _05608_);
  nand (_09136_, _05455_, _07209_);
  or (_09138_, _05455_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_09139_, _09138_, _09136_);
  and (_09141_, _09139_, _05641_);
  nand (_09143_, _05455_, _06943_);
  or (_09144_, _05455_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_09145_, _09144_, _09143_);
  and (_09146_, _09145_, _05640_);
  or (_09147_, _09146_, _09141_);
  and (_09149_, _09147_, _05670_);
  nand (_09151_, _05455_, _08271_);
  or (_09153_, _05455_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_09154_, _09153_, _09151_);
  and (_09156_, _09154_, _05641_);
  nand (_09157_, _05455_, _07992_);
  or (_09158_, _05455_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_09160_, _09158_, _09157_);
  and (_09161_, _09160_, _05640_);
  or (_09162_, _09161_, _09156_);
  and (_09163_, _09162_, _05684_);
  or (_09164_, _09163_, _09149_);
  or (_09165_, _09164_, _09135_);
  nor (_09166_, _09165_, _09121_);
  nor (_09167_, _09166_, _05639_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _09167_, _09107_);
  and (_09168_, _24615_, _23854_);
  not (_09169_, _09168_);
  and (_09170_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_09171_, _09168_, _23718_);
  or (_02844_, _09171_, _09170_);
  and (_09172_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_09173_, _08427_, _23755_);
  or (_02846_, _09173_, _09172_);
  and (_09174_, _05750_, word_in[16]);
  and (_09175_, _08438_, _05484_);
  and (_09176_, _08447_, _05473_);
  or (_09177_, _09176_, _09175_);
  and (_09178_, _08443_, _05477_);
  and (_09179_, _08451_, _05497_);
  or (_09180_, _09179_, _09178_);
  or (_09181_, _09180_, _09177_);
  or (_09182_, _09181_, _05706_);
  and (_09183_, _08459_, _05484_);
  and (_09184_, _08469_, _05473_);
  or (_09185_, _09184_, _09183_);
  and (_09186_, _08465_, _05477_);
  and (_09187_, _08473_, _05497_);
  or (_09189_, _09187_, _09186_);
  nor (_09190_, _09189_, _09185_);
  nand (_09191_, _09190_, _05706_);
  nand (_09192_, _09191_, _09182_);
  nor (_09193_, _09192_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _09193_, _09174_);
  and (_09195_, _05750_, word_in[17]);
  and (_09196_, _08484_, _05484_);
  and (_09197_, _08493_, _05473_);
  or (_09199_, _09197_, _09196_);
  and (_09200_, _08489_, _05477_);
  and (_09201_, _08497_, _05497_);
  or (_09203_, _09201_, _09200_);
  or (_09204_, _09203_, _09199_);
  or (_09206_, _09204_, _05706_);
  and (_09207_, _08516_, _05477_);
  and (_09208_, _08505_, _05484_);
  or (_09209_, _09208_, _09207_);
  and (_09210_, _08512_, _05473_);
  and (_09211_, _08522_, _05497_);
  or (_09212_, _09211_, _09210_);
  nor (_09213_, _09212_, _09209_);
  nand (_09214_, _09213_, _05706_);
  nand (_09215_, _09214_, _09206_);
  nor (_09216_, _09215_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _09216_, _09195_);
  and (_09217_, _05750_, word_in[18]);
  and (_09218_, _08537_, _05477_);
  and (_09219_, _08532_, _05484_);
  or (_09220_, _09219_, _09218_);
  and (_09221_, _08542_, _05473_);
  and (_09222_, _08547_, _05497_);
  or (_09223_, _09222_, _09221_);
  or (_09224_, _09223_, _09220_);
  or (_09225_, _09224_, _05706_);
  and (_09226_, _08555_, _05484_);
  and (_09227_, _08560_, _05473_);
  or (_09228_, _09227_, _09226_);
  and (_09229_, _08565_, _05477_);
  and (_09230_, _08571_, _05497_);
  or (_09231_, _09230_, _09229_);
  nor (_09232_, _09231_, _09228_);
  nand (_09234_, _09232_, _05706_);
  nand (_09236_, _09234_, _09225_);
  nor (_09237_, _09236_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _09237_, _09217_);
  and (_09238_, _05750_, word_in[19]);
  and (_09239_, _08581_, _05484_);
  and (_09240_, _08590_, _05473_);
  or (_09241_, _09240_, _09239_);
  and (_09243_, _08586_, _05477_);
  and (_09244_, _08596_, _05497_);
  or (_09245_, _09244_, _09243_);
  or (_09246_, _09245_, _09241_);
  or (_09247_, _09246_, _05706_);
  and (_09248_, _08603_, _05484_);
  and (_09249_, _08614_, _05473_);
  or (_09250_, _09249_, _09248_);
  and (_09252_, _08610_, _05477_);
  and (_09253_, _08618_, _05497_);
  or (_09254_, _09253_, _09252_);
  nor (_09255_, _09254_, _09250_);
  nand (_09256_, _09255_, _05706_);
  nand (_09257_, _09256_, _09247_);
  nor (_09258_, _09257_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _09258_, _09238_);
  and (_09259_, _05750_, word_in[20]);
  and (_09260_, _08634_, _05477_);
  and (_09261_, _08642_, _05484_);
  or (_09262_, _09261_, _09260_);
  and (_09263_, _08638_, _05473_);
  and (_09264_, _08629_, _05497_);
  or (_09265_, _09264_, _09263_);
  or (_09266_, _09265_, _09262_);
  or (_09267_, _09266_, _05706_);
  and (_09268_, _08664_, _05484_);
  and (_09269_, _08654_, _05473_);
  or (_09270_, _09269_, _09268_);
  and (_09272_, _08659_, _05477_);
  and (_09273_, _08649_, _05497_);
  or (_09274_, _09273_, _09272_);
  nor (_09275_, _09274_, _09270_);
  nand (_09276_, _09275_, _05706_);
  nand (_09277_, _09276_, _09267_);
  nor (_09278_, _09277_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _09278_, _09259_);
  and (_09279_, _05750_, word_in[21]);
  and (_09280_, _08687_, _05484_);
  and (_09282_, _08683_, _05473_);
  or (_09284_, _09282_, _09280_);
  and (_09286_, _08678_, _05477_);
  and (_09287_, _08673_, _05497_);
  or (_09288_, _09287_, _09286_);
  or (_09289_, _09288_, _09284_);
  or (_09290_, _09289_, _05706_);
  and (_09291_, _08711_, _05484_);
  and (_09292_, _08700_, _05473_);
  or (_09293_, _09292_, _09291_);
  and (_09294_, _08706_, _05477_);
  and (_09295_, _08694_, _05497_);
  or (_09296_, _09295_, _09294_);
  nor (_09297_, _09296_, _09293_);
  nand (_09298_, _09297_, _05706_);
  nand (_09299_, _09298_, _09290_);
  nor (_09300_, _09299_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _09300_, _09279_);
  and (_09301_, _05750_, word_in[22]);
  and (_09302_, _08724_, _05484_);
  and (_09303_, _08736_, _05473_);
  or (_09304_, _09303_, _09302_);
  and (_09306_, _08731_, _05477_);
  and (_09307_, _08740_, _05497_);
  or (_09308_, _09307_, _09306_);
  or (_09309_, _09308_, _09304_);
  or (_09310_, _09309_, _05706_);
  and (_09311_, _08753_, _05477_);
  and (_09312_, _08748_, _05484_);
  or (_09313_, _09312_, _09311_);
  and (_09314_, _08757_, _05473_);
  and (_09315_, _08763_, _05497_);
  or (_09316_, _09315_, _09314_);
  nor (_09317_, _09316_, _09313_);
  nand (_09318_, _09317_, _05706_);
  nand (_09319_, _09318_, _09310_);
  nor (_09320_, _09319_, _05750_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _09320_, _09301_);
  and (_09321_, _05808_, word_in[24]);
  and (_09322_, _08784_, _05641_);
  and (_09323_, _08779_, _05640_);
  or (_09324_, _09323_, _09322_);
  and (_09326_, _09324_, _05787_);
  and (_09327_, _08796_, _05641_);
  and (_09328_, _08792_, _05640_);
  or (_09330_, _09328_, _09327_);
  and (_09331_, _09330_, _05782_);
  and (_09332_, _08808_, _05641_);
  and (_09333_, _08803_, _05640_);
  or (_09334_, _09333_, _09332_);
  and (_09335_, _09334_, _05819_);
  and (_09336_, _08822_, _05641_);
  and (_09337_, _08816_, _05640_);
  or (_09338_, _09337_, _09336_);
  and (_09339_, _09338_, _05827_);
  or (_09340_, _09339_, _09335_);
  or (_09342_, _09340_, _09331_);
  nor (_09343_, _09342_, _09326_);
  nor (_09344_, _09343_, _05808_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _09344_, _09321_);
  and (_09345_, _05808_, word_in[25]);
  and (_09346_, _08851_, _05641_);
  and (_09348_, _08846_, _05640_);
  or (_09349_, _09348_, _09346_);
  and (_09350_, _09349_, _05782_);
  and (_09351_, _08838_, _05641_);
  and (_09352_, _08834_, _05640_);
  or (_09353_, _09352_, _09351_);
  and (_09354_, _09353_, _05787_);
  and (_09355_, _08862_, _05641_);
  and (_09356_, _08858_, _05640_);
  or (_09357_, _09356_, _09355_);
  and (_09358_, _09357_, _05819_);
  and (_09359_, _08872_, _05641_);
  and (_09360_, _08868_, _05640_);
  or (_09361_, _09360_, _09359_);
  and (_09363_, _09361_, _05827_);
  or (_09364_, _09363_, _09358_);
  or (_09365_, _09364_, _09354_);
  nor (_09367_, _09365_, _09350_);
  nor (_09368_, _09367_, _05808_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _09368_, _09345_);
  and (_09370_, _05808_, word_in[26]);
  and (_09371_, _08890_, _05641_);
  and (_09372_, _08885_, _05640_);
  or (_09373_, _09372_, _09371_);
  and (_09374_, _09373_, _05787_);
  and (_09375_, _08900_, _05641_);
  and (_09376_, _08896_, _05640_);
  or (_09377_, _09376_, _09375_);
  and (_09378_, _09377_, _05782_);
  and (_09379_, _08912_, _05641_);
  and (_09380_, _08908_, _05640_);
  or (_09381_, _09380_, _09379_);
  and (_09382_, _09381_, _05819_);
  and (_09383_, _08926_, _05641_);
  and (_09384_, _08920_, _05640_);
  or (_09385_, _09384_, _09383_);
  and (_09386_, _09385_, _05827_);
  or (_09387_, _09386_, _09382_);
  or (_09388_, _09387_, _09378_);
  nor (_09389_, _09388_, _09374_);
  nor (_09391_, _09389_, _05808_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _09391_, _09370_);
  and (_09393_, _05808_, word_in[27]);
  and (_09394_, _08960_, _05641_);
  and (_09395_, _08953_, _05640_);
  or (_09396_, _09395_, _09394_);
  and (_09397_, _09396_, _05782_);
  and (_09398_, _08946_, _05641_);
  and (_09399_, _08942_, _05640_);
  or (_09400_, _09399_, _09398_);
  and (_09401_, _09400_, _05787_);
  and (_09402_, _08975_, _05641_);
  and (_09403_, _08969_, _05640_);
  or (_09404_, _09403_, _09402_);
  and (_09405_, _09404_, _05819_);
  and (_09407_, _08987_, _05641_);
  and (_09408_, _08982_, _05640_);
  or (_09409_, _09408_, _09407_);
  and (_09410_, _09409_, _05827_);
  or (_09411_, _09410_, _09405_);
  or (_09412_, _09411_, _09401_);
  nor (_09413_, _09412_, _09397_);
  nor (_09414_, _09413_, _05808_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _09414_, _09393_);
  and (_09415_, _05808_, word_in[28]);
  and (_09416_, _09004_, _05641_);
  and (_09417_, _09000_, _05640_);
  or (_09418_, _09417_, _09416_);
  and (_09419_, _09418_, _05787_);
  and (_09420_, _09014_, _05641_);
  and (_09422_, _09010_, _05640_);
  or (_09423_, _09422_, _09420_);
  and (_09424_, _09423_, _05782_);
  and (_09425_, _09025_, _05641_);
  and (_09426_, _09021_, _05640_);
  or (_09427_, _09426_, _09425_);
  and (_09428_, _09427_, _05819_);
  and (_09429_, _09037_, _05641_);
  and (_09430_, _09033_, _05640_);
  or (_09431_, _09430_, _09429_);
  and (_09432_, _09431_, _05827_);
  or (_09433_, _09432_, _09428_);
  or (_09434_, _09433_, _09424_);
  nor (_09435_, _09434_, _09419_);
  nor (_09436_, _09435_, _05808_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _09436_, _09415_);
  and (_09437_, _05808_, word_in[29]);
  and (_09438_, _09068_, _05641_);
  and (_09440_, _09063_, _05640_);
  or (_09441_, _09440_, _09438_);
  and (_09442_, _09441_, _05782_);
  and (_09443_, _09055_, _05641_);
  and (_09444_, _09048_, _05640_);
  or (_09445_, _09444_, _09443_);
  and (_09446_, _09445_, _05787_);
  and (_09447_, _09082_, _05641_);
  and (_09448_, _09077_, _05640_);
  or (_09449_, _09448_, _09447_);
  and (_09450_, _09449_, _05819_);
  and (_09451_, _09095_, _05641_);
  and (_09453_, _09089_, _05640_);
  or (_09454_, _09453_, _09451_);
  and (_09455_, _09454_, _05827_);
  or (_09456_, _09455_, _09450_);
  or (_09457_, _09456_, _09446_);
  nor (_09458_, _09457_, _09442_);
  nor (_09459_, _09458_, _05808_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _09459_, _09437_);
  and (_09460_, _05808_, word_in[30]);
  and (_09461_, _09131_, _05641_);
  and (_09462_, _09125_, _05640_);
  or (_09463_, _09462_, _09461_);
  and (_09464_, _09463_, _05782_);
  and (_09465_, _09117_, _05641_);
  and (_09466_, _09111_, _05640_);
  or (_09467_, _09466_, _09465_);
  and (_09468_, _09467_, _05787_);
  and (_09469_, _09145_, _05641_);
  and (_09470_, _09139_, _05640_);
  or (_09471_, _09470_, _09469_);
  and (_09472_, _09471_, _05819_);
  and (_09473_, _09160_, _05641_);
  and (_09474_, _09154_, _05640_);
  or (_09475_, _09474_, _09473_);
  and (_09476_, _09475_, _05827_);
  or (_09477_, _09476_, _09472_);
  or (_09478_, _09477_, _09468_);
  nor (_09479_, _09478_, _09464_);
  nor (_09480_, _09479_, _05808_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _09480_, _09460_);
  and (_09481_, _24558_, _23641_);
  not (_09482_, _09481_);
  and (_09483_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_09484_, _09481_, _23791_);
  or (_02907_, _09484_, _09483_);
  nand (_09485_, _02077_, _23832_);
  and (_09486_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_09487_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_09488_, _09487_, _09486_);
  or (_09489_, _09488_, _02077_);
  and (_09491_, _09489_, _04740_);
  and (_09492_, _09491_, _09485_);
  and (_09493_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_09494_, _09493_, _09492_);
  and (_02930_, _09494_, _22761_);
  and (_09495_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_09496_, _09481_, _23838_);
  or (_27053_, _09496_, _09495_);
  or (_09497_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_09498_, _02078_);
  or (_09499_, _09498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_09500_, _09499_, _09497_);
  or (_09501_, _09500_, _02073_);
  nand (_09502_, _02073_, _23669_);
  and (_09503_, _09502_, _22761_);
  and (_02944_, _09503_, _09501_);
  and (_09504_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_09505_, _09481_, _23635_);
  or (_02946_, _09505_, _09504_);
  and (_09506_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_09508_, _03657_, _23755_);
  or (_27108_, _09508_, _09506_);
  and (_09509_, _24615_, _24103_);
  not (_09510_, _09509_);
  and (_09511_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and (_09512_, _09509_, _23676_);
  or (_02949_, _09512_, _09511_);
  and (_09513_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_09514_, _09481_, _23589_);
  or (_02952_, _09514_, _09513_);
  and (_09515_, _24615_, _23962_);
  not (_09516_, _09515_);
  and (_09517_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and (_09518_, _09515_, _23635_);
  or (_02955_, _09518_, _09517_);
  and (_09519_, _24615_, _24078_);
  not (_09520_, _09519_);
  and (_09521_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_09522_, _09519_, _23755_);
  or (_02959_, _09522_, _09521_);
  and (_09523_, _24558_, _24117_);
  not (_09524_, _09523_);
  and (_09525_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and (_09526_, _09523_, _23676_);
  or (_02965_, _09526_, _09525_);
  and (_09527_, _05351_, _05350_);
  and (_09528_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_09530_, _05387_, _05386_);
  and (_09531_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_09532_, _09531_, _09528_);
  and (_09533_, _09532_, _09527_);
  and (_09534_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_09535_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_09536_, _09535_, _09534_);
  and (_09537_, _09536_, _05352_);
  or (_09538_, _09537_, _09533_);
  and (_09539_, _09538_, _05373_);
  not (_09540_, _05373_);
  and (_09541_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_09542_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_09543_, _09542_, _09541_);
  and (_09544_, _09543_, _09527_);
  and (_09545_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_09547_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_09548_, _09547_, _09545_);
  and (_09549_, _09548_, _05352_);
  or (_09550_, _09549_, _09544_);
  and (_09551_, _09550_, _09540_);
  or (_09552_, _09551_, _05379_);
  or (_09553_, _09552_, _09539_);
  or (_09554_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_09555_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_09556_, _09555_, _05352_);
  and (_09557_, _09556_, _09554_);
  or (_09558_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_09559_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_09560_, _09559_, _09527_);
  and (_09561_, _09560_, _09558_);
  or (_09563_, _09561_, _09557_);
  and (_09564_, _09563_, _05373_);
  not (_09566_, _05379_);
  or (_09567_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_09568_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_09569_, _09568_, _05352_);
  and (_09570_, _09569_, _09567_);
  or (_09571_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_09572_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_09573_, _09572_, _09527_);
  and (_09574_, _09573_, _09571_);
  or (_09575_, _09574_, _09570_);
  and (_09576_, _09575_, _09540_);
  or (_09577_, _09576_, _09566_);
  or (_09578_, _09577_, _09564_);
  and (_09579_, _09578_, _09553_);
  or (_09580_, _09579_, _05361_);
  not (_09581_, _05361_);
  and (_09582_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_09584_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_09585_, _09584_, _09582_);
  and (_09586_, _09585_, _09527_);
  and (_09587_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_09588_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_09589_, _09588_, _09587_);
  and (_09590_, _09589_, _05352_);
  or (_09591_, _09590_, _09586_);
  and (_09592_, _09591_, _05373_);
  and (_09593_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_09594_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_09595_, _09594_, _09593_);
  and (_09596_, _09595_, _09527_);
  and (_09597_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_09598_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_09599_, _09598_, _09597_);
  and (_09600_, _09599_, _05352_);
  or (_09601_, _09600_, _09596_);
  and (_09602_, _09601_, _09540_);
  or (_09603_, _09602_, _05379_);
  or (_09604_, _09603_, _09592_);
  or (_09605_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_09606_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_09608_, _09606_, _09605_);
  and (_09609_, _09608_, _09527_);
  or (_09610_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_09611_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_09612_, _09611_, _09610_);
  and (_09613_, _09612_, _05352_);
  or (_09614_, _09613_, _09609_);
  and (_09615_, _09614_, _05373_);
  or (_09617_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_09618_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_09619_, _09618_, _09617_);
  and (_09620_, _09619_, _09527_);
  or (_09621_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_09622_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_09623_, _09622_, _09621_);
  and (_09624_, _09623_, _05352_);
  or (_09625_, _09624_, _09620_);
  and (_09626_, _09625_, _09540_);
  or (_09627_, _09626_, _09566_);
  or (_09628_, _09627_, _09615_);
  and (_09629_, _09628_, _09604_);
  or (_09630_, _09629_, _09581_);
  and (_09631_, _09630_, _05363_);
  and (_09633_, _09631_, _09580_);
  and (_09634_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_09635_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_09636_, _09635_, _09634_);
  and (_09637_, _09636_, _09527_);
  and (_09638_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_09639_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_09640_, _09639_, _09638_);
  and (_09641_, _09640_, _05352_);
  or (_09642_, _09641_, _09637_);
  or (_09643_, _09642_, _09540_);
  and (_09644_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_09645_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_09646_, _09645_, _09644_);
  and (_09647_, _09646_, _09527_);
  and (_09648_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_09649_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_09651_, _09649_, _09648_);
  and (_09652_, _09651_, _05352_);
  or (_09653_, _09652_, _09647_);
  or (_09654_, _09653_, _05373_);
  and (_09655_, _09654_, _09566_);
  and (_09656_, _09655_, _09643_);
  or (_09657_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_09658_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_09659_, _09658_, _09657_);
  and (_09660_, _09659_, _09527_);
  or (_09661_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_09662_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_09663_, _09662_, _09661_);
  and (_09664_, _09663_, _05352_);
  or (_09665_, _09664_, _09660_);
  or (_09666_, _09665_, _09540_);
  or (_09667_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_09669_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_09670_, _09669_, _09667_);
  and (_09671_, _09670_, _09527_);
  or (_09672_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_09673_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_09674_, _09673_, _09672_);
  and (_09675_, _09674_, _05352_);
  or (_09676_, _09675_, _09671_);
  or (_09677_, _09676_, _05373_);
  and (_09678_, _09677_, _05379_);
  and (_09679_, _09678_, _09666_);
  or (_09680_, _09679_, _09656_);
  or (_09681_, _09680_, _09581_);
  not (_09682_, _05363_);
  and (_09683_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_09684_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_09685_, _09684_, _09683_);
  and (_09686_, _09685_, _09527_);
  and (_09687_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_09688_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_09689_, _09688_, _09687_);
  and (_09690_, _09689_, _05352_);
  or (_09691_, _09690_, _09686_);
  or (_09692_, _09691_, _09540_);
  and (_09693_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_09694_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_09695_, _09694_, _09693_);
  and (_09696_, _09695_, _09527_);
  and (_09697_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_09698_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_09699_, _09698_, _09697_);
  and (_09700_, _09699_, _05352_);
  or (_09702_, _09700_, _09696_);
  or (_09703_, _09702_, _05373_);
  and (_09704_, _09703_, _09566_);
  and (_09705_, _09704_, _09692_);
  or (_09707_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_09708_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_09709_, _09708_, _05352_);
  and (_09710_, _09709_, _09707_);
  or (_09711_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_09712_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_09713_, _09712_, _09527_);
  and (_09714_, _09713_, _09711_);
  or (_09715_, _09714_, _09710_);
  or (_09716_, _09715_, _09540_);
  or (_09717_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_09718_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_09720_, _09718_, _05352_);
  and (_09721_, _09720_, _09717_);
  or (_09722_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_09723_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_09724_, _09723_, _09527_);
  and (_09726_, _09724_, _09722_);
  or (_09727_, _09726_, _09721_);
  or (_09728_, _09727_, _05373_);
  and (_09730_, _09728_, _05379_);
  and (_09732_, _09730_, _09716_);
  or (_09733_, _09732_, _09705_);
  or (_09734_, _09733_, _05361_);
  and (_09735_, _09734_, _09682_);
  and (_09736_, _09735_, _09681_);
  or (_09737_, _09736_, _09633_);
  or (_09738_, _09737_, _05357_);
  not (_09739_, _05357_);
  and (_09741_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_09742_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_09743_, _09742_, _09741_);
  and (_09744_, _09743_, _09527_);
  and (_09745_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_09747_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_09748_, _09747_, _09745_);
  and (_09749_, _09748_, _05352_);
  or (_09751_, _09749_, _09744_);
  and (_09753_, _09751_, _09540_);
  and (_09755_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_09756_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_09757_, _09756_, _09755_);
  and (_09758_, _09757_, _09527_);
  and (_09759_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_09760_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_09761_, _09760_, _09759_);
  and (_09763_, _09761_, _05352_);
  or (_09764_, _09763_, _09758_);
  and (_09765_, _09764_, _05373_);
  or (_09766_, _09765_, _09753_);
  and (_09768_, _09766_, _09566_);
  or (_09769_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_09770_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_09771_, _09770_, _09769_);
  and (_09772_, _09771_, _09527_);
  or (_09773_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_09774_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_09777_, _09774_, _09773_);
  and (_09778_, _09777_, _05352_);
  or (_09779_, _09778_, _09772_);
  and (_09780_, _09779_, _09540_);
  or (_09782_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_09783_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_09784_, _09783_, _09782_);
  and (_09785_, _09784_, _09527_);
  or (_09786_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_09787_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_09789_, _09787_, _09786_);
  and (_09790_, _09789_, _05352_);
  or (_09792_, _09790_, _09785_);
  and (_09793_, _09792_, _05373_);
  or (_09794_, _09793_, _09780_);
  and (_09795_, _09794_, _05379_);
  or (_09796_, _09795_, _09768_);
  or (_09797_, _09796_, _09581_);
  and (_09799_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_09800_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_09801_, _09800_, _09799_);
  and (_09802_, _09801_, _09527_);
  and (_09803_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_09804_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_09805_, _09804_, _09803_);
  and (_09807_, _09805_, _05352_);
  or (_09808_, _09807_, _09802_);
  and (_09809_, _09808_, _09540_);
  and (_09810_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_09812_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_09813_, _09812_, _09810_);
  and (_09814_, _09813_, _09527_);
  and (_09815_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_09817_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_09819_, _09817_, _09815_);
  and (_09820_, _09819_, _05352_);
  or (_09822_, _09820_, _09814_);
  and (_09824_, _09822_, _05373_);
  or (_09825_, _09824_, _09809_);
  and (_09826_, _09825_, _09566_);
  or (_09828_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_09829_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_09830_, _09829_, _05352_);
  and (_09831_, _09830_, _09828_);
  or (_09832_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_09833_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_09834_, _09833_, _09527_);
  and (_09836_, _09834_, _09832_);
  or (_09837_, _09836_, _09831_);
  and (_09839_, _09837_, _09540_);
  or (_09840_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_09842_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_09843_, _09842_, _05352_);
  and (_09844_, _09843_, _09840_);
  or (_09845_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_09846_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_09848_, _09846_, _09527_);
  and (_09849_, _09848_, _09845_);
  or (_09850_, _09849_, _09844_);
  and (_09851_, _09850_, _05373_);
  or (_09853_, _09851_, _09839_);
  and (_09855_, _09853_, _05379_);
  or (_09856_, _09855_, _09826_);
  or (_09857_, _09856_, _05361_);
  and (_09858_, _09857_, _05363_);
  and (_09859_, _09858_, _09797_);
  and (_09860_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_09862_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_09863_, _09862_, _09860_);
  and (_09864_, _09863_, _09527_);
  and (_09865_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_09866_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_09867_, _09866_, _09865_);
  and (_09868_, _09867_, _05352_);
  or (_09869_, _09868_, _09864_);
  or (_09870_, _09869_, _09540_);
  and (_09871_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_09872_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_09873_, _09872_, _09871_);
  and (_09874_, _09873_, _09527_);
  and (_09876_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_09877_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_09878_, _09877_, _09876_);
  and (_09880_, _09878_, _05352_);
  or (_09881_, _09880_, _09874_);
  or (_09882_, _09881_, _05373_);
  and (_09883_, _09882_, _09566_);
  and (_09884_, _09883_, _09870_);
  or (_09885_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_09886_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_09887_, _09886_, _05352_);
  and (_09888_, _09887_, _09885_);
  or (_09890_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_09891_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_09893_, _09891_, _09527_);
  and (_09895_, _09893_, _09890_);
  or (_09896_, _09895_, _09888_);
  or (_09898_, _09896_, _09540_);
  or (_09899_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_09901_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_09903_, _09901_, _05352_);
  and (_09904_, _09903_, _09899_);
  or (_09905_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_09906_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_09908_, _09906_, _09527_);
  and (_09909_, _09908_, _09905_);
  or (_09910_, _09909_, _09904_);
  or (_09911_, _09910_, _05373_);
  and (_09913_, _09911_, _05379_);
  and (_09914_, _09913_, _09898_);
  or (_09915_, _09914_, _09884_);
  or (_09916_, _09915_, _05361_);
  and (_09917_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_09918_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_09919_, _09918_, _09917_);
  and (_09921_, _09919_, _09527_);
  and (_09923_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_09924_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_09926_, _09924_, _09923_);
  and (_09927_, _09926_, _05352_);
  or (_09929_, _09927_, _09921_);
  or (_09930_, _09929_, _09540_);
  and (_09931_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_09933_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_09934_, _09933_, _09931_);
  and (_09936_, _09934_, _09527_);
  and (_09938_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_09940_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_09942_, _09940_, _09938_);
  and (_09943_, _09942_, _05352_);
  or (_09944_, _09943_, _09936_);
  or (_09945_, _09944_, _05373_);
  and (_09946_, _09945_, _09566_);
  and (_09948_, _09946_, _09930_);
  or (_09949_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_09951_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_09952_, _09951_, _09949_);
  and (_09953_, _09952_, _09527_);
  or (_09954_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_09955_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_09957_, _09955_, _09954_);
  and (_09958_, _09957_, _05352_);
  or (_09960_, _09958_, _09953_);
  or (_09961_, _09960_, _09540_);
  or (_09962_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_09964_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_09965_, _09964_, _09962_);
  and (_09966_, _09965_, _09527_);
  or (_09967_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_09968_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_09970_, _09968_, _09967_);
  and (_09971_, _09970_, _05352_);
  or (_09972_, _09971_, _09966_);
  or (_09973_, _09972_, _05373_);
  and (_09974_, _09973_, _05379_);
  and (_09975_, _09974_, _09961_);
  or (_09976_, _09975_, _09948_);
  or (_09977_, _09976_, _09581_);
  and (_09979_, _09977_, _09682_);
  and (_09980_, _09979_, _09916_);
  or (_09982_, _09980_, _09859_);
  or (_09984_, _09982_, _09739_);
  and (_09985_, _09984_, _26838_);
  and (_09986_, _09985_, _09738_);
  and (_09987_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_09989_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_09990_, _09989_, _09987_);
  and (_09991_, _09990_, _09527_);
  and (_09992_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_09993_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_09996_, _09993_, _09992_);
  and (_09998_, _09996_, _05352_);
  or (_09999_, _09998_, _09991_);
  or (_10000_, _09999_, _09540_);
  and (_10002_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_10003_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_10004_, _10003_, _10002_);
  and (_10005_, _10004_, _09527_);
  and (_10006_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_10007_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_10009_, _10007_, _10006_);
  and (_10010_, _10009_, _05352_);
  or (_10011_, _10010_, _10005_);
  or (_10012_, _10011_, _05373_);
  and (_10013_, _10012_, _09566_);
  and (_10014_, _10013_, _10000_);
  or (_10015_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_10016_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_10017_, _10016_, _10015_);
  and (_10018_, _10017_, _09527_);
  or (_10020_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_10021_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_10022_, _10021_, _10020_);
  and (_10023_, _10022_, _05352_);
  or (_10024_, _10023_, _10018_);
  or (_10026_, _10024_, _09540_);
  or (_10027_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_10028_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_10029_, _10028_, _10027_);
  and (_10031_, _10029_, _09527_);
  or (_10032_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_10033_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_10035_, _10033_, _10032_);
  and (_10037_, _10035_, _05352_);
  or (_10039_, _10037_, _10031_);
  or (_10040_, _10039_, _05373_);
  and (_10041_, _10040_, _05379_);
  and (_10042_, _10041_, _10026_);
  or (_10043_, _10042_, _10014_);
  and (_10044_, _10043_, _05361_);
  and (_10045_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_10047_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_10048_, _10047_, _10045_);
  and (_10049_, _10048_, _09527_);
  and (_10050_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and (_10051_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_10052_, _10051_, _10050_);
  and (_10053_, _10052_, _05352_);
  or (_10054_, _10053_, _10049_);
  or (_10055_, _10054_, _09540_);
  and (_10056_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_10057_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_10058_, _10057_, _10056_);
  and (_10059_, _10058_, _09527_);
  and (_10060_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_10061_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_10062_, _10061_, _10060_);
  and (_10063_, _10062_, _05352_);
  or (_10064_, _10063_, _10059_);
  or (_10065_, _10064_, _05373_);
  and (_10067_, _10065_, _09566_);
  and (_10068_, _10067_, _10055_);
  or (_10069_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_10071_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and (_10072_, _10071_, _05352_);
  and (_10074_, _10072_, _10069_);
  or (_10075_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_10076_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_10077_, _10076_, _09527_);
  and (_10078_, _10077_, _10075_);
  or (_10079_, _10078_, _10074_);
  or (_10081_, _10079_, _09540_);
  or (_10082_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_10083_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and (_10084_, _10083_, _05352_);
  and (_10085_, _10084_, _10082_);
  or (_10086_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_10087_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_10088_, _10087_, _09527_);
  and (_10090_, _10088_, _10086_);
  or (_10091_, _10090_, _10085_);
  or (_10093_, _10091_, _05373_);
  and (_10094_, _10093_, _05379_);
  and (_10095_, _10094_, _10081_);
  or (_10096_, _10095_, _10068_);
  and (_10097_, _10096_, _09581_);
  or (_10098_, _10097_, _10044_);
  and (_10099_, _10098_, _09682_);
  and (_10100_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and (_10101_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_10102_, _10101_, _10100_);
  and (_10103_, _10102_, _09527_);
  and (_10104_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_10106_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_10107_, _10106_, _10104_);
  and (_10108_, _10107_, _05352_);
  or (_10109_, _10108_, _10103_);
  and (_10111_, _10109_, _05373_);
  and (_10112_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and (_10113_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_10114_, _10113_, _10112_);
  and (_10115_, _10114_, _09527_);
  and (_10116_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_10117_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_10118_, _10117_, _10116_);
  and (_10119_, _10118_, _05352_);
  or (_10121_, _10119_, _10115_);
  and (_10122_, _10121_, _09540_);
  or (_10123_, _10122_, _10111_);
  and (_10125_, _10123_, _09566_);
  or (_10126_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_10128_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_10129_, _10128_, _05352_);
  and (_10130_, _10129_, _10126_);
  or (_10131_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_10132_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and (_10133_, _10132_, _09527_);
  and (_10134_, _10133_, _10131_);
  or (_10135_, _10134_, _10130_);
  and (_10137_, _10135_, _05373_);
  or (_10139_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_10140_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and (_10142_, _10140_, _05352_);
  and (_10144_, _10142_, _10139_);
  or (_10146_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_10147_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and (_10148_, _10147_, _09527_);
  and (_10149_, _10148_, _10146_);
  or (_10151_, _10149_, _10144_);
  and (_10152_, _10151_, _09540_);
  or (_10153_, _10152_, _10137_);
  and (_10154_, _10153_, _05379_);
  or (_10156_, _10154_, _10125_);
  and (_10157_, _10156_, _09581_);
  and (_10159_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_10161_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_10163_, _10161_, _10159_);
  and (_10164_, _10163_, _09527_);
  and (_10165_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_10166_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_10169_, _10166_, _10165_);
  and (_10170_, _10169_, _05352_);
  or (_10171_, _10170_, _10164_);
  and (_10173_, _10171_, _05373_);
  and (_10174_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and (_10176_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_10178_, _10176_, _10174_);
  and (_10179_, _10178_, _09527_);
  and (_10180_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_10181_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_10182_, _10181_, _10180_);
  and (_10183_, _10182_, _05352_);
  or (_10184_, _10183_, _10179_);
  and (_10186_, _10184_, _09540_);
  or (_10187_, _10186_, _10173_);
  and (_10188_, _10187_, _09566_);
  or (_10189_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_10190_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_10191_, _10190_, _10189_);
  and (_10192_, _10191_, _09527_);
  or (_10194_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_10195_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_10196_, _10195_, _10194_);
  and (_10197_, _10196_, _05352_);
  or (_10198_, _10197_, _10192_);
  and (_10199_, _10198_, _05373_);
  or (_10200_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_10201_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_10202_, _10201_, _10200_);
  and (_10204_, _10202_, _09527_);
  or (_10205_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_10206_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and (_10207_, _10206_, _10205_);
  and (_10208_, _10207_, _05352_);
  or (_10210_, _10208_, _10204_);
  and (_10211_, _10210_, _09540_);
  or (_10212_, _10211_, _10199_);
  and (_10214_, _10212_, _05379_);
  or (_10215_, _10214_, _10188_);
  and (_10217_, _10215_, _05361_);
  or (_10218_, _10217_, _10157_);
  and (_10220_, _10218_, _05363_);
  or (_10221_, _10220_, _10099_);
  or (_10222_, _10221_, _09739_);
  and (_10224_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_10225_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_10227_, _10225_, _10224_);
  and (_10228_, _10227_, _05352_);
  and (_10229_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_10230_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_10232_, _10230_, _10229_);
  and (_10234_, _10232_, _09527_);
  or (_10235_, _10234_, _10228_);
  or (_10236_, _10235_, _09540_);
  and (_10237_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_10238_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_10239_, _10238_, _10237_);
  and (_10240_, _10239_, _05352_);
  and (_10241_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and (_10242_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_10244_, _10242_, _10241_);
  and (_10245_, _10244_, _09527_);
  or (_10246_, _10245_, _10240_);
  or (_10247_, _10246_, _05373_);
  and (_10248_, _10247_, _09566_);
  and (_10249_, _10248_, _10236_);
  or (_10250_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_10251_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_10252_, _10251_, _09527_);
  and (_10253_, _10252_, _10250_);
  or (_10255_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_10256_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_10257_, _10256_, _05352_);
  and (_10258_, _10257_, _10255_);
  or (_10259_, _10258_, _10253_);
  or (_10260_, _10259_, _09540_);
  or (_10261_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_10262_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_10264_, _10262_, _09527_);
  and (_10265_, _10264_, _10261_);
  or (_10266_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_10267_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and (_10269_, _10267_, _05352_);
  and (_10270_, _10269_, _10266_);
  or (_10271_, _10270_, _10265_);
  or (_10272_, _10271_, _05373_);
  and (_10273_, _10272_, _05379_);
  and (_10274_, _10273_, _10260_);
  or (_10275_, _10274_, _10249_);
  and (_10276_, _10275_, _09581_);
  and (_10277_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_10278_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_10279_, _10278_, _09527_);
  or (_10280_, _10279_, _10277_);
  and (_10281_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_10282_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_10283_, _10282_, _05352_);
  or (_10284_, _10283_, _10281_);
  and (_10285_, _10284_, _10280_);
  or (_10286_, _10285_, _09540_);
  and (_10288_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and (_10289_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_10290_, _10289_, _09527_);
  or (_10291_, _10290_, _10288_);
  and (_10292_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_10293_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_10294_, _10293_, _05352_);
  or (_10295_, _10294_, _10292_);
  and (_10296_, _10295_, _10291_);
  or (_10297_, _10296_, _05373_);
  and (_10298_, _10297_, _09566_);
  and (_10299_, _10298_, _10286_);
  or (_10300_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_10301_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and (_10303_, _10301_, _10300_);
  or (_10304_, _10303_, _05352_);
  or (_10305_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_10306_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_10308_, _10306_, _10305_);
  or (_10309_, _10308_, _09527_);
  and (_10310_, _10309_, _10304_);
  or (_10311_, _10310_, _09540_);
  or (_10312_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_10313_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_10314_, _10313_, _10312_);
  or (_10315_, _10314_, _05352_);
  or (_10316_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_10317_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_10318_, _10317_, _10316_);
  or (_10319_, _10318_, _09527_);
  and (_10320_, _10319_, _10315_);
  or (_10321_, _10320_, _05373_);
  and (_10322_, _10321_, _05379_);
  and (_10323_, _10322_, _10311_);
  or (_10324_, _10323_, _10299_);
  and (_10325_, _10324_, _05361_);
  or (_10326_, _10325_, _10276_);
  and (_10327_, _10326_, _09682_);
  and (_10329_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_10330_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_10333_, _10330_, _10329_);
  and (_10334_, _10333_, _09527_);
  and (_10335_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_10336_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_10337_, _10336_, _10335_);
  and (_10338_, _10337_, _05352_);
  or (_10339_, _10338_, _10334_);
  and (_10340_, _10339_, _05373_);
  and (_10341_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_10342_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_10343_, _10342_, _10341_);
  and (_10344_, _10343_, _09527_);
  and (_10345_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and (_10346_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_10347_, _10346_, _10345_);
  and (_10349_, _10347_, _05352_);
  or (_10350_, _10349_, _10344_);
  and (_10351_, _10350_, _09540_);
  or (_10352_, _10351_, _10340_);
  and (_10353_, _10352_, _09566_);
  or (_10356_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_10357_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and (_10358_, _10357_, _10356_);
  and (_10359_, _10358_, _09527_);
  or (_10360_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_10361_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_10362_, _10361_, _10360_);
  and (_10363_, _10362_, _05352_);
  or (_10364_, _10363_, _10359_);
  and (_10365_, _10364_, _05373_);
  or (_10366_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_10367_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_10369_, _10367_, _10366_);
  and (_10370_, _10369_, _09527_);
  or (_10371_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_10372_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_10373_, _10372_, _10371_);
  and (_10375_, _10373_, _05352_);
  or (_10376_, _10375_, _10370_);
  and (_10377_, _10376_, _09540_);
  or (_10379_, _10377_, _10365_);
  and (_10381_, _10379_, _05379_);
  or (_10382_, _10381_, _10353_);
  and (_10383_, _10382_, _05361_);
  and (_10384_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_10385_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_10386_, _10385_, _10384_);
  and (_10387_, _10386_, _09527_);
  and (_10388_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_10389_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_10390_, _10389_, _10388_);
  and (_10392_, _10390_, _05352_);
  or (_10393_, _10392_, _10387_);
  and (_10394_, _10393_, _05373_);
  and (_10395_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_10396_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_10397_, _10396_, _10395_);
  and (_10398_, _10397_, _09527_);
  and (_10399_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_10400_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_10402_, _10400_, _10399_);
  and (_10403_, _10402_, _05352_);
  or (_10404_, _10403_, _10398_);
  and (_10405_, _10404_, _09540_);
  or (_10406_, _10405_, _10394_);
  and (_10407_, _10406_, _09566_);
  or (_10408_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_10409_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_10410_, _10409_, _10408_);
  and (_10411_, _10410_, _09527_);
  or (_10412_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_10413_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_10415_, _10413_, _10412_);
  and (_10416_, _10415_, _05352_);
  or (_10417_, _10416_, _10411_);
  and (_10419_, _10417_, _05373_);
  or (_10420_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_10421_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_10422_, _10421_, _10420_);
  and (_10423_, _10422_, _09527_);
  or (_10425_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_10426_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_10427_, _10426_, _10425_);
  and (_10428_, _10427_, _05352_);
  or (_10429_, _10428_, _10423_);
  and (_10430_, _10429_, _09540_);
  or (_10431_, _10430_, _10419_);
  and (_10432_, _10431_, _05379_);
  or (_10433_, _10432_, _10407_);
  and (_10434_, _10433_, _09581_);
  or (_10435_, _10434_, _10383_);
  and (_10436_, _10435_, _05363_);
  or (_10438_, _10436_, _10327_);
  or (_10439_, _10438_, _05357_);
  and (_10440_, _10439_, _04360_);
  and (_10441_, _10440_, _10222_);
  or (_10443_, _10441_, _09986_);
  or (_10444_, _10443_, _05401_);
  not (_10445_, _05401_);
  or (_10446_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_10448_, _10446_, _22761_);
  and (_02967_, _10448_, _10444_);
  or (_10449_, _25674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_10450_, _25674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_10452_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_10454_, _10452_, _25701_);
  nand (_10455_, _10454_, _10450_);
  and (_10456_, _10455_, _10449_);
  or (_10457_, _10456_, _25699_);
  nor (_10458_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_10459_, _10458_, _25667_);
  and (_10461_, _10459_, _10457_);
  and (_10462_, _25667_, _24763_);
  or (_10463_, _10462_, _25711_);
  or (_10464_, _10463_, _10461_);
  or (_10465_, _25716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_10466_, _10465_, _22761_);
  and (_02973_, _10466_, _10464_);
  and (_10467_, _25667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  not (_10468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_10470_, _25688_, _25674_);
  and (_10471_, _10470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_10472_, _10471_, _10468_);
  and (_10473_, _10471_, _10468_);
  or (_10474_, _10473_, _10472_);
  and (_10475_, _25703_, _25674_);
  and (_10476_, _10475_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_10477_, _10476_, _25701_);
  or (_10478_, _10477_, _25699_);
  or (_10479_, _10478_, _10474_);
  or (_10480_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_10481_, _10480_, _25712_);
  and (_10482_, _10481_, _10479_);
  or (_10483_, _10482_, _10467_);
  nor (_10484_, _25716_, _23628_);
  or (_10485_, _10484_, _10483_);
  and (_02992_, _10485_, _22761_);
  and (_10486_, _02436_, _23791_);
  and (_10487_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or (_02995_, _10487_, _10486_);
  and (_10488_, _02444_, _23838_);
  and (_10489_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_02997_, _10489_, _10488_);
  and (_10491_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  and (_10492_, _09523_, _23838_);
  or (_02999_, _10492_, _10491_);
  and (_10493_, _25696_, _06207_);
  or (_10494_, _10493_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_10495_, _10494_, _06195_);
  nand (_10496_, _03809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_10497_, _10496_, _06195_);
  or (_10498_, _10497_, _03810_);
  and (_10499_, _10498_, _10495_);
  or (_10501_, _10499_, _06202_);
  nand (_10502_, _06202_, _23748_);
  and (_10503_, _10502_, _22761_);
  and (_03002_, _10503_, _10501_);
  and (_10505_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and (_10506_, _09523_, _23982_);
  or (_27057_, _10506_, _10505_);
  and (_26869_[1], _24262_, _22761_);
  and (_10508_, _24567_, _23635_);
  and (_10509_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or (_03011_, _10509_, _10508_);
  and (_10510_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and (_10512_, _09523_, _23755_);
  or (_03020_, _10512_, _10510_);
  and (_10513_, _04692_, _23791_);
  and (_10514_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_03022_, _10514_, _10513_);
  and (_10515_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and (_10516_, _03657_, _23635_);
  or (_03026_, _10516_, _10515_);
  and (_10517_, _24558_, _24541_);
  not (_10518_, _10517_);
  and (_10519_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_10520_, _10517_, _23718_);
  or (_03036_, _10520_, _10519_);
  and (_10521_, _24214_, _23838_);
  and (_10522_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or (_03045_, _10522_, _10521_);
  and (_10524_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and (_10525_, _25294_, _23589_);
  or (_03049_, _10525_, _10524_);
  and (_10526_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_10527_, _10517_, _23838_);
  or (_27058_, _10527_, _10526_);
  and (_10529_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_10530_, _10517_, _23635_);
  or (_03060_, _10530_, _10529_);
  and (_10531_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and (_10532_, _25464_, _23791_);
  or (_27069_, _10532_, _10531_);
  and (_10533_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_10534_, _10517_, _23755_);
  or (_03071_, _10534_, _10533_);
  nand (_10535_, _22762_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_26914_, _10535_, _22761_);
  nand (_10537_, _26832_, _22761_);
  nor (_26918_, _10537_, _26676_);
  and (_10538_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and (_10539_, _04734_, _23755_);
  or (_03108_, _10539_, _10538_);
  and (_10540_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  and (_10541_, _04734_, _23635_);
  or (_03123_, _10541_, _10540_);
  and (_10542_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  and (_10543_, _02762_, _23982_);
  or (_03129_, _10543_, _10542_);
  and (_10544_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  and (_10545_, _04734_, _23982_);
  or (_03131_, _10545_, _10544_);
  or (_10547_, _01888_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_26911_[3], _10547_, _22761_);
  and (_10548_, _23864_, _23718_);
  and (_10549_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_03146_, _10549_, _10548_);
  and (_10550_, _03134_, _23838_);
  and (_10551_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or (_03153_, _10551_, _10550_);
  and (_10552_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  and (_10553_, _04599_, _23791_);
  or (_27121_, _10553_, _10552_);
  and (_10555_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_10556_, _06040_, _23982_);
  or (_03164_, _10556_, _10555_);
  and (_10557_, _04733_, _23854_);
  not (_10558_, _10557_);
  and (_10559_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  and (_10560_, _10557_, _23755_);
  or (_03172_, _10560_, _10559_);
  and (_10562_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_10563_, _02858_, _23718_);
  or (_03182_, _10563_, _10562_);
  and (_10564_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_10565_, _24616_, _23982_);
  or (_03186_, _10565_, _10564_);
  and (_10566_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_10568_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_10570_, _10568_, _10566_);
  and (_10571_, _10570_, _09527_);
  and (_10572_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_10573_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_10574_, _10573_, _10572_);
  and (_10575_, _10574_, _05352_);
  or (_10577_, _10575_, _10571_);
  and (_10578_, _10577_, _05373_);
  and (_10580_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_10581_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_10582_, _10581_, _10580_);
  and (_10583_, _10582_, _09527_);
  and (_10584_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_10585_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_10587_, _10585_, _10584_);
  and (_10588_, _10587_, _05352_);
  or (_10589_, _10588_, _10583_);
  and (_10590_, _10589_, _09540_);
  or (_10591_, _10590_, _05379_);
  or (_10593_, _10591_, _10578_);
  or (_10594_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_10595_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_10596_, _10595_, _05352_);
  and (_10597_, _10596_, _10594_);
  or (_10598_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_10599_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_10600_, _10599_, _09527_);
  and (_10601_, _10600_, _10598_);
  or (_10602_, _10601_, _10597_);
  and (_10603_, _10602_, _05373_);
  or (_10604_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_10605_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_10606_, _10605_, _05352_);
  and (_10608_, _10606_, _10604_);
  or (_10610_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_10612_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_10613_, _10612_, _09527_);
  and (_10614_, _10613_, _10610_);
  or (_10615_, _10614_, _10608_);
  and (_10617_, _10615_, _09540_);
  or (_10618_, _10617_, _09566_);
  or (_10619_, _10618_, _10603_);
  and (_10620_, _10619_, _10593_);
  or (_10621_, _10620_, _05361_);
  and (_10623_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_10624_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_10625_, _10624_, _10623_);
  and (_10626_, _10625_, _09527_);
  and (_10627_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_10629_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_10631_, _10629_, _10627_);
  and (_10632_, _10631_, _05352_);
  or (_10633_, _10632_, _10626_);
  and (_10634_, _10633_, _05373_);
  and (_10635_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_10636_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_10637_, _10636_, _10635_);
  and (_10638_, _10637_, _09527_);
  and (_10640_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_10641_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_10642_, _10641_, _10640_);
  and (_10643_, _10642_, _05352_);
  or (_10644_, _10643_, _10638_);
  and (_10645_, _10644_, _09540_);
  or (_10646_, _10645_, _05379_);
  or (_10647_, _10646_, _10634_);
  or (_10648_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_10649_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_10651_, _10649_, _10648_);
  and (_10652_, _10651_, _09527_);
  or (_10654_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_10655_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_10657_, _10655_, _10654_);
  and (_10658_, _10657_, _05352_);
  or (_10659_, _10658_, _10652_);
  and (_10660_, _10659_, _05373_);
  or (_10661_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_10662_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_10663_, _10662_, _10661_);
  and (_10664_, _10663_, _09527_);
  or (_10665_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_10666_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_10667_, _10666_, _10665_);
  and (_10668_, _10667_, _05352_);
  or (_10670_, _10668_, _10664_);
  and (_10671_, _10670_, _09540_);
  or (_10672_, _10671_, _09566_);
  or (_10674_, _10672_, _10660_);
  and (_10675_, _10674_, _10647_);
  or (_10677_, _10675_, _09581_);
  and (_10678_, _10677_, _05363_);
  and (_10680_, _10678_, _10621_);
  and (_10681_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_10682_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_10683_, _10682_, _10681_);
  and (_10684_, _10683_, _09527_);
  and (_10685_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_10686_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_10687_, _10686_, _10685_);
  and (_10689_, _10687_, _05352_);
  or (_10690_, _10689_, _10684_);
  or (_10691_, _10690_, _09540_);
  and (_10692_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_10693_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_10694_, _10693_, _10692_);
  and (_10695_, _10694_, _09527_);
  and (_10696_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_10697_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_10698_, _10697_, _10696_);
  and (_10699_, _10698_, _05352_);
  or (_10700_, _10699_, _10695_);
  or (_10701_, _10700_, _05373_);
  and (_10702_, _10701_, _09566_);
  and (_10703_, _10702_, _10691_);
  or (_10704_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_10705_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_10706_, _10705_, _10704_);
  and (_10707_, _10706_, _09527_);
  or (_10708_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_10709_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_10711_, _10709_, _10708_);
  and (_10712_, _10711_, _05352_);
  or (_10714_, _10712_, _10707_);
  or (_10715_, _10714_, _09540_);
  or (_10717_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_10719_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_10720_, _10719_, _10717_);
  and (_10722_, _10720_, _09527_);
  or (_10723_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_10725_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_10726_, _10725_, _10723_);
  and (_10728_, _10726_, _05352_);
  or (_10730_, _10728_, _10722_);
  or (_10731_, _10730_, _05373_);
  and (_10732_, _10731_, _05379_);
  and (_10733_, _10732_, _10715_);
  or (_10734_, _10733_, _10703_);
  or (_10735_, _10734_, _09581_);
  and (_10736_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_10738_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_10739_, _10738_, _10736_);
  and (_10740_, _10739_, _09527_);
  and (_10741_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_10743_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_10744_, _10743_, _10741_);
  and (_10746_, _10744_, _05352_);
  or (_10747_, _10746_, _10740_);
  or (_10748_, _10747_, _09540_);
  and (_10749_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_10750_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_10752_, _10750_, _10749_);
  and (_10753_, _10752_, _09527_);
  and (_10755_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_10757_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_10759_, _10757_, _10755_);
  and (_10760_, _10759_, _05352_);
  or (_10761_, _10760_, _10753_);
  or (_10763_, _10761_, _05373_);
  and (_10764_, _10763_, _09566_);
  and (_10765_, _10764_, _10748_);
  or (_10766_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_10767_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_10768_, _10767_, _05352_);
  and (_10769_, _10768_, _10766_);
  or (_10770_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_10771_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_10772_, _10771_, _09527_);
  and (_10773_, _10772_, _10770_);
  or (_10774_, _10773_, _10769_);
  or (_10775_, _10774_, _09540_);
  or (_10776_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_10778_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_10779_, _10778_, _05352_);
  and (_10781_, _10779_, _10776_);
  or (_10783_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_10784_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_10785_, _10784_, _09527_);
  and (_10786_, _10785_, _10783_);
  or (_10788_, _10786_, _10781_);
  or (_10789_, _10788_, _05373_);
  and (_10790_, _10789_, _05379_);
  and (_10791_, _10790_, _10775_);
  or (_10793_, _10791_, _10765_);
  or (_10794_, _10793_, _05361_);
  and (_10795_, _10794_, _09682_);
  and (_10796_, _10795_, _10735_);
  or (_10797_, _10796_, _10680_);
  or (_10798_, _10797_, _05357_);
  and (_10799_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_10800_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_10801_, _10800_, _10799_);
  and (_10803_, _10801_, _09527_);
  and (_10804_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_10805_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_10806_, _10805_, _10804_);
  and (_10808_, _10806_, _05352_);
  or (_10810_, _10808_, _10803_);
  and (_10812_, _10810_, _09540_);
  and (_10814_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_10816_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_10817_, _10816_, _10814_);
  and (_10819_, _10817_, _09527_);
  and (_10820_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_10821_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_10822_, _10821_, _10820_);
  and (_10824_, _10822_, _05352_);
  or (_10825_, _10824_, _10819_);
  and (_10826_, _10825_, _05373_);
  or (_10827_, _10826_, _10812_);
  and (_10829_, _10827_, _09566_);
  or (_10831_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_10833_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_10834_, _10833_, _10831_);
  and (_10836_, _10834_, _09527_);
  or (_10837_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_10839_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_10841_, _10839_, _10837_);
  and (_10842_, _10841_, _05352_);
  or (_10844_, _10842_, _10836_);
  and (_10846_, _10844_, _09540_);
  or (_10847_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_10848_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_10850_, _10848_, _10847_);
  and (_10851_, _10850_, _09527_);
  or (_10852_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_10853_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_10854_, _10853_, _10852_);
  and (_10855_, _10854_, _05352_);
  or (_10856_, _10855_, _10851_);
  and (_10857_, _10856_, _05373_);
  or (_10858_, _10857_, _10846_);
  and (_10859_, _10858_, _05379_);
  or (_10860_, _10859_, _10829_);
  or (_10862_, _10860_, _09581_);
  and (_10863_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and (_10864_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_10865_, _10864_, _10863_);
  and (_10867_, _10865_, _09527_);
  and (_10868_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and (_10870_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_10871_, _10870_, _10868_);
  and (_10873_, _10871_, _05352_);
  or (_10875_, _10873_, _10867_);
  and (_10877_, _10875_, _09540_);
  and (_10879_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_10881_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_10883_, _10881_, _10879_);
  and (_10884_, _10883_, _09527_);
  and (_10885_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and (_10886_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_10887_, _10886_, _10885_);
  and (_10889_, _10887_, _05352_);
  or (_10891_, _10889_, _10884_);
  and (_10892_, _10891_, _05373_);
  or (_10893_, _10892_, _10877_);
  and (_10894_, _10893_, _09566_);
  or (_10896_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_10898_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and (_10900_, _10898_, _05352_);
  and (_10901_, _10900_, _10896_);
  or (_10903_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_10906_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and (_10907_, _10906_, _09527_);
  and (_10908_, _10907_, _10903_);
  or (_10909_, _10908_, _10901_);
  and (_10910_, _10909_, _09540_);
  or (_10911_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_10912_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_10913_, _10912_, _05352_);
  and (_10914_, _10913_, _10911_);
  or (_10915_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_10916_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and (_10917_, _10916_, _09527_);
  and (_10918_, _10917_, _10915_);
  or (_10919_, _10918_, _10914_);
  and (_10920_, _10919_, _05373_);
  or (_10921_, _10920_, _10910_);
  and (_10922_, _10921_, _05379_);
  or (_10923_, _10922_, _10894_);
  or (_10924_, _10923_, _05361_);
  and (_10925_, _10924_, _05363_);
  and (_10926_, _10925_, _10862_);
  and (_10927_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_10928_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_10930_, _10928_, _10927_);
  and (_10931_, _10930_, _09527_);
  and (_10932_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_10933_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_10934_, _10933_, _10932_);
  and (_10935_, _10934_, _05352_);
  or (_10936_, _10935_, _10931_);
  or (_10937_, _10936_, _09540_);
  and (_10938_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_10939_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_10940_, _10939_, _10938_);
  and (_10941_, _10940_, _09527_);
  and (_10942_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_10943_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_10944_, _10943_, _10942_);
  and (_10946_, _10944_, _05352_);
  or (_10947_, _10946_, _10941_);
  or (_10948_, _10947_, _05373_);
  and (_10949_, _10948_, _09566_);
  and (_10950_, _10949_, _10937_);
  or (_10951_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_10952_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_10953_, _10952_, _05352_);
  and (_10954_, _10953_, _10951_);
  or (_10955_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_10956_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_10957_, _10956_, _09527_);
  and (_10958_, _10957_, _10955_);
  or (_10959_, _10958_, _10954_);
  or (_10960_, _10959_, _09540_);
  or (_10961_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_10962_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_10964_, _10962_, _05352_);
  and (_10965_, _10964_, _10961_);
  or (_10966_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_10967_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_10968_, _10967_, _09527_);
  and (_10969_, _10968_, _10966_);
  or (_10970_, _10969_, _10965_);
  or (_10971_, _10970_, _05373_);
  and (_10972_, _10971_, _05379_);
  and (_10973_, _10972_, _10960_);
  or (_10974_, _10973_, _10950_);
  or (_10975_, _10974_, _05361_);
  and (_10976_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_10978_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_10979_, _10978_, _10976_);
  and (_10981_, _10979_, _09527_);
  and (_10982_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_10983_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_10984_, _10983_, _10982_);
  and (_10985_, _10984_, _05352_);
  or (_10986_, _10985_, _10981_);
  or (_10987_, _10986_, _09540_);
  and (_10988_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_10989_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_10990_, _10989_, _10988_);
  and (_10991_, _10990_, _09527_);
  and (_10992_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_10993_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_10994_, _10993_, _10992_);
  and (_10995_, _10994_, _05352_);
  or (_10996_, _10995_, _10991_);
  or (_10997_, _10996_, _05373_);
  and (_10998_, _10997_, _09566_);
  and (_10999_, _10998_, _10987_);
  or (_11000_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_11001_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_11002_, _11001_, _11000_);
  and (_11003_, _11002_, _09527_);
  or (_11004_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_11005_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_11006_, _11005_, _11004_);
  and (_11007_, _11006_, _05352_);
  or (_11008_, _11007_, _11003_);
  or (_11009_, _11008_, _09540_);
  or (_11010_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_11011_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_11012_, _11011_, _11010_);
  and (_11013_, _11012_, _09527_);
  or (_11014_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_11015_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_11016_, _11015_, _11014_);
  and (_11017_, _11016_, _05352_);
  or (_11018_, _11017_, _11013_);
  or (_11019_, _11018_, _05373_);
  and (_11020_, _11019_, _05379_);
  and (_11021_, _11020_, _11009_);
  or (_11022_, _11021_, _10999_);
  or (_11023_, _11022_, _09581_);
  and (_11024_, _11023_, _09682_);
  and (_11025_, _11024_, _10975_);
  or (_11026_, _11025_, _10926_);
  or (_11027_, _11026_, _09739_);
  and (_11028_, _11027_, _26838_);
  and (_11029_, _11028_, _10798_);
  and (_11030_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_11032_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_11033_, _11032_, _11030_);
  and (_11034_, _11033_, _05352_);
  and (_11036_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_11037_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_11038_, _11037_, _11036_);
  and (_11039_, _11038_, _09527_);
  or (_11040_, _11039_, _11034_);
  or (_11042_, _11040_, _09540_);
  and (_11044_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_11045_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_11046_, _11045_, _11044_);
  and (_11047_, _11046_, _05352_);
  and (_11049_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_11050_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_11052_, _11050_, _11049_);
  and (_11053_, _11052_, _09527_);
  or (_11054_, _11053_, _11047_);
  or (_11055_, _11054_, _05373_);
  and (_11056_, _11055_, _09566_);
  and (_11058_, _11056_, _11042_);
  or (_11059_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_11060_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_11062_, _11060_, _09527_);
  and (_11064_, _11062_, _11059_);
  or (_11066_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_11067_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and (_11069_, _11067_, _05352_);
  and (_11070_, _11069_, _11066_);
  or (_11071_, _11070_, _11064_);
  or (_11072_, _11071_, _09540_);
  or (_11073_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_11074_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_11075_, _11074_, _09527_);
  and (_11076_, _11075_, _11073_);
  or (_11077_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_11078_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_11080_, _11078_, _05352_);
  and (_11081_, _11080_, _11077_);
  or (_11082_, _11081_, _11076_);
  or (_11084_, _11082_, _05373_);
  and (_11086_, _11084_, _05379_);
  and (_11087_, _11086_, _11072_);
  or (_11088_, _11087_, _11058_);
  and (_11089_, _11088_, _09581_);
  and (_11091_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_11092_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_11093_, _11092_, _09527_);
  or (_11094_, _11093_, _11091_);
  and (_11095_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_11096_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_11098_, _11096_, _05352_);
  or (_11099_, _11098_, _11095_);
  and (_11101_, _11099_, _11094_);
  or (_11103_, _11101_, _09540_);
  and (_11105_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_11106_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_11107_, _11106_, _09527_);
  or (_11109_, _11107_, _11105_);
  and (_11110_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_11113_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_11115_, _11113_, _05352_);
  or (_11117_, _11115_, _11110_);
  and (_11118_, _11117_, _11109_);
  or (_11120_, _11118_, _05373_);
  and (_11121_, _11120_, _09566_);
  and (_11122_, _11121_, _11103_);
  or (_11124_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_11126_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_11127_, _11126_, _11124_);
  or (_11128_, _11127_, _05352_);
  or (_11130_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_11131_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_11133_, _11131_, _11130_);
  or (_11134_, _11133_, _09527_);
  and (_11135_, _11134_, _11128_);
  or (_11136_, _11135_, _09540_);
  or (_11138_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_11140_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_11142_, _11140_, _11138_);
  or (_11145_, _11142_, _05352_);
  or (_11146_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_11148_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_11150_, _11148_, _11146_);
  or (_11152_, _11150_, _09527_);
  and (_11153_, _11152_, _11145_);
  or (_11155_, _11153_, _05373_);
  and (_11156_, _11155_, _05379_);
  and (_11157_, _11156_, _11136_);
  or (_11158_, _11157_, _11122_);
  and (_11160_, _11158_, _05361_);
  or (_11162_, _11160_, _11089_);
  and (_11163_, _11162_, _09682_);
  or (_11164_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_11165_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_11166_, _11165_, _11164_);
  and (_11167_, _11166_, _09527_);
  or (_11169_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_11171_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_11172_, _11171_, _11169_);
  and (_11173_, _11172_, _05352_);
  or (_11174_, _11173_, _11167_);
  and (_11175_, _11174_, _09540_);
  or (_11176_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_11177_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_11178_, _11177_, _11176_);
  and (_11179_, _11178_, _09527_);
  or (_11181_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_11183_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_11184_, _11183_, _11181_);
  and (_11185_, _11184_, _05352_);
  or (_11186_, _11185_, _11179_);
  and (_11188_, _11186_, _05373_);
  or (_11189_, _11188_, _11175_);
  and (_11190_, _11189_, _05379_);
  and (_11191_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_11193_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_11194_, _11193_, _11191_);
  and (_11195_, _11194_, _09527_);
  and (_11197_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_11198_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_11199_, _11198_, _11197_);
  and (_11200_, _11199_, _05352_);
  or (_11202_, _11200_, _11195_);
  and (_11203_, _11202_, _09540_);
  and (_11204_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_11205_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_11207_, _11205_, _11204_);
  and (_11208_, _11207_, _09527_);
  and (_11209_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_11210_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_11211_, _11210_, _11209_);
  and (_11212_, _11211_, _05352_);
  or (_11214_, _11212_, _11208_);
  and (_11215_, _11214_, _05373_);
  or (_11216_, _11215_, _11203_);
  and (_11218_, _11216_, _09566_);
  or (_11219_, _11218_, _11190_);
  and (_11220_, _11219_, _05361_);
  or (_11221_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_11223_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  and (_11224_, _11223_, _11221_);
  and (_11225_, _11224_, _09527_);
  or (_11227_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_11228_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  and (_11229_, _11228_, _11227_);
  and (_11230_, _11229_, _05352_);
  or (_11231_, _11230_, _11225_);
  and (_11232_, _11231_, _09540_);
  or (_11233_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_11234_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and (_11236_, _11234_, _11233_);
  and (_11238_, _11236_, _09527_);
  or (_11239_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or (_11241_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  and (_11243_, _11241_, _11239_);
  and (_11244_, _11243_, _05352_);
  or (_11246_, _11244_, _11238_);
  and (_11248_, _11246_, _05373_);
  or (_11249_, _11248_, _11232_);
  and (_11250_, _11249_, _05379_);
  and (_11251_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and (_11252_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_11253_, _11252_, _11251_);
  and (_11254_, _11253_, _09527_);
  and (_11256_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and (_11258_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or (_11259_, _11258_, _11256_);
  and (_11260_, _11259_, _05352_);
  or (_11261_, _11260_, _11254_);
  and (_11262_, _11261_, _09540_);
  and (_11264_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  and (_11266_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_11267_, _11266_, _11264_);
  and (_11268_, _11267_, _09527_);
  and (_11269_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  and (_11270_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or (_11271_, _11270_, _11269_);
  and (_11272_, _11271_, _05352_);
  or (_11273_, _11272_, _11268_);
  and (_11274_, _11273_, _05373_);
  or (_11275_, _11274_, _11262_);
  and (_11276_, _11275_, _09566_);
  or (_11277_, _11276_, _11250_);
  and (_11278_, _11277_, _09581_);
  or (_11279_, _11278_, _11220_);
  and (_11281_, _11279_, _05363_);
  or (_11282_, _11281_, _11163_);
  or (_11284_, _11282_, _09739_);
  and (_11286_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and (_11288_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_11290_, _11288_, _11286_);
  and (_11292_, _11290_, _05352_);
  and (_11293_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_11295_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_11296_, _11295_, _11293_);
  and (_11298_, _11296_, _09527_);
  or (_11299_, _11298_, _11292_);
  or (_11301_, _11299_, _09540_);
  and (_11302_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and (_11303_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_11304_, _11303_, _11302_);
  and (_11306_, _11304_, _05352_);
  and (_11308_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_11309_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_11311_, _11309_, _11308_);
  and (_11313_, _11311_, _09527_);
  or (_11314_, _11313_, _11306_);
  or (_11315_, _11314_, _05373_);
  and (_11316_, _11315_, _09566_);
  and (_11318_, _11316_, _11301_);
  or (_11319_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_11321_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_11322_, _11321_, _09527_);
  and (_11323_, _11322_, _11319_);
  or (_11324_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_11326_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and (_11327_, _11326_, _05352_);
  and (_11328_, _11327_, _11324_);
  or (_11330_, _11328_, _11323_);
  or (_11332_, _11330_, _09540_);
  or (_11333_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_11334_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_11335_, _11334_, _09527_);
  and (_11336_, _11335_, _11333_);
  or (_11337_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_11338_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_11339_, _11338_, _05352_);
  and (_11340_, _11339_, _11337_);
  or (_11341_, _11340_, _11336_);
  or (_11342_, _11341_, _05373_);
  and (_11343_, _11342_, _05379_);
  and (_11345_, _11343_, _11332_);
  or (_11347_, _11345_, _11318_);
  and (_11348_, _11347_, _09581_);
  and (_11349_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and (_11350_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_11351_, _11350_, _09527_);
  or (_11353_, _11351_, _11349_);
  and (_11354_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_11357_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_11358_, _11357_, _05352_);
  or (_11359_, _11358_, _11354_);
  and (_11360_, _11359_, _11353_);
  or (_11361_, _11360_, _09540_);
  and (_11362_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_11363_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_11365_, _11363_, _09527_);
  or (_11367_, _11365_, _11362_);
  and (_11368_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_11369_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_11371_, _11369_, _05352_);
  or (_11373_, _11371_, _11368_);
  and (_11374_, _11373_, _11367_);
  or (_11375_, _11374_, _05373_);
  and (_11376_, _11375_, _09566_);
  and (_11377_, _11376_, _11361_);
  or (_11378_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_11379_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and (_11381_, _11379_, _11378_);
  or (_11383_, _11381_, _05352_);
  or (_11384_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_11385_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_11387_, _11385_, _11384_);
  or (_11389_, _11387_, _09527_);
  and (_11390_, _11389_, _11383_);
  or (_11391_, _11390_, _09540_);
  or (_11393_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_11395_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_11396_, _11395_, _11393_);
  or (_11398_, _11396_, _05352_);
  or (_11399_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_11400_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and (_11401_, _11400_, _11399_);
  or (_11402_, _11401_, _09527_);
  and (_11404_, _11402_, _11398_);
  or (_11406_, _11404_, _05373_);
  and (_11407_, _11406_, _05379_);
  and (_11409_, _11407_, _11391_);
  or (_11411_, _11409_, _11377_);
  and (_11413_, _11411_, _05361_);
  or (_11414_, _11413_, _11348_);
  and (_11415_, _11414_, _09682_);
  and (_11416_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_11417_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_11418_, _11417_, _11416_);
  and (_11419_, _11418_, _09527_);
  and (_11420_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and (_11421_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_11423_, _11421_, _11420_);
  and (_11425_, _11423_, _05352_);
  or (_11426_, _11425_, _11419_);
  and (_11427_, _11426_, _05373_);
  and (_11429_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_11430_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_11432_, _11430_, _11429_);
  and (_11433_, _11432_, _09527_);
  and (_11434_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_11436_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_11437_, _11436_, _11434_);
  and (_11438_, _11437_, _05352_);
  or (_11439_, _11438_, _11433_);
  and (_11440_, _11439_, _09540_);
  or (_11441_, _11440_, _11427_);
  and (_11442_, _11441_, _09566_);
  or (_11443_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_11444_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_11445_, _11444_, _11443_);
  and (_11446_, _11445_, _09527_);
  or (_11448_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_11449_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_11451_, _11449_, _11448_);
  and (_11452_, _11451_, _05352_);
  or (_11453_, _11452_, _11446_);
  and (_11454_, _11453_, _05373_);
  or (_11455_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_11456_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_11457_, _11456_, _11455_);
  and (_11458_, _11457_, _09527_);
  or (_11459_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_11461_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_11462_, _11461_, _11459_);
  and (_11463_, _11462_, _05352_);
  or (_11464_, _11463_, _11458_);
  and (_11465_, _11464_, _09540_);
  or (_11466_, _11465_, _11454_);
  and (_11467_, _11466_, _05379_);
  or (_11468_, _11467_, _11442_);
  and (_11469_, _11468_, _05361_);
  and (_11470_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_11471_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_11472_, _11471_, _11470_);
  and (_11473_, _11472_, _09527_);
  and (_11474_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_11475_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_11476_, _11475_, _11474_);
  and (_11477_, _11476_, _05352_);
  or (_11478_, _11477_, _11473_);
  and (_11479_, _11478_, _05373_);
  and (_11480_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_11481_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_11483_, _11481_, _11480_);
  and (_11484_, _11483_, _09527_);
  and (_11486_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_11487_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_11488_, _11487_, _11486_);
  and (_11489_, _11488_, _05352_);
  or (_11491_, _11489_, _11484_);
  and (_11493_, _11491_, _09540_);
  or (_11494_, _11493_, _11479_);
  and (_11496_, _11494_, _09566_);
  or (_11497_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_11498_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_11499_, _11498_, _11497_);
  and (_11500_, _11499_, _09527_);
  or (_11502_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_11503_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_11504_, _11503_, _11502_);
  and (_11505_, _11504_, _05352_);
  or (_11506_, _11505_, _11500_);
  and (_11507_, _11506_, _05373_);
  or (_11508_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_11509_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_11511_, _11509_, _11508_);
  and (_11512_, _11511_, _09527_);
  or (_11513_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_11514_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_11515_, _11514_, _11513_);
  and (_11517_, _11515_, _05352_);
  or (_11518_, _11517_, _11512_);
  and (_11519_, _11518_, _09540_);
  or (_11520_, _11519_, _11507_);
  and (_11521_, _11520_, _05379_);
  or (_11522_, _11521_, _11496_);
  and (_11524_, _11522_, _09581_);
  or (_11525_, _11524_, _11469_);
  and (_11526_, _11525_, _05363_);
  or (_11527_, _11526_, _11415_);
  or (_11528_, _11527_, _05357_);
  and (_11530_, _11528_, _04360_);
  and (_11531_, _11530_, _11284_);
  or (_11533_, _11531_, _11029_);
  or (_11535_, _11533_, _05401_);
  or (_11537_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_11538_, _11537_, _22761_);
  and (_03190_, _11538_, _11535_);
  and (_11539_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  and (_11540_, _09509_, _23589_);
  or (_03194_, _11540_, _11539_);
  and (_11541_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_11542_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_11543_, _11542_, _11541_);
  and (_11544_, _11543_, _05352_);
  and (_11545_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_11546_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_11547_, _11546_, _11545_);
  and (_11548_, _11547_, _09527_);
  or (_11549_, _11548_, _11544_);
  or (_11551_, _11549_, _09540_);
  and (_11552_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_11553_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_11555_, _11553_, _11552_);
  and (_11556_, _11555_, _05352_);
  and (_11557_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_11559_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_11560_, _11559_, _11557_);
  and (_11562_, _11560_, _09527_);
  or (_11564_, _11562_, _11556_);
  or (_11565_, _11564_, _05373_);
  and (_11566_, _11565_, _09566_);
  and (_11568_, _11566_, _11551_);
  or (_11570_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_11571_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_11572_, _11571_, _09527_);
  and (_11573_, _11572_, _11570_);
  or (_11575_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_11576_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and (_11578_, _11576_, _05352_);
  and (_11579_, _11578_, _11575_);
  or (_11580_, _11579_, _11573_);
  or (_11581_, _11580_, _09540_);
  or (_11582_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_11583_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_11584_, _11583_, _09527_);
  and (_11585_, _11584_, _11582_);
  or (_11587_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_11589_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and (_11590_, _11589_, _05352_);
  and (_11592_, _11590_, _11587_);
  or (_11593_, _11592_, _11585_);
  or (_11594_, _11593_, _05373_);
  and (_11595_, _11594_, _05379_);
  and (_11596_, _11595_, _11581_);
  or (_11598_, _11596_, _11568_);
  or (_11599_, _11598_, _05361_);
  and (_11600_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_11601_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_11602_, _11601_, _09527_);
  or (_11604_, _11602_, _11600_);
  and (_11606_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_11607_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_11608_, _11607_, _05352_);
  or (_11609_, _11608_, _11606_);
  and (_11611_, _11609_, _11604_);
  or (_11612_, _11611_, _09540_);
  and (_11613_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and (_11614_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_11615_, _11614_, _09527_);
  or (_11616_, _11615_, _11613_);
  and (_11617_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_11618_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_11619_, _11618_, _05352_);
  or (_11620_, _11619_, _11617_);
  and (_11621_, _11620_, _11616_);
  or (_11622_, _11621_, _05373_);
  and (_11623_, _11622_, _09566_);
  and (_11624_, _11623_, _11612_);
  or (_11625_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_11626_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_11627_, _11626_, _11625_);
  or (_11628_, _11627_, _05352_);
  or (_11629_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_11630_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_11631_, _11630_, _11629_);
  or (_11632_, _11631_, _09527_);
  and (_11633_, _11632_, _11628_);
  or (_11634_, _11633_, _09540_);
  or (_11635_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_11636_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_11637_, _11636_, _11635_);
  or (_11640_, _11637_, _05352_);
  or (_11641_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_11643_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_11645_, _11643_, _11641_);
  or (_11647_, _11645_, _09527_);
  and (_11648_, _11647_, _11640_);
  or (_11649_, _11648_, _05373_);
  and (_11651_, _11649_, _05379_);
  and (_11652_, _11651_, _11634_);
  or (_11653_, _11652_, _11624_);
  or (_11655_, _11653_, _09581_);
  and (_11656_, _11655_, _09682_);
  and (_11657_, _11656_, _11599_);
  and (_11658_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_11659_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_11660_, _11659_, _11658_);
  and (_11661_, _11660_, _09527_);
  and (_11662_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_11663_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_11664_, _11663_, _11662_);
  and (_11665_, _11664_, _05352_);
  or (_11666_, _11665_, _11661_);
  and (_11667_, _11666_, _05373_);
  and (_11668_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_11669_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_11670_, _11669_, _11668_);
  and (_11671_, _11670_, _09527_);
  and (_11672_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_11673_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_11674_, _11673_, _11672_);
  and (_11675_, _11674_, _05352_);
  or (_11676_, _11675_, _11671_);
  and (_11677_, _11676_, _09540_);
  or (_11678_, _11677_, _11667_);
  and (_11679_, _11678_, _09566_);
  or (_11681_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_11682_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_11683_, _11682_, _11681_);
  and (_11684_, _11683_, _09527_);
  or (_11686_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_11689_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_11690_, _11689_, _11686_);
  and (_11692_, _11690_, _05352_);
  or (_11693_, _11692_, _11684_);
  and (_11694_, _11693_, _05373_);
  or (_11695_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_11696_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_11697_, _11696_, _11695_);
  and (_11699_, _11697_, _09527_);
  or (_11700_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_11702_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_11704_, _11702_, _11700_);
  and (_11705_, _11704_, _05352_);
  or (_11706_, _11705_, _11699_);
  and (_11707_, _11706_, _09540_);
  or (_11708_, _11707_, _11694_);
  and (_11709_, _11708_, _05379_);
  or (_11710_, _11709_, _11679_);
  and (_11711_, _11710_, _09581_);
  and (_11712_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_11713_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_11714_, _11713_, _11712_);
  and (_11715_, _11714_, _09527_);
  and (_11716_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_11717_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_11718_, _11717_, _11716_);
  and (_11719_, _11718_, _05352_);
  or (_11720_, _11719_, _11715_);
  and (_11722_, _11720_, _05373_);
  and (_11723_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_11724_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_11725_, _11724_, _11723_);
  and (_11726_, _11725_, _09527_);
  and (_11727_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and (_11728_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_11729_, _11728_, _11727_);
  and (_11730_, _11729_, _05352_);
  or (_11731_, _11730_, _11726_);
  and (_11733_, _11731_, _09540_);
  or (_11735_, _11733_, _11722_);
  and (_11736_, _11735_, _09566_);
  or (_11737_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_11738_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and (_11739_, _11738_, _11737_);
  and (_11740_, _11739_, _09527_);
  or (_11741_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_11742_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_11743_, _11742_, _11741_);
  and (_11744_, _11743_, _05352_);
  or (_11745_, _11744_, _11740_);
  and (_11747_, _11745_, _05373_);
  or (_11748_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_11749_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and (_11750_, _11749_, _11748_);
  and (_11751_, _11750_, _09527_);
  or (_11752_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_11754_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_11756_, _11754_, _11752_);
  and (_11758_, _11756_, _05352_);
  or (_11759_, _11758_, _11751_);
  and (_11760_, _11759_, _09540_);
  or (_11761_, _11760_, _11747_);
  and (_11763_, _11761_, _05379_);
  or (_11765_, _11763_, _11736_);
  and (_11767_, _11765_, _05361_);
  or (_11768_, _11767_, _11711_);
  and (_11769_, _11768_, _05363_);
  or (_11770_, _11769_, _11657_);
  or (_11771_, _11770_, _05357_);
  and (_11772_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_11773_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_11775_, _11773_, _11772_);
  and (_11776_, _11775_, _09527_);
  and (_11777_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_11778_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_11780_, _11778_, _11777_);
  and (_11781_, _11780_, _05352_);
  or (_11782_, _11781_, _11776_);
  or (_11783_, _11782_, _09540_);
  and (_11785_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_11787_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_11788_, _11787_, _11785_);
  and (_11789_, _11788_, _09527_);
  and (_11790_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_11791_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_11792_, _11791_, _11790_);
  and (_11793_, _11792_, _05352_);
  or (_11794_, _11793_, _11789_);
  or (_11795_, _11794_, _05373_);
  and (_11797_, _11795_, _09566_);
  and (_11799_, _11797_, _11783_);
  or (_11800_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_11801_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_11802_, _11801_, _05352_);
  and (_11804_, _11802_, _11800_);
  or (_11805_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_11806_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_11807_, _11806_, _09527_);
  and (_11809_, _11807_, _11805_);
  or (_11810_, _11809_, _11804_);
  or (_11812_, _11810_, _09540_);
  or (_11813_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_11814_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and (_11815_, _11814_, _05352_);
  and (_11817_, _11815_, _11813_);
  or (_11818_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_11819_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and (_11820_, _11819_, _09527_);
  and (_11821_, _11820_, _11818_);
  or (_11822_, _11821_, _11817_);
  or (_11823_, _11822_, _05373_);
  and (_11824_, _11823_, _05379_);
  and (_11825_, _11824_, _11812_);
  or (_11826_, _11825_, _11799_);
  and (_11827_, _11826_, _09581_);
  and (_11828_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_11829_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_11830_, _11829_, _11828_);
  and (_11831_, _11830_, _09527_);
  and (_11832_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_11833_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_11834_, _11833_, _11832_);
  and (_11835_, _11834_, _05352_);
  or (_11836_, _11835_, _11831_);
  or (_11838_, _11836_, _09540_);
  and (_11840_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_11842_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_11843_, _11842_, _11840_);
  and (_11844_, _11843_, _09527_);
  and (_11845_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_11846_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_11848_, _11846_, _11845_);
  and (_11849_, _11848_, _05352_);
  or (_11850_, _11849_, _11844_);
  or (_11851_, _11850_, _05373_);
  and (_11852_, _11851_, _09566_);
  and (_11854_, _11852_, _11838_);
  or (_11855_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_11857_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_11858_, _11857_, _11855_);
  and (_11860_, _11858_, _09527_);
  or (_11861_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_11862_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_11863_, _11862_, _11861_);
  and (_11865_, _11863_, _05352_);
  or (_11866_, _11865_, _11860_);
  or (_11867_, _11866_, _09540_);
  or (_11868_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_11870_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_11871_, _11870_, _11868_);
  and (_11872_, _11871_, _09527_);
  or (_11873_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_11874_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_11875_, _11874_, _11873_);
  and (_11876_, _11875_, _05352_);
  or (_11878_, _11876_, _11872_);
  or (_11880_, _11878_, _05373_);
  and (_11881_, _11880_, _05379_);
  and (_11883_, _11881_, _11867_);
  or (_11884_, _11883_, _11854_);
  and (_11885_, _11884_, _05361_);
  or (_11887_, _11885_, _11827_);
  and (_11889_, _11887_, _09682_);
  or (_11890_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_11892_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and (_11893_, _11892_, _11890_);
  and (_11894_, _11893_, _09527_);
  or (_11895_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_11896_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_11897_, _11896_, _11895_);
  and (_11899_, _11897_, _05352_);
  or (_11900_, _11899_, _11894_);
  and (_11901_, _11900_, _09540_);
  or (_11902_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_11903_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_11904_, _11903_, _11902_);
  and (_11905_, _11904_, _09527_);
  or (_11906_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_11907_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_11908_, _11907_, _11906_);
  and (_11909_, _11908_, _05352_);
  or (_11910_, _11909_, _11905_);
  and (_11912_, _11910_, _05373_);
  or (_11914_, _11912_, _11901_);
  and (_11916_, _11914_, _05379_);
  and (_11918_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and (_11920_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_11922_, _11920_, _11918_);
  and (_11923_, _11922_, _09527_);
  and (_11924_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and (_11925_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_11926_, _11925_, _11924_);
  and (_11927_, _11926_, _05352_);
  or (_11928_, _11927_, _11923_);
  and (_11929_, _11928_, _09540_);
  and (_11930_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and (_11931_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_11932_, _11931_, _11930_);
  and (_11933_, _11932_, _09527_);
  and (_11934_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_11936_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_11937_, _11936_, _11934_);
  and (_11938_, _11937_, _05352_);
  or (_11939_, _11938_, _11933_);
  and (_11940_, _11939_, _05373_);
  or (_11942_, _11940_, _11929_);
  and (_11944_, _11942_, _09566_);
  or (_11946_, _11944_, _11916_);
  and (_11948_, _11946_, _05361_);
  or (_11950_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_11951_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_11953_, _11951_, _05352_);
  and (_11954_, _11953_, _11950_);
  or (_11956_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_11958_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_11959_, _11958_, _09527_);
  and (_11960_, _11959_, _11956_);
  or (_11961_, _11960_, _11954_);
  and (_11963_, _11961_, _09540_);
  or (_11964_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_11965_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_11966_, _11965_, _05352_);
  and (_11967_, _11966_, _11964_);
  or (_11968_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_11969_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and (_11970_, _11969_, _09527_);
  and (_11971_, _11970_, _11968_);
  or (_11973_, _11971_, _11967_);
  and (_11975_, _11973_, _05373_);
  or (_11976_, _11975_, _11963_);
  and (_11978_, _11976_, _05379_);
  and (_11979_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and (_11980_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_11981_, _11980_, _11979_);
  and (_11982_, _11981_, _09527_);
  and (_11984_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_11986_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_11987_, _11986_, _11984_);
  and (_11989_, _11987_, _05352_);
  or (_11991_, _11989_, _11982_);
  and (_11993_, _11991_, _09540_);
  and (_11994_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_11995_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_11997_, _11995_, _11994_);
  and (_11999_, _11997_, _09527_);
  and (_12001_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_12003_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_12004_, _12003_, _12001_);
  and (_12006_, _12004_, _05352_);
  or (_12007_, _12006_, _11999_);
  and (_12008_, _12007_, _05373_);
  or (_12010_, _12008_, _11993_);
  and (_12011_, _12010_, _09566_);
  or (_12012_, _12011_, _11978_);
  and (_12013_, _12012_, _09581_);
  or (_12014_, _12013_, _11948_);
  and (_12015_, _12014_, _05363_);
  or (_12016_, _12015_, _11889_);
  or (_12017_, _12016_, _09739_);
  and (_12018_, _12017_, _11771_);
  or (_12019_, _12018_, _26838_);
  and (_12020_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_12021_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_12022_, _12021_, _12020_);
  and (_12023_, _12022_, _09527_);
  and (_12024_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_12025_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_12026_, _12025_, _12024_);
  and (_12027_, _12026_, _05352_);
  or (_12029_, _12027_, _12023_);
  or (_12031_, _12029_, _09540_);
  and (_12032_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_12033_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_12034_, _12033_, _12032_);
  and (_12035_, _12034_, _09527_);
  and (_12036_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_12037_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_12038_, _12037_, _12036_);
  and (_12039_, _12038_, _05352_);
  or (_12040_, _12039_, _12035_);
  or (_12041_, _12040_, _05373_);
  and (_12042_, _12041_, _09566_);
  and (_12043_, _12042_, _12031_);
  or (_12044_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_12046_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_12047_, _12046_, _12044_);
  and (_12048_, _12047_, _09527_);
  or (_12049_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_12050_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_12051_, _12050_, _12049_);
  and (_12052_, _12051_, _05352_);
  or (_12053_, _12052_, _12048_);
  or (_12054_, _12053_, _09540_);
  or (_12055_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_12056_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_12057_, _12056_, _12055_);
  and (_12058_, _12057_, _09527_);
  or (_12059_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_12060_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_12061_, _12060_, _12059_);
  and (_12062_, _12061_, _05352_);
  or (_12063_, _12062_, _12058_);
  or (_12064_, _12063_, _05373_);
  and (_12065_, _12064_, _05379_);
  and (_12066_, _12065_, _12054_);
  or (_12067_, _12066_, _12043_);
  and (_12068_, _12067_, _05361_);
  and (_12069_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_12070_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_12071_, _12070_, _12069_);
  and (_12072_, _12071_, _09527_);
  and (_12073_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_12074_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_12075_, _12074_, _12073_);
  and (_12076_, _12075_, _05352_);
  or (_12077_, _12076_, _12072_);
  or (_12078_, _12077_, _09540_);
  and (_12079_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_12080_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_12081_, _12080_, _12079_);
  and (_12082_, _12081_, _09527_);
  and (_12083_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_12084_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_12085_, _12084_, _12083_);
  and (_12086_, _12085_, _05352_);
  or (_12087_, _12086_, _12082_);
  or (_12088_, _12087_, _05373_);
  and (_12089_, _12088_, _09566_);
  and (_12090_, _12089_, _12078_);
  or (_12091_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_12092_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_12093_, _12092_, _05352_);
  and (_12094_, _12093_, _12091_);
  or (_12095_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_12097_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_12098_, _12097_, _09527_);
  and (_12099_, _12098_, _12095_);
  or (_12100_, _12099_, _12094_);
  or (_12101_, _12100_, _09540_);
  or (_12102_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_12103_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_12104_, _12103_, _05352_);
  and (_12105_, _12104_, _12102_);
  or (_12106_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_12107_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_12108_, _12107_, _09527_);
  and (_12110_, _12108_, _12106_);
  or (_12111_, _12110_, _12105_);
  or (_12112_, _12111_, _05373_);
  and (_12113_, _12112_, _05379_);
  and (_12114_, _12113_, _12101_);
  or (_12115_, _12114_, _12090_);
  and (_12116_, _12115_, _09581_);
  or (_12117_, _12116_, _12068_);
  and (_12118_, _12117_, _09682_);
  and (_12119_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_12120_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_12121_, _12120_, _12119_);
  and (_12122_, _12121_, _09527_);
  and (_12123_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_12124_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_12125_, _12124_, _12123_);
  and (_12126_, _12125_, _05352_);
  or (_12127_, _12126_, _12122_);
  and (_12128_, _12127_, _05373_);
  and (_12129_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_12130_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_12131_, _12130_, _12129_);
  and (_12132_, _12131_, _09527_);
  and (_12133_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_12134_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_12135_, _12134_, _12133_);
  and (_12136_, _12135_, _05352_);
  or (_12137_, _12136_, _12132_);
  and (_12138_, _12137_, _09540_);
  or (_12139_, _12138_, _12128_);
  and (_12140_, _12139_, _09566_);
  or (_12141_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_12142_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_12143_, _12142_, _05352_);
  and (_12144_, _12143_, _12141_);
  or (_12145_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_12146_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_12147_, _12146_, _09527_);
  and (_12148_, _12147_, _12145_);
  or (_12149_, _12148_, _12144_);
  and (_12150_, _12149_, _05373_);
  or (_12151_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_12152_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_12154_, _12152_, _05352_);
  and (_12155_, _12154_, _12151_);
  or (_12156_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_12157_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_12159_, _12157_, _09527_);
  and (_12161_, _12159_, _12156_);
  or (_12163_, _12161_, _12155_);
  and (_12165_, _12163_, _09540_);
  or (_12166_, _12165_, _12150_);
  and (_12168_, _12166_, _05379_);
  or (_12170_, _12168_, _12140_);
  and (_12171_, _12170_, _09581_);
  and (_12173_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_12174_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_12176_, _12174_, _12173_);
  and (_12177_, _12176_, _09527_);
  and (_12178_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_12179_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_12180_, _12179_, _12178_);
  and (_12181_, _12180_, _05352_);
  or (_12182_, _12181_, _12177_);
  and (_12183_, _12182_, _05373_);
  and (_12184_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_12185_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_12187_, _12185_, _12184_);
  and (_12188_, _12187_, _09527_);
  and (_12189_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_12190_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_12192_, _12190_, _12189_);
  and (_12193_, _12192_, _05352_);
  or (_12194_, _12193_, _12188_);
  and (_12195_, _12194_, _09540_);
  or (_12196_, _12195_, _12183_);
  and (_12197_, _12196_, _09566_);
  or (_12199_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_12200_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_12201_, _12200_, _12199_);
  and (_12202_, _12201_, _09527_);
  or (_12203_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_12204_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_12205_, _12204_, _12203_);
  and (_12206_, _12205_, _05352_);
  or (_12207_, _12206_, _12202_);
  and (_12208_, _12207_, _05373_);
  or (_12209_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_12210_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_12212_, _12210_, _12209_);
  and (_12213_, _12212_, _09527_);
  or (_12214_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_12215_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_12216_, _12215_, _12214_);
  and (_12217_, _12216_, _05352_);
  or (_12218_, _12217_, _12213_);
  and (_12220_, _12218_, _09540_);
  or (_12221_, _12220_, _12208_);
  and (_12222_, _12221_, _05379_);
  or (_12223_, _12222_, _12197_);
  and (_12224_, _12223_, _05361_);
  or (_12225_, _12224_, _12171_);
  and (_12226_, _12225_, _05363_);
  or (_12227_, _12226_, _12118_);
  or (_12228_, _12227_, _05357_);
  and (_12229_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_12230_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_12231_, _12230_, _12229_);
  and (_12232_, _12231_, _09527_);
  and (_12233_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_12234_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_12235_, _12234_, _12233_);
  and (_12236_, _12235_, _05352_);
  or (_12237_, _12236_, _12232_);
  or (_12239_, _12237_, _09540_);
  and (_12240_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_12241_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_12242_, _12241_, _12240_);
  and (_12243_, _12242_, _09527_);
  and (_12244_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_12245_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_12246_, _12245_, _12244_);
  and (_12247_, _12246_, _05352_);
  or (_12248_, _12247_, _12243_);
  or (_12249_, _12248_, _05373_);
  and (_12250_, _12249_, _09566_);
  and (_12251_, _12250_, _12239_);
  or (_12252_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_12253_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_12254_, _12253_, _05352_);
  and (_12255_, _12254_, _12252_);
  or (_12256_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_12257_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_12258_, _12257_, _09527_);
  and (_12259_, _12258_, _12256_);
  or (_12260_, _12259_, _12255_);
  or (_12261_, _12260_, _09540_);
  or (_12262_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_12263_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_12264_, _12263_, _05352_);
  and (_12265_, _12264_, _12262_);
  or (_12266_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_12267_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_12268_, _12267_, _09527_);
  and (_12269_, _12268_, _12266_);
  or (_12270_, _12269_, _12265_);
  or (_12271_, _12270_, _05373_);
  and (_12272_, _12271_, _05379_);
  and (_12273_, _12272_, _12261_);
  or (_12274_, _12273_, _12251_);
  and (_12275_, _12274_, _09581_);
  and (_12276_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_12277_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_12278_, _12277_, _12276_);
  and (_12279_, _12278_, _09527_);
  and (_12280_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_12281_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_12282_, _12281_, _12280_);
  and (_12283_, _12282_, _05352_);
  or (_12284_, _12283_, _12279_);
  or (_12285_, _12284_, _09540_);
  and (_12286_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_12287_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_12288_, _12287_, _12286_);
  and (_12289_, _12288_, _09527_);
  and (_12290_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_12291_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_12292_, _12291_, _12290_);
  and (_12293_, _12292_, _05352_);
  or (_12294_, _12293_, _12289_);
  or (_12295_, _12294_, _05373_);
  and (_12296_, _12295_, _09566_);
  and (_12297_, _12296_, _12285_);
  or (_12298_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_12300_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_12301_, _12300_, _12298_);
  and (_12302_, _12301_, _09527_);
  or (_12303_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_12304_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_12305_, _12304_, _12303_);
  and (_12306_, _12305_, _05352_);
  or (_12307_, _12306_, _12302_);
  or (_12308_, _12307_, _09540_);
  or (_12309_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_12310_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_12311_, _12310_, _12309_);
  and (_12312_, _12311_, _09527_);
  or (_12313_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_12314_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_12315_, _12314_, _12313_);
  and (_12316_, _12315_, _05352_);
  or (_12317_, _12316_, _12312_);
  or (_12318_, _12317_, _05373_);
  and (_12319_, _12318_, _05379_);
  and (_12320_, _12319_, _12308_);
  or (_12321_, _12320_, _12297_);
  and (_12322_, _12321_, _05361_);
  or (_12323_, _12322_, _12275_);
  and (_12324_, _12323_, _09682_);
  or (_12325_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_12326_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_12327_, _12326_, _12325_);
  and (_12328_, _12327_, _09527_);
  or (_12329_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_12330_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_12331_, _12330_, _12329_);
  and (_12332_, _12331_, _05352_);
  or (_12333_, _12332_, _12328_);
  and (_12334_, _12333_, _09540_);
  or (_12335_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_12336_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_12337_, _12336_, _12335_);
  and (_12338_, _12337_, _09527_);
  or (_12339_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_12340_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_12341_, _12340_, _12339_);
  and (_12342_, _12341_, _05352_);
  or (_12343_, _12342_, _12338_);
  and (_12344_, _12343_, _05373_);
  or (_12345_, _12344_, _12334_);
  and (_12346_, _12345_, _05379_);
  and (_12347_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_12348_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_12349_, _12348_, _12347_);
  and (_12350_, _12349_, _09527_);
  and (_12351_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_12352_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_12353_, _12352_, _12351_);
  and (_12354_, _12353_, _05352_);
  or (_12355_, _12354_, _12350_);
  and (_12356_, _12355_, _09540_);
  and (_12357_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_12358_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_12359_, _12358_, _12357_);
  and (_12360_, _12359_, _09527_);
  and (_12361_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_12362_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_12363_, _12362_, _12361_);
  and (_12364_, _12363_, _05352_);
  or (_12365_, _12364_, _12360_);
  and (_12366_, _12365_, _05373_);
  or (_12367_, _12366_, _12356_);
  and (_12368_, _12367_, _09566_);
  or (_12369_, _12368_, _12346_);
  and (_12370_, _12369_, _05361_);
  or (_12372_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_12373_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and (_12374_, _12373_, _05352_);
  and (_12375_, _12374_, _12372_);
  or (_12376_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_12377_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and (_12378_, _12377_, _09527_);
  and (_12379_, _12378_, _12376_);
  or (_12380_, _12379_, _12375_);
  and (_12381_, _12380_, _09540_);
  or (_12382_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_12383_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and (_12384_, _12383_, _05352_);
  and (_12385_, _12384_, _12382_);
  or (_12386_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_12387_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and (_12388_, _12387_, _09527_);
  and (_12389_, _12388_, _12386_);
  or (_12390_, _12389_, _12385_);
  and (_12391_, _12390_, _05373_);
  or (_12392_, _12391_, _12381_);
  and (_12393_, _12392_, _05379_);
  and (_12394_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and (_12395_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_12396_, _12395_, _12394_);
  and (_12397_, _12396_, _09527_);
  and (_12398_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and (_12399_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_12400_, _12399_, _12398_);
  and (_12401_, _12400_, _05352_);
  or (_12402_, _12401_, _12397_);
  and (_12403_, _12402_, _09540_);
  and (_12405_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and (_12406_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_12407_, _12406_, _12405_);
  and (_12408_, _12407_, _09527_);
  and (_12409_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and (_12410_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_12411_, _12410_, _12409_);
  and (_12412_, _12411_, _05352_);
  or (_12413_, _12412_, _12408_);
  and (_12414_, _12413_, _05373_);
  or (_12415_, _12414_, _12403_);
  and (_12416_, _12415_, _09566_);
  or (_12417_, _12416_, _12393_);
  and (_12418_, _12417_, _09581_);
  or (_12419_, _12418_, _12370_);
  and (_12420_, _12419_, _05363_);
  or (_12421_, _12420_, _12324_);
  or (_12422_, _12421_, _09739_);
  and (_12424_, _12422_, _12228_);
  or (_12425_, _12424_, _04360_);
  and (_12426_, _12425_, _12019_);
  or (_12427_, _12426_, _05401_);
  or (_12428_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_12429_, _12428_, _22761_);
  and (_03197_, _12429_, _12427_);
  and (_12430_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  and (_12431_, _10557_, _23635_);
  or (_03200_, _12431_, _12430_);
  and (_12432_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  and (_12433_, _02840_, _23982_);
  or (_27100_, _12433_, _12432_);
  and (_12435_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_12436_, _06040_, _23838_);
  or (_03209_, _12436_, _12435_);
  and (_12437_, _25301_, _23838_);
  and (_12438_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_03224_, _12438_, _12437_);
  and (_12439_, _02225_, _23718_);
  and (_12440_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_27089_, _12440_, _12439_);
  and (_12441_, _24089_, _23635_);
  and (_12442_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_03230_, _12442_, _12441_);
  and (_12443_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_12444_, _24559_, _23755_);
  or (_03240_, _12444_, _12443_);
  and (_12445_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  and (_12446_, _04734_, _23676_);
  or (_03243_, _12446_, _12445_);
  and (_12447_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and (_12448_, _25294_, _23838_);
  or (_03252_, _12448_, _12447_);
  and (_12450_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_12451_, _25619_, _23718_);
  or (_03258_, _12451_, _12450_);
  and (_12452_, _23864_, _23755_);
  and (_12453_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_03268_, _12453_, _12452_);
  and (_12455_, _06009_, _23676_);
  and (_12456_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_03289_, _12456_, _12455_);
  and (_12459_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and (_12460_, _25464_, _23718_);
  or (_27070_, _12460_, _12459_);
  and (_12461_, _03006_, _23676_);
  and (_12462_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or (_27082_, _12462_, _12461_);
  and (_12463_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and (_12465_, _10557_, _23676_);
  or (_03333_, _12465_, _12463_);
  and (_12466_, _02459_, _23589_);
  and (_12467_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or (_03339_, _12467_, _12466_);
  and (_12468_, _04733_, _23797_);
  not (_12469_, _12468_);
  and (_12470_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_12471_, _12468_, _23589_);
  or (_03342_, _12471_, _12470_);
  and (_12472_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_12473_, _12468_, _23755_);
  or (_03347_, _12473_, _12472_);
  and (_12474_, _03183_, _23849_);
  not (_12475_, _12474_);
  and (_12476_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_12477_, _12474_, _23791_);
  or (_03366_, _12477_, _12476_);
  and (_12478_, _03183_, _23803_);
  not (_12479_, _12478_);
  and (_12481_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_12482_, _12478_, _23718_);
  or (_03371_, _12482_, _12481_);
  and (_12484_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  and (_12485_, _10557_, _23838_);
  or (_03377_, _12485_, _12484_);
  and (_12486_, _03183_, _23842_);
  not (_12487_, _12486_);
  and (_12488_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  and (_12489_, _12486_, _23982_);
  or (_03387_, _12489_, _12488_);
  and (_12490_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  and (_12491_, _12486_, _23718_);
  or (_27138_, _12491_, _12490_);
  and (_03390_, t1_i, _22761_);
  and (_12492_, _03183_, _23854_);
  not (_12493_, _12492_);
  and (_12494_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and (_12496_, _12492_, _23589_);
  or (_03398_, _12496_, _12494_);
  and (_12498_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and (_12499_, _10557_, _23718_);
  or (_03401_, _12499_, _12498_);
  and (_12500_, _03183_, _23797_);
  not (_12501_, _12500_);
  and (_12502_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_12503_, _12500_, _23755_);
  or (_03419_, _12503_, _12502_);
  and (_12505_, _24078_, _23028_);
  and (_12507_, _12505_, _23982_);
  not (_12508_, _12505_);
  and (_12509_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_03422_, _12509_, _12507_);
  and (_12510_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_12511_, _12500_, _23718_);
  or (_03428_, _12511_, _12510_);
  and (_12512_, _03183_, _24768_);
  not (_12513_, _12512_);
  and (_12514_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_12515_, _12512_, _23589_);
  or (_03444_, _12515_, _12514_);
  and (_12516_, _05322_, _23797_);
  and (_12517_, _12516_, _23589_);
  not (_12519_, _12516_);
  and (_12520_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or (_03451_, _12520_, _12517_);
  and (_12521_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_12522_, _12512_, _23718_);
  or (_03458_, _12522_, _12521_);
  and (_26869_[0], _24409_, _22761_);
  and (_12524_, _03183_, _24541_);
  not (_12525_, _12524_);
  and (_12526_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and (_12527_, _12524_, _23755_);
  or (_03465_, _12527_, _12526_);
  and (_12528_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  and (_12529_, _12524_, _23838_);
  or (_03468_, _12529_, _12528_);
  and (_12530_, _03183_, _23641_);
  not (_12531_, _12530_);
  and (_12533_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  and (_12534_, _12530_, _23755_);
  or (_03481_, _12534_, _12533_);
  and (_12535_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_12536_, _12468_, _23718_);
  or (_03484_, _12536_, _12535_);
  and (_26869_[2], _24288_, _22761_);
  and (_12537_, _12505_, _23838_);
  and (_12538_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_03488_, _12538_, _12537_);
  and (_12539_, _03183_, _23863_);
  not (_12540_, _12539_);
  and (_12542_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  and (_12543_, _12539_, _23755_);
  or (_03500_, _12543_, _12542_);
  and (_12544_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_12545_, _12468_, _23791_);
  or (_03502_, _12545_, _12544_);
  and (_12547_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and (_12548_, _12539_, _23791_);
  or (_03520_, _12548_, _12547_);
  and (_12549_, _03183_, _24103_);
  not (_12550_, _12549_);
  and (_12551_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_12552_, _12549_, _23755_);
  or (_03523_, _12552_, _12551_);
  and (_12553_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_12554_, _12549_, _23676_);
  or (_03542_, _12554_, _12553_);
  and (_12556_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and (_12557_, _12524_, _23676_);
  or (_27134_, _12557_, _12556_);
  and (_12558_, _03183_, _24117_);
  not (_12560_, _12558_);
  and (_12561_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_12562_, _12558_, _23589_);
  or (_03551_, _12562_, _12561_);
  and (_12565_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_12566_, _12558_, _23635_);
  or (_27133_, _12566_, _12565_);
  and (_12567_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_12569_, _04776_, _23718_);
  or (_27033_, _12569_, _12567_);
  and (_12571_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_12572_, _12558_, _23718_);
  or (_03559_, _12572_, _12571_);
  and (_12573_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_12574_, _12468_, _23635_);
  or (_03561_, _12574_, _12573_);
  and (_12576_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_12577_, _12478_, _23982_);
  or (_03575_, _12577_, _12576_);
  and (_12579_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  and (_12580_, _12486_, _23755_);
  or (_03578_, _12580_, _12579_);
  and (_12581_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  and (_12582_, _12492_, _23982_);
  or (_03581_, _12582_, _12581_);
  and (_12583_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  and (_12584_, _12492_, _23791_);
  or (_03585_, _12584_, _12583_);
  and (_12585_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_12586_, _12468_, _23982_);
  or (_27029_, _12586_, _12585_);
  and (_12587_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_12588_, _12468_, _23838_);
  or (_03590_, _12588_, _12587_);
  and (_12589_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_12590_, _12512_, _23982_);
  or (_03598_, _12590_, _12589_);
  and (_12592_, _12505_, _23718_);
  and (_12593_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_27263_, _12593_, _12592_);
  and (_12595_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  and (_12597_, _12530_, _23791_);
  or (_27130_, _12597_, _12595_);
  and (_12599_, _04733_, _24768_);
  not (_12600_, _12599_);
  and (_12601_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_12603_, _12599_, _23838_);
  or (_03640_, _12603_, _12601_);
  and (_12605_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_12606_, _12549_, _23718_);
  or (_03642_, _12606_, _12605_);
  and (_12608_, _04692_, _23718_);
  and (_12609_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_03649_, _12609_, _12608_);
  and (_12610_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_12611_, _03657_, _23982_);
  or (_03661_, _12611_, _12610_);
  and (_12612_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_12613_, _12599_, _23635_);
  or (_03668_, _12613_, _12612_);
  and (_12615_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_12617_, _12599_, _23982_);
  or (_03673_, _12617_, _12615_);
  and (_12618_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_12619_, _12500_, _23838_);
  or (_03676_, _12619_, _12618_);
  nand (_12620_, _24311_, _22767_);
  or (_12621_, _22767_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_12622_, _12621_, _22761_);
  and (_26873_[3], _12622_, _12620_);
  and (_12624_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_12625_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_12627_, _12625_, _12624_);
  and (_12628_, _12627_, _05352_);
  and (_12629_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_12630_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_12632_, _12630_, _12629_);
  and (_12634_, _12632_, _09527_);
  or (_12635_, _12634_, _12628_);
  or (_12636_, _12635_, _09540_);
  and (_12637_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_12638_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_12639_, _12638_, _12637_);
  and (_12640_, _12639_, _05352_);
  and (_12641_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and (_12642_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_12644_, _12642_, _12641_);
  and (_12646_, _12644_, _09527_);
  or (_12648_, _12646_, _12640_);
  or (_12650_, _12648_, _05373_);
  and (_12651_, _12650_, _09566_);
  and (_12652_, _12651_, _12636_);
  or (_12653_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_12654_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_12655_, _12654_, _09527_);
  and (_12656_, _12655_, _12653_);
  or (_12657_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_12658_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and (_12659_, _12658_, _05352_);
  and (_12660_, _12659_, _12657_);
  or (_12661_, _12660_, _12656_);
  or (_12662_, _12661_, _09540_);
  or (_12663_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_12664_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_12665_, _12664_, _09527_);
  and (_12666_, _12665_, _12663_);
  or (_12667_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_12668_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and (_12669_, _12668_, _05352_);
  and (_12670_, _12669_, _12667_);
  or (_12671_, _12670_, _12666_);
  or (_12672_, _12671_, _05373_);
  and (_12673_, _12672_, _05379_);
  and (_12674_, _12673_, _12662_);
  or (_12675_, _12674_, _12652_);
  or (_12676_, _12675_, _05361_);
  and (_12677_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_12678_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_12679_, _12678_, _09527_);
  or (_12680_, _12679_, _12677_);
  and (_12681_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_12682_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_12683_, _12682_, _05352_);
  or (_12684_, _12683_, _12681_);
  and (_12685_, _12684_, _12680_);
  or (_12686_, _12685_, _09540_);
  and (_12687_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and (_12688_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_12689_, _12688_, _09527_);
  or (_12690_, _12689_, _12687_);
  and (_12691_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_12692_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_12693_, _12692_, _05352_);
  or (_12694_, _12693_, _12691_);
  and (_12695_, _12694_, _12690_);
  or (_12696_, _12695_, _05373_);
  and (_12697_, _12696_, _09566_);
  and (_12698_, _12697_, _12686_);
  or (_12699_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_12700_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_12701_, _12700_, _12699_);
  or (_12702_, _12701_, _05352_);
  or (_12703_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_12704_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_12705_, _12704_, _12703_);
  or (_12706_, _12705_, _09527_);
  and (_12707_, _12706_, _12702_);
  or (_12708_, _12707_, _09540_);
  or (_12709_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_12710_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and (_12711_, _12710_, _12709_);
  or (_12712_, _12711_, _05352_);
  or (_12713_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_12714_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_12715_, _12714_, _12713_);
  or (_12716_, _12715_, _09527_);
  and (_12717_, _12716_, _12712_);
  or (_12718_, _12717_, _05373_);
  and (_12719_, _12718_, _05379_);
  and (_12720_, _12719_, _12708_);
  or (_12721_, _12720_, _12698_);
  or (_12722_, _12721_, _09581_);
  and (_12723_, _12722_, _09682_);
  and (_12724_, _12723_, _12676_);
  and (_12725_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_12726_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_12727_, _12726_, _12725_);
  and (_12728_, _12727_, _09527_);
  and (_12729_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_12730_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_12731_, _12730_, _12729_);
  and (_12732_, _12731_, _05352_);
  or (_12733_, _12732_, _12728_);
  and (_12734_, _12733_, _05373_);
  and (_12735_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_12736_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_12737_, _12736_, _12735_);
  and (_12738_, _12737_, _09527_);
  and (_12739_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_12740_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_12741_, _12740_, _12739_);
  and (_12742_, _12741_, _05352_);
  or (_12743_, _12742_, _12738_);
  and (_12744_, _12743_, _09540_);
  or (_12745_, _12744_, _12734_);
  and (_12746_, _12745_, _09566_);
  or (_12747_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_12748_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_12749_, _12748_, _12747_);
  and (_12750_, _12749_, _09527_);
  or (_12751_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_12752_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_12753_, _12752_, _12751_);
  and (_12754_, _12753_, _05352_);
  or (_12755_, _12754_, _12750_);
  and (_12756_, _12755_, _05373_);
  or (_12757_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_12758_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_12759_, _12758_, _12757_);
  and (_12760_, _12759_, _09527_);
  or (_12761_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_12762_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_12763_, _12762_, _12761_);
  and (_12764_, _12763_, _05352_);
  or (_12765_, _12764_, _12760_);
  and (_12766_, _12765_, _09540_);
  or (_12767_, _12766_, _12756_);
  and (_12768_, _12767_, _05379_);
  or (_12769_, _12768_, _12746_);
  and (_12770_, _12769_, _09581_);
  and (_12771_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and (_12772_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_12773_, _12772_, _12771_);
  and (_12774_, _12773_, _09527_);
  and (_12775_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_12776_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_12777_, _12776_, _12775_);
  and (_12778_, _12777_, _05352_);
  or (_12779_, _12778_, _12774_);
  and (_12780_, _12779_, _05373_);
  and (_12781_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_12782_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_12783_, _12782_, _12781_);
  and (_12784_, _12783_, _09527_);
  and (_12785_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_12786_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_12787_, _12786_, _12785_);
  and (_12788_, _12787_, _05352_);
  or (_12789_, _12788_, _12784_);
  and (_12790_, _12789_, _09540_);
  or (_12791_, _12790_, _12780_);
  and (_12792_, _12791_, _09566_);
  or (_12793_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_12794_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and (_12795_, _12794_, _12793_);
  and (_12796_, _12795_, _09527_);
  or (_12797_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_12798_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_12799_, _12798_, _12797_);
  and (_12800_, _12799_, _05352_);
  or (_12801_, _12800_, _12796_);
  and (_12802_, _12801_, _05373_);
  or (_12803_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_12804_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_12805_, _12804_, _12803_);
  and (_12806_, _12805_, _09527_);
  or (_12807_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_12808_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_12809_, _12808_, _12807_);
  and (_12810_, _12809_, _05352_);
  or (_12811_, _12810_, _12806_);
  and (_12812_, _12811_, _09540_);
  or (_12813_, _12812_, _12802_);
  and (_12814_, _12813_, _05379_);
  or (_12815_, _12814_, _12792_);
  and (_12816_, _12815_, _05361_);
  or (_12817_, _12816_, _12770_);
  and (_12818_, _12817_, _05363_);
  or (_12819_, _12818_, _12724_);
  or (_12820_, _12819_, _05357_);
  and (_12821_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and (_12822_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_12823_, _12822_, _12821_);
  and (_12824_, _12823_, _09527_);
  and (_12825_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_12826_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_12827_, _12826_, _12825_);
  and (_12828_, _12827_, _05352_);
  or (_12829_, _12828_, _12824_);
  or (_12830_, _12829_, _09540_);
  and (_12831_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and (_12832_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_12833_, _12832_, _12831_);
  and (_12834_, _12833_, _09527_);
  and (_12835_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_12836_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_12837_, _12836_, _12835_);
  and (_12838_, _12837_, _05352_);
  or (_12839_, _12838_, _12834_);
  or (_12840_, _12839_, _05373_);
  and (_12841_, _12840_, _09566_);
  and (_12842_, _12841_, _12830_);
  or (_12843_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_12844_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_12845_, _12844_, _05352_);
  and (_12846_, _12845_, _12843_);
  or (_12847_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_12848_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_12849_, _12848_, _09527_);
  and (_12850_, _12849_, _12847_);
  or (_12851_, _12850_, _12846_);
  or (_12852_, _12851_, _09540_);
  or (_12853_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_12854_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_12855_, _12854_, _05352_);
  and (_12856_, _12855_, _12853_);
  or (_12857_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_12858_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and (_12859_, _12858_, _09527_);
  and (_12860_, _12859_, _12857_);
  or (_12861_, _12860_, _12856_);
  or (_12862_, _12861_, _05373_);
  and (_12863_, _12862_, _05379_);
  and (_12864_, _12863_, _12852_);
  or (_12865_, _12864_, _12842_);
  and (_12866_, _12865_, _09581_);
  and (_12867_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_12868_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_12869_, _12868_, _12867_);
  and (_12870_, _12869_, _09527_);
  and (_12871_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_12872_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_12873_, _12872_, _12871_);
  and (_12874_, _12873_, _05352_);
  or (_12875_, _12874_, _12870_);
  or (_12876_, _12875_, _09540_);
  and (_12877_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_12878_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_12879_, _12878_, _12877_);
  and (_12880_, _12879_, _09527_);
  and (_12881_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_12882_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_12883_, _12882_, _12881_);
  and (_12884_, _12883_, _05352_);
  or (_12885_, _12884_, _12880_);
  or (_12886_, _12885_, _05373_);
  and (_12887_, _12886_, _09566_);
  and (_12888_, _12887_, _12876_);
  or (_12889_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_12890_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_12891_, _12890_, _12889_);
  and (_12892_, _12891_, _09527_);
  or (_12893_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_12894_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_12895_, _12894_, _12893_);
  and (_12896_, _12895_, _05352_);
  or (_12897_, _12896_, _12892_);
  or (_12898_, _12897_, _09540_);
  or (_12899_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_12900_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_12901_, _12900_, _12899_);
  and (_12902_, _12901_, _09527_);
  or (_12903_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_12904_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_12905_, _12904_, _12903_);
  and (_12906_, _12905_, _05352_);
  or (_12907_, _12906_, _12902_);
  or (_12908_, _12907_, _05373_);
  and (_12909_, _12908_, _05379_);
  and (_12910_, _12909_, _12898_);
  or (_12911_, _12910_, _12888_);
  and (_12912_, _12911_, _05361_);
  or (_12913_, _12912_, _12866_);
  and (_12914_, _12913_, _09682_);
  or (_12915_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_12916_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_12917_, _12916_, _12915_);
  and (_12918_, _12917_, _09527_);
  or (_12919_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_12920_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and (_12921_, _12920_, _12919_);
  and (_12922_, _12921_, _05352_);
  or (_12923_, _12922_, _12918_);
  and (_12924_, _12923_, _09540_);
  or (_12925_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_12926_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_12927_, _12926_, _12925_);
  and (_12928_, _12927_, _09527_);
  or (_12929_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_12930_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and (_12931_, _12930_, _12929_);
  and (_12932_, _12931_, _05352_);
  or (_12933_, _12932_, _12928_);
  and (_12934_, _12933_, _05373_);
  or (_12935_, _12934_, _12924_);
  and (_12936_, _12935_, _05379_);
  and (_12937_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_12938_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_12939_, _12938_, _12937_);
  and (_12940_, _12939_, _09527_);
  and (_12941_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and (_12942_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_12943_, _12942_, _12941_);
  and (_12944_, _12943_, _05352_);
  or (_12945_, _12944_, _12940_);
  and (_12946_, _12945_, _09540_);
  and (_12947_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_12948_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_12949_, _12948_, _12947_);
  and (_12950_, _12949_, _09527_);
  and (_12951_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and (_12952_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_12953_, _12952_, _12951_);
  and (_12954_, _12953_, _05352_);
  or (_12955_, _12954_, _12950_);
  and (_12956_, _12955_, _05373_);
  or (_12957_, _12956_, _12946_);
  and (_12958_, _12957_, _09566_);
  or (_12959_, _12958_, _12936_);
  and (_12960_, _12959_, _05361_);
  or (_12961_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_12962_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and (_12963_, _12962_, _05352_);
  and (_12964_, _12963_, _12961_);
  or (_12965_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_12966_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and (_12967_, _12966_, _09527_);
  and (_12968_, _12967_, _12965_);
  or (_12969_, _12968_, _12964_);
  and (_12970_, _12969_, _09540_);
  or (_12971_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_12972_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and (_12973_, _12972_, _05352_);
  and (_12974_, _12973_, _12971_);
  or (_12975_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_12976_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and (_12977_, _12976_, _09527_);
  and (_12978_, _12977_, _12975_);
  or (_12979_, _12978_, _12974_);
  and (_12980_, _12979_, _05373_);
  or (_12981_, _12980_, _12970_);
  and (_12982_, _12981_, _05379_);
  and (_12983_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and (_12984_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_12985_, _12984_, _12983_);
  and (_12986_, _12985_, _09527_);
  and (_12987_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and (_12988_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_12989_, _12988_, _12987_);
  and (_12990_, _12989_, _05352_);
  or (_12991_, _12990_, _12986_);
  and (_12992_, _12991_, _09540_);
  and (_12993_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and (_12994_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_12995_, _12994_, _12993_);
  and (_12996_, _12995_, _09527_);
  and (_12997_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and (_12998_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_12999_, _12998_, _12997_);
  and (_13000_, _12999_, _05352_);
  or (_13001_, _13000_, _12996_);
  and (_13002_, _13001_, _05373_);
  or (_13003_, _13002_, _12992_);
  and (_13004_, _13003_, _09566_);
  or (_13005_, _13004_, _12982_);
  and (_13006_, _13005_, _09581_);
  or (_13007_, _13006_, _12960_);
  and (_13008_, _13007_, _05363_);
  or (_13009_, _13008_, _12914_);
  or (_13010_, _13009_, _09739_);
  and (_13011_, _13010_, _12820_);
  or (_13012_, _13011_, _26838_);
  and (_13013_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_13014_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_13015_, _13014_, _13013_);
  and (_13016_, _13015_, _09527_);
  and (_13017_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_13018_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_13019_, _13018_, _13017_);
  and (_13020_, _13019_, _05352_);
  or (_13021_, _13020_, _13016_);
  or (_13022_, _13021_, _09540_);
  and (_13023_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_13024_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_13025_, _13024_, _13023_);
  and (_13026_, _13025_, _09527_);
  and (_13027_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_13028_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_13029_, _13028_, _13027_);
  and (_13030_, _13029_, _05352_);
  or (_13031_, _13030_, _13026_);
  or (_13032_, _13031_, _05373_);
  and (_13033_, _13032_, _09566_);
  and (_13034_, _13033_, _13022_);
  or (_13035_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_13036_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_13037_, _13036_, _13035_);
  and (_13038_, _13037_, _09527_);
  or (_13039_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_13040_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_13041_, _13040_, _13039_);
  and (_13042_, _13041_, _05352_);
  or (_13043_, _13042_, _13038_);
  or (_13044_, _13043_, _09540_);
  or (_13045_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_13046_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_13047_, _13046_, _13045_);
  and (_13048_, _13047_, _09527_);
  or (_13049_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_13050_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_13051_, _13050_, _13049_);
  and (_13052_, _13051_, _05352_);
  or (_13053_, _13052_, _13048_);
  or (_13054_, _13053_, _05373_);
  and (_13055_, _13054_, _05379_);
  and (_13056_, _13055_, _13044_);
  or (_13057_, _13056_, _13034_);
  and (_13058_, _13057_, _05361_);
  and (_13059_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_13060_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_13061_, _13060_, _13059_);
  and (_13062_, _13061_, _09527_);
  and (_13063_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_13064_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_13065_, _13064_, _13063_);
  and (_13066_, _13065_, _05352_);
  or (_13067_, _13066_, _13062_);
  or (_13068_, _13067_, _09540_);
  and (_13069_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_13070_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_13071_, _13070_, _13069_);
  and (_13072_, _13071_, _09527_);
  and (_13073_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_13074_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_13075_, _13074_, _13073_);
  and (_13076_, _13075_, _05352_);
  or (_13077_, _13076_, _13072_);
  or (_13078_, _13077_, _05373_);
  and (_13079_, _13078_, _09566_);
  and (_13080_, _13079_, _13068_);
  or (_13081_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_13082_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_13083_, _13082_, _05352_);
  and (_13084_, _13083_, _13081_);
  or (_13085_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_13086_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_13087_, _13086_, _09527_);
  and (_13088_, _13087_, _13085_);
  or (_13089_, _13088_, _13084_);
  or (_13090_, _13089_, _09540_);
  or (_13091_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_13092_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_13093_, _13092_, _05352_);
  and (_13094_, _13093_, _13091_);
  or (_13095_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_13096_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_13097_, _13096_, _09527_);
  and (_13098_, _13097_, _13095_);
  or (_13099_, _13098_, _13094_);
  or (_13100_, _13099_, _05373_);
  and (_13101_, _13100_, _05379_);
  and (_13102_, _13101_, _13090_);
  or (_13103_, _13102_, _13080_);
  and (_13104_, _13103_, _09581_);
  or (_13105_, _13104_, _13058_);
  and (_13106_, _13105_, _09682_);
  and (_13107_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and (_13108_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_13109_, _13108_, _13107_);
  and (_13110_, _13109_, _09527_);
  and (_13111_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_13112_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_13113_, _13112_, _13111_);
  and (_13114_, _13113_, _05352_);
  or (_13115_, _13114_, _13110_);
  and (_13116_, _13115_, _05373_);
  and (_13117_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_13118_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_13119_, _13118_, _13117_);
  and (_13120_, _13119_, _09527_);
  and (_13121_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_13122_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_13123_, _13122_, _13121_);
  and (_13124_, _13123_, _05352_);
  or (_13125_, _13124_, _13120_);
  and (_13126_, _13125_, _09540_);
  or (_13127_, _13126_, _13116_);
  and (_13128_, _13127_, _09566_);
  or (_13129_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_13130_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_13131_, _13130_, _05352_);
  and (_13132_, _13131_, _13129_);
  or (_13133_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_13134_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_13135_, _13134_, _09527_);
  and (_13136_, _13135_, _13133_);
  or (_13137_, _13136_, _13132_);
  and (_13138_, _13137_, _05373_);
  or (_13139_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_13140_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and (_13141_, _13140_, _05352_);
  and (_13142_, _13141_, _13139_);
  or (_13143_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_13144_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_13145_, _13144_, _09527_);
  and (_13146_, _13145_, _13143_);
  or (_13147_, _13146_, _13142_);
  and (_13148_, _13147_, _09540_);
  or (_13149_, _13148_, _13138_);
  and (_13150_, _13149_, _05379_);
  or (_13151_, _13150_, _13128_);
  and (_13152_, _13151_, _09581_);
  and (_13153_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_13154_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_13155_, _13154_, _13153_);
  and (_13156_, _13155_, _09527_);
  and (_13157_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_13158_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_13159_, _13158_, _13157_);
  and (_13160_, _13159_, _05352_);
  or (_13161_, _13160_, _13156_);
  and (_13162_, _13161_, _05373_);
  and (_13163_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_13164_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_13165_, _13164_, _13163_);
  and (_13166_, _13165_, _09527_);
  and (_13167_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_13168_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_13169_, _13168_, _13167_);
  and (_13170_, _13169_, _05352_);
  or (_13171_, _13170_, _13166_);
  and (_13172_, _13171_, _09540_);
  or (_13173_, _13172_, _13162_);
  and (_13174_, _13173_, _09566_);
  or (_13175_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_13176_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_13177_, _13176_, _13175_);
  and (_13178_, _13177_, _09527_);
  or (_13179_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_13180_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_13181_, _13180_, _13179_);
  and (_13182_, _13181_, _05352_);
  or (_13183_, _13182_, _13178_);
  and (_13184_, _13183_, _05373_);
  or (_13185_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_13186_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_13187_, _13186_, _13185_);
  and (_13188_, _13187_, _09527_);
  or (_13189_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_13190_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_13191_, _13190_, _13189_);
  and (_13192_, _13191_, _05352_);
  or (_13193_, _13192_, _13188_);
  and (_13194_, _13193_, _09540_);
  or (_13195_, _13194_, _13184_);
  and (_13196_, _13195_, _05379_);
  or (_13197_, _13196_, _13174_);
  and (_13198_, _13197_, _05361_);
  or (_13199_, _13198_, _13152_);
  and (_13200_, _13199_, _05363_);
  or (_13201_, _13200_, _13106_);
  or (_13202_, _13201_, _05357_);
  and (_13203_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_13204_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_13205_, _13204_, _13203_);
  and (_13206_, _13205_, _09527_);
  and (_13207_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_13208_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_13209_, _13208_, _13207_);
  and (_13210_, _13209_, _05352_);
  or (_13211_, _13210_, _13206_);
  or (_13212_, _13211_, _09540_);
  and (_13213_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_13214_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_13215_, _13214_, _13213_);
  and (_13216_, _13215_, _09527_);
  and (_13217_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_13218_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_13219_, _13218_, _13217_);
  and (_13220_, _13219_, _05352_);
  or (_13221_, _13220_, _13216_);
  or (_13222_, _13221_, _05373_);
  and (_13223_, _13222_, _09566_);
  and (_13224_, _13223_, _13212_);
  or (_13225_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_13226_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_13227_, _13226_, _05352_);
  and (_13228_, _13227_, _13225_);
  or (_13229_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_13230_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_13231_, _13230_, _09527_);
  and (_13232_, _13231_, _13229_);
  or (_13233_, _13232_, _13228_);
  or (_13234_, _13233_, _09540_);
  or (_13235_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_13236_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_13237_, _13236_, _05352_);
  and (_13238_, _13237_, _13235_);
  or (_13239_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_13240_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_13241_, _13240_, _09527_);
  and (_13242_, _13241_, _13239_);
  or (_13243_, _13242_, _13238_);
  or (_13244_, _13243_, _05373_);
  and (_13245_, _13244_, _05379_);
  and (_13246_, _13245_, _13234_);
  or (_13247_, _13246_, _13224_);
  and (_13248_, _13247_, _09581_);
  and (_13249_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_13250_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_13251_, _13250_, _13249_);
  and (_13252_, _13251_, _09527_);
  and (_13253_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_13254_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_13255_, _13254_, _13253_);
  and (_13256_, _13255_, _05352_);
  or (_13257_, _13256_, _13252_);
  or (_13258_, _13257_, _09540_);
  and (_13259_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_13260_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_13261_, _13260_, _13259_);
  and (_13262_, _13261_, _09527_);
  and (_13263_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_13264_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_13265_, _13264_, _13263_);
  and (_13266_, _13265_, _05352_);
  or (_13267_, _13266_, _13262_);
  or (_13268_, _13267_, _05373_);
  and (_13269_, _13268_, _09566_);
  and (_13270_, _13269_, _13258_);
  or (_13271_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_13272_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_13273_, _13272_, _13271_);
  and (_13274_, _13273_, _09527_);
  or (_13275_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_13276_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_13277_, _13276_, _13275_);
  and (_13278_, _13277_, _05352_);
  or (_13279_, _13278_, _13274_);
  or (_13280_, _13279_, _09540_);
  or (_13281_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_13282_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_13283_, _13282_, _13281_);
  and (_13284_, _13283_, _09527_);
  or (_13285_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_13286_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_13287_, _13286_, _13285_);
  and (_13288_, _13287_, _05352_);
  or (_13289_, _13288_, _13284_);
  or (_13290_, _13289_, _05373_);
  and (_13291_, _13290_, _05379_);
  and (_13292_, _13291_, _13280_);
  or (_13293_, _13292_, _13270_);
  and (_13294_, _13293_, _05361_);
  or (_13295_, _13294_, _13248_);
  and (_13296_, _13295_, _09682_);
  or (_13297_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_13298_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_13299_, _13298_, _13297_);
  and (_13300_, _13299_, _09527_);
  or (_13301_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_13302_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_13303_, _13302_, _13301_);
  and (_13304_, _13303_, _05352_);
  or (_13305_, _13304_, _13300_);
  and (_13306_, _13305_, _09540_);
  or (_13307_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_13308_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_13309_, _13308_, _13307_);
  and (_13310_, _13309_, _09527_);
  or (_13311_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_13312_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_13313_, _13312_, _13311_);
  and (_13314_, _13313_, _05352_);
  or (_13315_, _13314_, _13310_);
  and (_13316_, _13315_, _05373_);
  or (_13317_, _13316_, _13306_);
  and (_13318_, _13317_, _05379_);
  and (_13319_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_13320_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_13321_, _13320_, _13319_);
  and (_13322_, _13321_, _09527_);
  and (_13323_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_13324_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_13325_, _13324_, _13323_);
  and (_13326_, _13325_, _05352_);
  or (_13327_, _13326_, _13322_);
  and (_13328_, _13327_, _09540_);
  and (_13329_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_13330_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_13331_, _13330_, _13329_);
  and (_13332_, _13331_, _09527_);
  and (_13333_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_13334_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_13335_, _13334_, _13333_);
  and (_13336_, _13335_, _05352_);
  or (_13337_, _13336_, _13332_);
  and (_13338_, _13337_, _05373_);
  or (_13339_, _13338_, _13328_);
  and (_13340_, _13339_, _09566_);
  or (_13341_, _13340_, _13318_);
  and (_13342_, _13341_, _05361_);
  or (_13343_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_13344_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_13345_, _13344_, _05352_);
  and (_13346_, _13345_, _13343_);
  or (_13347_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_13348_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_13349_, _13348_, _09527_);
  and (_13350_, _13349_, _13347_);
  or (_13351_, _13350_, _13346_);
  and (_13352_, _13351_, _09540_);
  or (_13353_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_13354_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_13355_, _13354_, _05352_);
  and (_13356_, _13355_, _13353_);
  or (_13357_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_13358_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_13359_, _13358_, _09527_);
  and (_13360_, _13359_, _13357_);
  or (_13361_, _13360_, _13356_);
  and (_13362_, _13361_, _05373_);
  or (_13363_, _13362_, _13352_);
  and (_13364_, _13363_, _05379_);
  and (_13365_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_13366_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_13367_, _13366_, _13365_);
  and (_13368_, _13367_, _09527_);
  and (_13369_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_13370_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_13371_, _13370_, _13369_);
  and (_13372_, _13371_, _05352_);
  or (_13373_, _13372_, _13368_);
  and (_13374_, _13373_, _09540_);
  and (_13375_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_13376_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_13377_, _13376_, _13375_);
  and (_13378_, _13377_, _09527_);
  and (_13379_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_13380_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_13381_, _13380_, _13379_);
  and (_13382_, _13381_, _05352_);
  or (_13383_, _13382_, _13378_);
  and (_13384_, _13383_, _05373_);
  or (_13385_, _13384_, _13374_);
  and (_13386_, _13385_, _09566_);
  or (_13387_, _13386_, _13364_);
  and (_13388_, _13387_, _09581_);
  or (_13389_, _13388_, _13342_);
  and (_13390_, _13389_, _05363_);
  or (_13391_, _13390_, _13296_);
  or (_13392_, _13391_, _09739_);
  and (_13393_, _13392_, _13202_);
  or (_13394_, _13393_, _04360_);
  and (_13395_, _13394_, _13012_);
  or (_13396_, _13395_, _05401_);
  or (_13397_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_13398_, _13397_, _22761_);
  and (_27317_[1], _13398_, _13396_);
  and (_13399_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_13400_, _03657_, _23838_);
  or (_03689_, _13400_, _13399_);
  and (_13401_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  and (_13402_, _12539_, _23838_);
  or (_03693_, _13402_, _13401_);
  and (_13403_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_13404_, _12558_, _23791_);
  or (_27132_, _13404_, _13403_);
  and (_13405_, _03134_, _23676_);
  and (_13406_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or (_03739_, _13406_, _13405_);
  and (_13407_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_13408_, _12599_, _23589_);
  or (_03741_, _13408_, _13407_);
  and (_13409_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  and (_13410_, _12530_, _23589_);
  or (_03748_, _13410_, _13409_);
  and (_13411_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_13412_, _12558_, _23676_);
  or (_03751_, _13412_, _13411_);
  and (_13413_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_13414_, _12599_, _23755_);
  or (_03762_, _13414_, _13413_);
  and (_13415_, _03134_, _23791_);
  and (_13416_, _03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or (_03765_, _13416_, _13415_);
  and (_13417_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_13418_, _12558_, _23838_);
  or (_03768_, _13418_, _13417_);
  and (_13419_, _03006_, _23838_);
  and (_13420_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or (_03771_, _13420_, _13419_);
  and (_03784_, t0_i, _22761_);
  and (_13421_, _02225_, _23755_);
  and (_13422_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_03786_, _13422_, _13421_);
  nand (_13423_, _02077_, _23914_);
  and (_13424_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_13425_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_13426_, _13425_, _13424_);
  or (_13427_, _13426_, _02077_);
  and (_13428_, _13427_, _04740_);
  and (_13429_, _13428_, _13423_);
  and (_13430_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_13431_, _13430_, _13429_);
  and (_03788_, _13431_, _22761_);
  and (_13432_, _03006_, _23791_);
  and (_13433_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or (_03807_, _13433_, _13432_);
  and (_13434_, _04733_, _24541_);
  not (_13435_, _13434_);
  and (_13436_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  and (_13437_, _13434_, _23635_);
  or (_03813_, _13437_, _13436_);
  or (_13438_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  not (_13439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_13440_, _02078_, _13439_);
  and (_13441_, _13440_, _13438_);
  and (_13442_, _13441_, _04740_);
  nor (_13443_, _04740_, _23784_);
  or (_13444_, _13443_, _13442_);
  and (_03815_, _13444_, _22761_);
  and (_13445_, _03006_, _23589_);
  and (_13446_, _03008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or (_03818_, _13446_, _13445_);
  and (_13447_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_13448_, _12558_, _23982_);
  or (_03820_, _13448_, _13447_);
  and (_13449_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and (_13450_, _13434_, _23755_);
  or (_27028_, _13450_, _13449_);
  and (_13451_, _12560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_13452_, _12558_, _23755_);
  or (_03835_, _13452_, _13451_);
  and (_13453_, _23864_, _23791_);
  and (_13454_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_27083_, _13454_, _13453_);
  and (_13455_, _23838_, _23601_);
  and (_13456_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or (_03842_, _13456_, _13455_);
  and (_13457_, _23864_, _23635_);
  and (_13458_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_03845_, _13458_, _13457_);
  and (_13459_, _23982_, _23864_);
  and (_13460_, _23866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_03851_, _13460_, _13459_);
  and (_13461_, _02225_, _23589_);
  and (_13462_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_03856_, _13462_, _13461_);
  and (_13463_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_13464_, _12549_, _23791_);
  or (_03870_, _13464_, _13463_);
  and (_13465_, _02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and (_13466_, _02762_, _23589_);
  or (_03873_, _13466_, _13465_);
  and (_13467_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_13468_, _12549_, _23838_);
  or (_03904_, _13468_, _13467_);
  and (_13469_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and (_13470_, _02233_, _23982_);
  or (_03906_, _13470_, _13469_);
  and (_13471_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_13472_, _12549_, _23982_);
  or (_03913_, _13472_, _13471_);
  and (_13473_, _02018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_13474_, _02017_, _23635_);
  or (_27064_, _13474_, _13473_);
  and (_13475_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_13476_, _12549_, _23635_);
  or (_03926_, _13476_, _13475_);
  and (_13477_, _12550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_13478_, _12549_, _23589_);
  or (_27127_, _13478_, _13477_);
  and (_13479_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_13480_, _25619_, _23791_);
  or (_03933_, _13480_, _13479_);
  and (_13481_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_13482_, _12599_, _23791_);
  or (_03936_, _13482_, _13481_);
  and (_13483_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_13484_, _12599_, _23676_);
  or (_03948_, _13484_, _13483_);
  and (_13485_, _05322_, _24541_);
  and (_13486_, _13485_, _23589_);
  not (_13487_, _13485_);
  and (_13488_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_03953_, _13488_, _13486_);
  and (_13489_, _06044_, _23755_);
  and (_13490_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_03957_, _13490_, _13489_);
  and (_13491_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_13492_, _25619_, _23635_);
  or (_03959_, _13492_, _13491_);
  and (_13493_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and (_13494_, _12539_, _23676_);
  or (_03962_, _13494_, _13493_);
  and (_13495_, _25620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_13496_, _25619_, _23982_);
  or (_27065_, _13496_, _13495_);
  and (_13497_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  and (_13498_, _12539_, _23718_);
  or (_27128_, _13498_, _13497_);
  and (_13499_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  and (_13500_, _12539_, _23982_);
  or (_27129_, _13500_, _13499_);
  and (_13501_, _25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and (_13502_, _25464_, _23755_);
  or (_03970_, _13502_, _13501_);
  and (_13503_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and (_13504_, _25294_, _23718_);
  or (_03995_, _13504_, _13503_);
  and (_13505_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  and (_13506_, _12539_, _23635_);
  or (_03999_, _13506_, _13505_);
  and (_13507_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and (_13508_, _25294_, _23676_);
  or (_04008_, _13508_, _13507_);
  and (_13509_, _12540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  and (_13510_, _12539_, _23589_);
  or (_04021_, _13510_, _13509_);
  and (_13511_, _25295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and (_13512_, _25294_, _23635_);
  or (_04024_, _13512_, _13511_);
  and (_13513_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_13514_, _24559_, _23635_);
  or (_04029_, _13514_, _13513_);
  and (_13515_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and (_13516_, _12530_, _23676_);
  or (_04032_, _13516_, _13515_);
  nand (_13517_, _24363_, _22767_);
  or (_13518_, _22767_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_13519_, _13518_, _22761_);
  and (_26873_[6], _13519_, _13517_);
  and (_13520_, _24560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_13521_, _24559_, _23718_);
  or (_04038_, _13521_, _13520_);
  and (_13522_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and (_13523_, _12530_, _23718_);
  or (_04041_, _13523_, _13522_);
  and (_13524_, _04733_, _24117_);
  not (_13525_, _13524_);
  and (_13526_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_13527_, _13524_, _23589_);
  or (_04044_, _13527_, _13526_);
  and (_13528_, _24214_, _23676_);
  and (_13529_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or (_04047_, _13529_, _13528_);
  and (_13530_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and (_13531_, _12530_, _23838_);
  or (_04050_, _13531_, _13530_);
  and (_13532_, _24093_, _23676_);
  and (_13533_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_04053_, _13533_, _13532_);
  and (_13534_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_13535_, _13524_, _23755_);
  or (_04058_, _13535_, _13534_);
  nand (_13536_, _23927_, _23832_);
  and (_13537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor (_13538_, _13537_, _23921_);
  not (_13539_, _13538_);
  and (_13540_, _13539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_13541_, _24165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not (_13542_, _13537_);
  and (_13543_, _23940_, _23938_);
  and (_13544_, _13543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_13545_, _13543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_13546_, _13545_, _13544_);
  and (_13547_, _13546_, _13542_);
  nor (_13548_, _13547_, _13541_);
  nor (_13549_, _13548_, _23921_);
  or (_13550_, _13549_, _13540_);
  or (_13551_, _13550_, _23927_);
  and (_13552_, _13551_, _22761_);
  and (_04060_, _13552_, _13536_);
  and (_13553_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_13554_, _13524_, _23635_);
  or (_04063_, _13554_, _13553_);
  and (_13555_, _24214_, _23755_);
  and (_13556_, _24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or (_27076_, _13556_, _13555_);
  and (_13557_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  and (_13558_, _12530_, _23982_);
  or (_27131_, _13558_, _13557_);
  and (_13559_, _06009_, _23635_);
  and (_13560_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_04082_, _13560_, _13559_);
  and (_13561_, _24093_, _23755_);
  and (_13562_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_04084_, _13562_, _13561_);
  and (_13563_, _13539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_13564_, _23948_, _23943_);
  and (_13565_, _24148_, _13564_);
  and (_13566_, _23938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_13567_, _23938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_13568_, _13567_, _13566_);
  and (_13569_, _13568_, _13542_);
  nor (_13570_, _13569_, _13565_);
  nor (_13571_, _13570_, _23921_);
  or (_13572_, _13571_, _23927_);
  or (_13573_, _13572_, _13563_);
  nand (_13574_, _23927_, _23669_);
  and (_13575_, _13574_, _22761_);
  and (_04087_, _13575_, _13573_);
  and (_13576_, _24093_, _23838_);
  and (_13577_, _24095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_04090_, _13577_, _13576_);
  or (_13578_, _23928_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_13579_, _13578_, _22761_);
  and (_13580_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_13581_, _13580_, _23950_);
  nand (_13582_, _13581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_13583_, _13581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_13584_, _13583_, _13582_);
  nor (_13585_, _13584_, _23921_);
  and (_13586_, _23921_, _24763_);
  or (_13587_, _13586_, _13585_);
  or (_13588_, _13587_, _23927_);
  and (_04094_, _13588_, _13579_);
  or (_13589_, _02962_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_13590_, _13589_, _02981_);
  and (_13591_, _13590_, _02993_);
  nor (_13592_, _02991_, _26569_);
  or (_13593_, _13592_, rst);
  or (_26872_[0], _13593_, _13591_);
  and (_13594_, _24089_, _23982_);
  and (_13595_, _24091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_04099_, _13595_, _13594_);
  and (_13596_, _12531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  and (_13597_, _12530_, _23635_);
  or (_04102_, _13597_, _13596_);
  and (_13598_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  and (_13599_, _12524_, _23791_);
  or (_27135_, _13599_, _13598_);
  nand (_13600_, _23994_, _23832_);
  nor (_13601_, _24048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_13602_, _24048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_13603_, _13602_, _13601_);
  and (_13604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_13605_, _13604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_13606_, _13605_, _24050_);
  and (_13607_, _13606_, _23997_);
  and (_13608_, _13607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_13609_, _13608_, _13603_);
  nor (_13610_, _13609_, _23988_);
  and (_13611_, _23988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_13612_, _13611_, _13610_);
  or (_13613_, _13612_, _23994_);
  and (_13614_, _13613_, _22761_);
  and (_04110_, _13614_, _13600_);
  and (_13615_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and (_13616_, _12524_, _23718_);
  or (_04113_, _13616_, _13615_);
  and (_13617_, _07101_, _23676_);
  and (_13618_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or (_04117_, _13618_, _13617_);
  and (_13619_, _23644_, _23635_);
  and (_13620_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_04120_, _13620_, _13619_);
  and (_13621_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  and (_13622_, _12524_, _23982_);
  or (_04125_, _13622_, _13621_);
  and (_13623_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  and (_13624_, _13434_, _23718_);
  or (_04127_, _13624_, _13623_);
  not (_13625_, _23988_);
  or (_13626_, _13625_, _23709_);
  and (_13627_, _24026_, _24000_);
  or (_13628_, _13627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_13629_, _13606_, _24001_);
  not (_13630_, _13629_);
  and (_13631_, _13630_, _23998_);
  and (_13632_, _13631_, _13628_);
  not (_13633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_13634_, _24050_, _24000_);
  nand (_13635_, _13634_, _13633_);
  and (_13636_, _24050_, _24001_);
  nor (_13637_, _13636_, _24054_);
  and (_13638_, _13637_, _13635_);
  and (_13639_, _24039_, _24000_);
  and (_13640_, _13639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor (_13641_, _13640_, _13633_);
  and (_13642_, _13640_, _13633_);
  or (_13643_, _13642_, _13641_);
  and (_13644_, _13643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_13645_, _13644_, _13638_);
  or (_13646_, _13645_, _13632_);
  or (_13647_, _13646_, _23988_);
  and (_13648_, _13647_, _23995_);
  and (_13649_, _13648_, _13626_);
  and (_13650_, _23994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_13651_, _13650_, _13649_);
  and (_04133_, _13651_, _22761_);
  or (_13652_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_13653_, _13652_, _22761_);
  not (_13654_, _23889_);
  or (_13655_, _13654_, _23709_);
  and (_04135_, _13655_, _13653_);
  and (_13656_, _07101_, _23718_);
  and (_13657_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or (_04137_, _13657_, _13656_);
  and (_13658_, _02225_, _23791_);
  and (_13659_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_27088_, _13659_, _13658_);
  and (_13660_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  and (_13661_, _12524_, _23635_);
  or (_04144_, _13661_, _13660_);
  and (_13662_, _12525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  and (_13663_, _12524_, _23589_);
  or (_04164_, _13663_, _13662_);
  and (_13664_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_13665_, _12512_, _23676_);
  or (_27136_, _13665_, _13664_);
  and (_13666_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and (_13667_, _13434_, _23791_);
  or (_04173_, _13667_, _13666_);
  and (_13668_, _24567_, _23589_);
  and (_13669_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or (_04176_, _13669_, _13668_);
  and (_13670_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and (_13671_, _13434_, _23676_);
  or (_04185_, _13671_, _13670_);
  and (_13672_, _24769_, _23755_);
  and (_13673_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or (_04189_, _13673_, _13672_);
  and (_13674_, _24769_, _23838_);
  and (_13675_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or (_04192_, _13675_, _13674_);
  and (_13676_, _24597_, _23982_);
  and (_13677_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or (_04198_, _13677_, _13676_);
  and (_13678_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_13679_, _12512_, _23791_);
  or (_04201_, _13679_, _13678_);
  and (_13680_, _24597_, _23718_);
  and (_13681_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or (_04209_, _13681_, _13680_);
  and (_13682_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_13683_, _12512_, _23838_);
  or (_27137_, _13683_, _13682_);
  and (_13684_, _25301_, _23718_);
  and (_13685_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_04213_, _13685_, _13684_);
  and (_13686_, _24597_, _23589_);
  and (_13687_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or (_04218_, _13687_, _13686_);
  and (_13688_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_13689_, _12512_, _23635_);
  or (_04221_, _13689_, _13688_);
  and (_13690_, _24583_, _24541_);
  and (_13691_, _13690_, _23676_);
  not (_13692_, _13690_);
  and (_13693_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_04225_, _13693_, _13691_);
  and (_13694_, _25301_, _23589_);
  and (_13695_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_04233_, _13695_, _13694_);
  and (_13696_, _24583_, _24117_);
  and (_13697_, _13696_, _23589_);
  not (_13698_, _13696_);
  and (_13699_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or (_04236_, _13699_, _13697_);
  and (_13700_, _12513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_13701_, _12512_, _23755_);
  or (_04244_, _13701_, _13700_);
  and (_13702_, _02444_, _23635_);
  and (_13703_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_27092_, _13703_, _13702_);
  and (_13704_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_13705_, _12500_, _23676_);
  or (_04249_, _13705_, _13704_);
  and (_13706_, _23849_, _23643_);
  and (_13707_, _13706_, _23676_);
  not (_13708_, _13706_);
  and (_13709_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or (_27097_, _13709_, _13707_);
  and (_13710_, _02436_, _23635_);
  and (_13711_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or (_27094_, _13711_, _13710_);
  and (_13712_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_13713_, _13524_, _23676_);
  or (_04275_, _13713_, _13712_);
  and (_13714_, _13706_, _23589_);
  and (_13715_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or (_04281_, _13715_, _13714_);
  and (_13716_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_13717_, _12500_, _23791_);
  or (_04283_, _13717_, _13716_);
  and (_13718_, _04733_, _23641_);
  not (_13719_, _13718_);
  and (_13720_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and (_13721_, _13718_, _23589_);
  or (_04286_, _13721_, _13720_);
  and (_13722_, _13706_, _23982_);
  and (_13723_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or (_04288_, _13723_, _13722_);
  and (_13724_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_13725_, _12500_, _23982_);
  or (_04292_, _13725_, _13724_);
  and (_13726_, _13690_, _23635_);
  and (_13727_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_04298_, _13727_, _13726_);
  and (_13728_, _06009_, _23982_);
  and (_13729_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_04301_, _13729_, _13728_);
  and (_13730_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  and (_13731_, _02840_, _23838_);
  or (_27099_, _13731_, _13730_);
  and (_13732_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_13733_, _12500_, _23635_);
  or (_04307_, _13733_, _13732_);
  and (_13734_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  and (_13735_, _02840_, _23791_);
  or (_04311_, _13735_, _13734_);
  and (_13736_, _24583_, _23854_);
  and (_13737_, _13736_, _23791_);
  not (_13738_, _13736_);
  and (_13739_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_04317_, _13739_, _13737_);
  or (_13740_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_13741_, _13740_, _22761_);
  nand (_13742_, _23889_, _23585_);
  and (_04320_, _13742_, _13741_);
  and (_13743_, _12501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_13744_, _12500_, _23589_);
  or (_04322_, _13744_, _13743_);
  and (_13745_, _13736_, _23838_);
  and (_13747_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_04324_, _13747_, _13745_);
  and (_13748_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_13749_, _09519_, _23676_);
  or (_04328_, _13749_, _13748_);
  and (_13750_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and (_13751_, _02840_, _23589_);
  or (_04331_, _13751_, _13750_);
  and (_13752_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and (_13753_, _12492_, _23676_);
  or (_04333_, _13753_, _13752_);
  and (_13754_, _13690_, _23838_);
  and (_13755_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_27189_, _13755_, _13754_);
  and (_13756_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  and (_13757_, _12492_, _23718_);
  or (_04346_, _13757_, _13756_);
  and (_13758_, _13690_, _23718_);
  and (_13759_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_27188_, _13759_, _13758_);
  and (_13760_, _23652_, _23589_);
  and (_13761_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_04354_, _13761_, _13760_);
  and (_13762_, _13690_, _23791_);
  and (_13763_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_27187_, _13763_, _13762_);
  and (_13764_, _24615_, _23594_);
  not (_13765_, _13764_);
  and (_13766_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  and (_13767_, _13764_, _23718_);
  or (_04373_, _13767_, _13766_);
  and (_13768_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  and (_13769_, _12492_, _23838_);
  or (_04377_, _13769_, _13768_);
  and (_13770_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_13771_, _13524_, _23838_);
  or (_04380_, _13771_, _13770_);
  and (_13772_, _13696_, _23676_);
  and (_13773_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or (_04389_, _13773_, _13772_);
  and (_13774_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  and (_13775_, _12492_, _23635_);
  or (_04392_, _13775_, _13774_);
  and (_13776_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_13777_, _13524_, _23718_);
  or (_04396_, _13777_, _13776_);
  and (_13778_, _13696_, _23791_);
  and (_13779_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or (_04399_, _13779_, _13778_);
  and (_13780_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  and (_13782_, _13764_, _23635_);
  or (_27106_, _13782_, _13780_);
  and (_13783_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_13784_, _13524_, _23791_);
  or (_27027_, _13784_, _13783_);
  and (_13785_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  and (_13786_, _09509_, _23755_);
  or (_04404_, _13786_, _13785_);
  and (_13787_, _12493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  and (_13788_, _12492_, _23755_);
  or (_04412_, _13788_, _13787_);
  and (_13789_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  and (_13790_, _09509_, _23838_);
  or (_04417_, _13790_, _13789_);
  and (_13791_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and (_13792_, _12486_, _23676_);
  or (_04420_, _13792_, _13791_);
  and (_13793_, _03658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_13794_, _03657_, _23718_);
  or (_04431_, _13794_, _13793_);
  or (_13795_, _24409_, _02363_);
  or (_13796_, _22767_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_13797_, _13796_, _22761_);
  and (_26873_[0], _13797_, _13795_);
  and (_13798_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_13799_, _24616_, _23838_);
  or (_04438_, _13799_, _13798_);
  and (_13800_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  and (_13801_, _12486_, _23791_);
  or (_04441_, _13801_, _13800_);
  and (_13802_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and (_13803_, _24616_, _23676_);
  or (_04445_, _13803_, _13802_);
  and (_13804_, _13696_, _23838_);
  and (_13805_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or (_04462_, _13805_, _13804_);
  and (_13806_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  and (_13807_, _02450_, _23718_);
  or (_27110_, _13807_, _13806_);
  and (_13808_, _13696_, _23635_);
  and (_13809_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or (_27170_, _13809_, _13808_);
  and (_13810_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and (_13811_, _12486_, _23838_);
  or (_27139_, _13811_, _13810_);
  and (_13812_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  and (_13813_, _13718_, _23791_);
  or (_04471_, _13813_, _13812_);
  and (_13814_, _24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_13815_, _24616_, _23589_);
  or (_04475_, _13815_, _13814_);
  and (_13816_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and (_13817_, _12486_, _23635_);
  or (_04478_, _13817_, _13816_);
  and (_13818_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_13819_, _02858_, _23791_);
  or (_04482_, _13819_, _13818_);
  and (_13820_, _13696_, _23982_);
  and (_13821_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or (_04485_, _13821_, _13820_);
  and (_13822_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  and (_13823_, _13718_, _23676_);
  or (_04490_, _13823_, _13822_);
  and (_13824_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  and (_13825_, _02450_, _23755_);
  or (_04492_, _13825_, _13824_);
  and (_13826_, _24768_, _24615_);
  not (_13827_, _13826_);
  and (_13828_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and (_13829_, _13826_, _23676_);
  or (_04495_, _13829_, _13828_);
  and (_13830_, _12487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  and (_13831_, _12486_, _23589_);
  or (_04498_, _13831_, _13830_);
  and (_13832_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and (_13833_, _09168_, _23635_);
  or (_04503_, _13833_, _13832_);
  and (_13834_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_13835_, _12478_, _23676_);
  or (_04523_, _13835_, _13834_);
  and (_13836_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  and (_13837_, _13826_, _23982_);
  or (_27114_, _13837_, _13836_);
  and (_13838_, _24615_, _23797_);
  not (_13839_, _13838_);
  and (_13840_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  and (_13841_, _13838_, _23838_);
  or (_04531_, _13841_, _13840_);
  and (_13842_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_13843_, _12478_, _23791_);
  or (_04536_, _13843_, _13842_);
  and (_13844_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and (_13845_, _13838_, _23676_);
  or (_04540_, _13845_, _13844_);
  and (_13846_, _24583_, _23797_);
  and (_13847_, _13846_, _23589_);
  not (_13848_, _13846_);
  and (_13849_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or (_04543_, _13849_, _13847_);
  and (_13850_, _13736_, _23589_);
  and (_13851_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_04546_, _13851_, _13850_);
  and (_13852_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and (_13853_, _13718_, _23718_);
  or (_04548_, _13853_, _13852_);
  and (_13854_, _13736_, _23982_);
  and (_13855_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_04550_, _13855_, _13854_);
  and (_13856_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_13857_, _12478_, _23838_);
  or (_04553_, _13857_, _13856_);
  and (_13858_, _13736_, _23755_);
  and (_13859_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_04555_, _13859_, _13858_);
  and (_13860_, _02277_, _23718_);
  and (_13861_, _02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or (_27186_, _13861_, _13860_);
  and (_13862_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_13863_, _12478_, _23635_);
  or (_04567_, _13863_, _13862_);
  and (_13864_, _24583_, _23641_);
  and (_13865_, _13864_, _23755_);
  not (_13866_, _13864_);
  and (_13867_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_27152_, _13867_, _13865_);
  and (_13868_, _24622_, _23838_);
  and (_13869_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_04574_, _13869_, _13868_);
  and (_13870_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_13871_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_13872_, _13871_, _13870_);
  and (_13873_, _13872_, _05352_);
  and (_13874_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_13875_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_13876_, _13875_, _13874_);
  and (_13877_, _13876_, _09527_);
  or (_13878_, _13877_, _13873_);
  or (_13879_, _13878_, _09540_);
  and (_13880_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_13881_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_13882_, _13881_, _13880_);
  and (_13883_, _13882_, _05352_);
  and (_13884_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_13885_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_13886_, _13885_, _13884_);
  and (_13887_, _13886_, _09527_);
  or (_13888_, _13887_, _13883_);
  or (_13889_, _13888_, _05373_);
  and (_13890_, _13889_, _09566_);
  and (_13891_, _13890_, _13879_);
  or (_13892_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_13893_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_13894_, _13893_, _09527_);
  and (_13895_, _13894_, _13892_);
  or (_13896_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_13897_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_13898_, _13897_, _05352_);
  and (_13899_, _13898_, _13896_);
  or (_13900_, _13899_, _13895_);
  or (_13901_, _13900_, _09540_);
  or (_13903_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_13904_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_13905_, _13904_, _09527_);
  and (_13906_, _13905_, _13903_);
  or (_13907_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_13908_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_13909_, _13908_, _05352_);
  and (_13910_, _13909_, _13907_);
  or (_13911_, _13910_, _13906_);
  or (_13912_, _13911_, _05373_);
  and (_13913_, _13912_, _05379_);
  and (_13914_, _13913_, _13901_);
  or (_13915_, _13914_, _13891_);
  or (_13916_, _13915_, _05361_);
  and (_13917_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_13918_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_13919_, _13918_, _09527_);
  or (_13920_, _13919_, _13917_);
  and (_13921_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_13922_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_13923_, _13922_, _05352_);
  or (_13924_, _13923_, _13921_);
  and (_13925_, _13924_, _13920_);
  or (_13926_, _13925_, _09540_);
  and (_13927_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_13928_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_13929_, _13928_, _09527_);
  or (_13930_, _13929_, _13927_);
  and (_13931_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_13932_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_13933_, _13932_, _05352_);
  or (_13934_, _13933_, _13931_);
  and (_13935_, _13934_, _13930_);
  or (_13936_, _13935_, _05373_);
  and (_13937_, _13936_, _09566_);
  and (_13938_, _13937_, _13926_);
  or (_13939_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_13940_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_13941_, _13940_, _13939_);
  or (_13942_, _13941_, _05352_);
  or (_13943_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_13944_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_13945_, _13944_, _13943_);
  or (_13946_, _13945_, _09527_);
  and (_13947_, _13946_, _13942_);
  or (_13948_, _13947_, _09540_);
  or (_13949_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_13950_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and (_13951_, _13950_, _13949_);
  or (_13952_, _13951_, _05352_);
  or (_13953_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_13954_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_13955_, _13954_, _13953_);
  or (_13956_, _13955_, _09527_);
  and (_13957_, _13956_, _13952_);
  or (_13958_, _13957_, _05373_);
  and (_13959_, _13958_, _05379_);
  and (_13960_, _13959_, _13948_);
  or (_13961_, _13960_, _13938_);
  or (_13962_, _13961_, _09581_);
  and (_13963_, _13962_, _09682_);
  and (_13964_, _13963_, _13916_);
  and (_13965_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_13966_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_13967_, _13966_, _13965_);
  and (_13968_, _13967_, _09527_);
  and (_13969_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_13970_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_13971_, _13970_, _13969_);
  and (_13972_, _13971_, _05352_);
  or (_13973_, _13972_, _13968_);
  and (_13974_, _13973_, _05373_);
  and (_13975_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_13976_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_13977_, _13976_, _13975_);
  and (_13978_, _13977_, _09527_);
  and (_13979_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_13980_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_13981_, _13980_, _13979_);
  and (_13982_, _13981_, _05352_);
  or (_13983_, _13982_, _13978_);
  and (_13984_, _13983_, _09540_);
  or (_13985_, _13984_, _13974_);
  and (_13986_, _13985_, _09566_);
  or (_13987_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_13988_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_13989_, _13988_, _13987_);
  and (_13990_, _13989_, _09527_);
  or (_13991_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_13992_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_13993_, _13992_, _13991_);
  and (_13994_, _13993_, _05352_);
  or (_13995_, _13994_, _13990_);
  and (_13996_, _13995_, _05373_);
  or (_13997_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_13998_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_13999_, _13998_, _13997_);
  and (_14000_, _13999_, _09527_);
  or (_14001_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_14002_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_14003_, _14002_, _14001_);
  and (_14004_, _14003_, _05352_);
  or (_14005_, _14004_, _14000_);
  and (_14006_, _14005_, _09540_);
  or (_14007_, _14006_, _13996_);
  and (_14008_, _14007_, _05379_);
  or (_14009_, _14008_, _13986_);
  and (_14010_, _14009_, _09581_);
  and (_14011_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and (_14012_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_14013_, _14012_, _14011_);
  and (_14014_, _14013_, _09527_);
  and (_14015_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_14016_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_14017_, _14016_, _14015_);
  and (_14018_, _14017_, _05352_);
  or (_14019_, _14018_, _14014_);
  and (_14020_, _14019_, _05373_);
  and (_14021_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and (_14022_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_14023_, _14022_, _14021_);
  and (_14024_, _14023_, _09527_);
  and (_14025_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and (_14026_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_14027_, _14026_, _14025_);
  and (_14028_, _14027_, _05352_);
  or (_14029_, _14028_, _14024_);
  and (_14030_, _14029_, _09540_);
  or (_14031_, _14030_, _14020_);
  and (_14032_, _14031_, _09566_);
  or (_14033_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_14034_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and (_14035_, _14034_, _14033_);
  and (_14036_, _14035_, _09527_);
  or (_14037_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_14038_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_14039_, _14038_, _14037_);
  and (_14040_, _14039_, _05352_);
  or (_14041_, _14040_, _14036_);
  and (_14042_, _14041_, _05373_);
  or (_14043_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_14044_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and (_14045_, _14044_, _14043_);
  and (_14046_, _14045_, _09527_);
  or (_14047_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_14048_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_14049_, _14048_, _14047_);
  and (_14050_, _14049_, _05352_);
  or (_14051_, _14050_, _14046_);
  and (_14052_, _14051_, _09540_);
  or (_14053_, _14052_, _14042_);
  and (_14054_, _14053_, _05379_);
  or (_14055_, _14054_, _14032_);
  and (_14056_, _14055_, _05361_);
  or (_14057_, _14056_, _14010_);
  and (_14058_, _14057_, _05363_);
  or (_14059_, _14058_, _13964_);
  or (_14060_, _14059_, _05357_);
  and (_14061_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and (_14062_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_14063_, _14062_, _14061_);
  and (_14064_, _14063_, _09527_);
  and (_14065_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_14066_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_14067_, _14066_, _14065_);
  and (_14068_, _14067_, _05352_);
  or (_14069_, _14068_, _14064_);
  or (_14070_, _14069_, _09540_);
  and (_14071_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_14072_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_14073_, _14072_, _14071_);
  and (_14074_, _14073_, _09527_);
  and (_14075_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and (_14076_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_14077_, _14076_, _14075_);
  and (_14078_, _14077_, _05352_);
  or (_14079_, _14078_, _14074_);
  or (_14080_, _14079_, _05373_);
  and (_14081_, _14080_, _09566_);
  and (_14082_, _14081_, _14070_);
  or (_14083_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_14084_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_14085_, _14084_, _05352_);
  and (_14086_, _14085_, _14083_);
  or (_14087_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_14088_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_14089_, _14088_, _09527_);
  and (_14090_, _14089_, _14087_);
  or (_14091_, _14090_, _14086_);
  or (_14092_, _14091_, _09540_);
  or (_14093_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_14094_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_14095_, _14094_, _05352_);
  and (_14096_, _14095_, _14093_);
  or (_14097_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_14098_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_14099_, _14098_, _09527_);
  and (_14100_, _14099_, _14097_);
  or (_14101_, _14100_, _14096_);
  or (_14102_, _14101_, _05373_);
  and (_14103_, _14102_, _05379_);
  and (_14104_, _14103_, _14092_);
  or (_14105_, _14104_, _14082_);
  and (_14106_, _14105_, _09581_);
  and (_14107_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_14108_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_14109_, _14108_, _14107_);
  and (_14110_, _14109_, _09527_);
  and (_14111_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_14112_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_14113_, _14112_, _14111_);
  and (_14114_, _14113_, _05352_);
  or (_14115_, _14114_, _14110_);
  or (_14116_, _14115_, _09540_);
  and (_14117_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_14118_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_14119_, _14118_, _14117_);
  and (_14120_, _14119_, _09527_);
  and (_14121_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_14122_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_14123_, _14122_, _14121_);
  and (_14124_, _14123_, _05352_);
  or (_14125_, _14124_, _14120_);
  or (_14126_, _14125_, _05373_);
  and (_14127_, _14126_, _09566_);
  and (_14128_, _14127_, _14116_);
  or (_14129_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_14130_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_14131_, _14130_, _14129_);
  and (_14132_, _14131_, _09527_);
  or (_14133_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_14134_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_14135_, _14134_, _14133_);
  and (_14136_, _14135_, _05352_);
  or (_14137_, _14136_, _14132_);
  or (_14138_, _14137_, _09540_);
  or (_14139_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_14140_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_14141_, _14140_, _14139_);
  and (_14142_, _14141_, _09527_);
  or (_14143_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_14144_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_14145_, _14144_, _14143_);
  and (_14146_, _14145_, _05352_);
  or (_14147_, _14146_, _14142_);
  or (_14148_, _14147_, _05373_);
  and (_14149_, _14148_, _05379_);
  and (_14150_, _14149_, _14138_);
  or (_14151_, _14150_, _14128_);
  and (_14152_, _14151_, _05361_);
  or (_14153_, _14152_, _14106_);
  and (_14154_, _14153_, _09682_);
  or (_14155_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_14156_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_14157_, _14156_, _14155_);
  and (_14158_, _14157_, _09527_);
  or (_14159_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_14160_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and (_14161_, _14160_, _14159_);
  and (_14162_, _14161_, _05352_);
  or (_14163_, _14162_, _14158_);
  and (_14164_, _14163_, _09540_);
  or (_14165_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_14166_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_14167_, _14166_, _14165_);
  and (_14168_, _14167_, _09527_);
  or (_14169_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_14170_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_14171_, _14170_, _14169_);
  and (_14172_, _14171_, _05352_);
  or (_14173_, _14172_, _14168_);
  and (_14174_, _14173_, _05373_);
  or (_14175_, _14174_, _14164_);
  and (_14176_, _14175_, _05379_);
  and (_14177_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_14178_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_14179_, _14178_, _14177_);
  and (_14180_, _14179_, _09527_);
  and (_14181_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_14182_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_14183_, _14182_, _14181_);
  and (_14184_, _14183_, _05352_);
  or (_14185_, _14184_, _14180_);
  and (_14186_, _14185_, _09540_);
  and (_14187_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_14188_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_14189_, _14188_, _14187_);
  and (_14190_, _14189_, _09527_);
  and (_14191_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and (_14192_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_14193_, _14192_, _14191_);
  and (_14194_, _14193_, _05352_);
  or (_14195_, _14194_, _14190_);
  and (_14196_, _14195_, _05373_);
  or (_14197_, _14196_, _14186_);
  and (_14198_, _14197_, _09566_);
  or (_14199_, _14198_, _14176_);
  and (_14200_, _14199_, _05361_);
  or (_14201_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_14202_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and (_14203_, _14202_, _05352_);
  and (_14204_, _14203_, _14201_);
  or (_14205_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_14206_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_14207_, _14206_, _09527_);
  and (_14208_, _14207_, _14205_);
  or (_14209_, _14208_, _14204_);
  and (_14210_, _14209_, _09540_);
  or (_14211_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_14212_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and (_14213_, _14212_, _05352_);
  and (_14214_, _14213_, _14211_);
  or (_14215_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_14216_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and (_14217_, _14216_, _09527_);
  and (_14218_, _14217_, _14215_);
  or (_14219_, _14218_, _14214_);
  and (_14220_, _14219_, _05373_);
  or (_14221_, _14220_, _14210_);
  and (_14222_, _14221_, _05379_);
  and (_14223_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_14224_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_14225_, _14224_, _14223_);
  and (_14226_, _14225_, _09527_);
  and (_14227_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_14228_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_14229_, _14228_, _14227_);
  and (_14230_, _14229_, _05352_);
  or (_14231_, _14230_, _14226_);
  and (_14232_, _14231_, _09540_);
  and (_14233_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_14234_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_14235_, _14234_, _14233_);
  and (_14236_, _14235_, _09527_);
  and (_14237_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_14238_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_14239_, _14238_, _14237_);
  and (_14240_, _14239_, _05352_);
  or (_14241_, _14240_, _14236_);
  and (_14242_, _14241_, _05373_);
  or (_14243_, _14242_, _14232_);
  and (_14244_, _14243_, _09566_);
  or (_14245_, _14244_, _14222_);
  and (_14246_, _14245_, _09581_);
  or (_14247_, _14246_, _14200_);
  and (_14248_, _14247_, _05363_);
  or (_14249_, _14248_, _14154_);
  or (_14250_, _14249_, _09739_);
  and (_14251_, _14250_, _14060_);
  or (_14252_, _14251_, _26838_);
  and (_14253_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_14254_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_14255_, _14254_, _14253_);
  and (_14256_, _14255_, _09527_);
  and (_14257_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_14258_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_14259_, _14258_, _14257_);
  and (_14260_, _14259_, _05352_);
  or (_14261_, _14260_, _14256_);
  or (_14262_, _14261_, _09540_);
  and (_14263_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_14264_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_14265_, _14264_, _14263_);
  and (_14266_, _14265_, _09527_);
  and (_14267_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_14268_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_14269_, _14268_, _14267_);
  and (_14270_, _14269_, _05352_);
  or (_14271_, _14270_, _14266_);
  or (_14272_, _14271_, _05373_);
  and (_14273_, _14272_, _09566_);
  and (_14274_, _14273_, _14262_);
  or (_14275_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_14276_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_14277_, _14276_, _14275_);
  and (_14278_, _14277_, _09527_);
  or (_14279_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_14280_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_14281_, _14280_, _14279_);
  and (_14282_, _14281_, _05352_);
  or (_14283_, _14282_, _14278_);
  or (_14284_, _14283_, _09540_);
  or (_14285_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_14286_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_14287_, _14286_, _14285_);
  and (_14288_, _14287_, _09527_);
  or (_14289_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_14290_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_14291_, _14290_, _14289_);
  and (_14292_, _14291_, _05352_);
  or (_14293_, _14292_, _14288_);
  or (_14294_, _14293_, _05373_);
  and (_14295_, _14294_, _05379_);
  and (_14296_, _14295_, _14284_);
  or (_14297_, _14296_, _14274_);
  and (_14298_, _14297_, _05361_);
  and (_14299_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_14300_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_14301_, _14300_, _14299_);
  and (_14302_, _14301_, _09527_);
  and (_14303_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_14304_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_14305_, _14304_, _14303_);
  and (_14306_, _14305_, _05352_);
  or (_14307_, _14306_, _14302_);
  or (_14308_, _14307_, _09540_);
  and (_14309_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_14310_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_14311_, _14310_, _14309_);
  and (_14312_, _14311_, _09527_);
  and (_14313_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_14314_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_14315_, _14314_, _14313_);
  and (_14316_, _14315_, _05352_);
  or (_14317_, _14316_, _14312_);
  or (_14318_, _14317_, _05373_);
  and (_14319_, _14318_, _09566_);
  and (_14320_, _14319_, _14308_);
  or (_14321_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_14322_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_14323_, _14322_, _05352_);
  and (_14324_, _14323_, _14321_);
  or (_14325_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_14326_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_14327_, _14326_, _09527_);
  and (_14328_, _14327_, _14325_);
  or (_14329_, _14328_, _14324_);
  or (_14330_, _14329_, _09540_);
  or (_14331_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_14332_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_14333_, _14332_, _05352_);
  and (_14334_, _14333_, _14331_);
  or (_14335_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_14336_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_14337_, _14336_, _09527_);
  and (_14338_, _14337_, _14335_);
  or (_14339_, _14338_, _14334_);
  or (_14340_, _14339_, _05373_);
  and (_14341_, _14340_, _05379_);
  and (_14342_, _14341_, _14330_);
  or (_14344_, _14342_, _14320_);
  and (_14345_, _14344_, _09581_);
  or (_14346_, _14345_, _14298_);
  and (_14347_, _14346_, _09682_);
  and (_14348_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_14349_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_14350_, _14349_, _14348_);
  and (_14351_, _14350_, _09527_);
  and (_14352_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_14353_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_14354_, _14353_, _14352_);
  and (_14355_, _14354_, _05352_);
  or (_14356_, _14355_, _14351_);
  and (_14357_, _14356_, _05373_);
  and (_14358_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_14359_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_14360_, _14359_, _14358_);
  and (_14361_, _14360_, _09527_);
  and (_14362_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_14363_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_14364_, _14363_, _14362_);
  and (_14365_, _14364_, _05352_);
  or (_14366_, _14365_, _14361_);
  and (_14367_, _14366_, _09540_);
  or (_14368_, _14367_, _14357_);
  and (_14369_, _14368_, _09566_);
  or (_14370_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_14371_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_14372_, _14371_, _05352_);
  and (_14373_, _14372_, _14370_);
  or (_14375_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_14376_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and (_14377_, _14376_, _09527_);
  and (_14378_, _14377_, _14375_);
  or (_14379_, _14378_, _14373_);
  and (_14380_, _14379_, _05373_);
  or (_14381_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_14382_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and (_14383_, _14382_, _05352_);
  and (_14384_, _14383_, _14381_);
  or (_14385_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_14386_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_14387_, _14386_, _09527_);
  and (_14388_, _14387_, _14385_);
  or (_14389_, _14388_, _14384_);
  and (_14390_, _14389_, _09540_);
  or (_14391_, _14390_, _14380_);
  and (_14392_, _14391_, _05379_);
  or (_14393_, _14392_, _14369_);
  and (_14394_, _14393_, _09581_);
  and (_14395_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_14396_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_14397_, _14396_, _14395_);
  and (_14398_, _14397_, _09527_);
  and (_14399_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_14400_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_14401_, _14400_, _14399_);
  and (_14402_, _14401_, _05352_);
  or (_14403_, _14402_, _14398_);
  and (_14404_, _14403_, _05373_);
  and (_14405_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_14406_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_14407_, _14406_, _14405_);
  and (_14408_, _14407_, _09527_);
  and (_14409_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_14410_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_14411_, _14410_, _14409_);
  and (_14412_, _14411_, _05352_);
  or (_14413_, _14412_, _14408_);
  and (_14414_, _14413_, _09540_);
  or (_14415_, _14414_, _14404_);
  and (_14416_, _14415_, _09566_);
  or (_14417_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_14418_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_14419_, _14418_, _14417_);
  and (_14420_, _14419_, _09527_);
  or (_14421_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_14422_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_14423_, _14422_, _14421_);
  and (_14424_, _14423_, _05352_);
  or (_14425_, _14424_, _14420_);
  and (_14426_, _14425_, _05373_);
  or (_14427_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_14428_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_14429_, _14428_, _14427_);
  and (_14430_, _14429_, _09527_);
  or (_14431_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_14432_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_14433_, _14432_, _14431_);
  and (_14434_, _14433_, _05352_);
  or (_14435_, _14434_, _14430_);
  and (_14436_, _14435_, _09540_);
  or (_14437_, _14436_, _14426_);
  and (_14438_, _14437_, _05379_);
  or (_14439_, _14438_, _14416_);
  and (_14440_, _14439_, _05361_);
  or (_14441_, _14440_, _14394_);
  and (_14442_, _14441_, _05363_);
  or (_14443_, _14442_, _14347_);
  or (_14444_, _14443_, _05357_);
  and (_14445_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_14446_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_14447_, _14446_, _14445_);
  and (_14448_, _14447_, _09527_);
  and (_14449_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_14450_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_14451_, _14450_, _14449_);
  and (_14452_, _14451_, _05352_);
  or (_14453_, _14452_, _14448_);
  or (_14454_, _14453_, _09540_);
  and (_14455_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_14456_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_14457_, _14456_, _14455_);
  and (_14458_, _14457_, _09527_);
  and (_14459_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_14460_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_14461_, _14460_, _14459_);
  and (_14462_, _14461_, _05352_);
  or (_14463_, _14462_, _14458_);
  or (_14464_, _14463_, _05373_);
  and (_14465_, _14464_, _09566_);
  and (_14466_, _14465_, _14454_);
  or (_14467_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_14468_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_14469_, _14468_, _05352_);
  and (_14470_, _14469_, _14467_);
  or (_14471_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_14472_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_14473_, _14472_, _09527_);
  and (_14474_, _14473_, _14471_);
  or (_14475_, _14474_, _14470_);
  or (_14476_, _14475_, _09540_);
  or (_14477_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_14478_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_14479_, _14478_, _05352_);
  and (_14480_, _14479_, _14477_);
  or (_14481_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_14482_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_14483_, _14482_, _09527_);
  and (_14484_, _14483_, _14481_);
  or (_14485_, _14484_, _14480_);
  or (_14486_, _14485_, _05373_);
  and (_14487_, _14486_, _05379_);
  and (_14488_, _14487_, _14476_);
  or (_14489_, _14488_, _14466_);
  and (_14490_, _14489_, _09581_);
  and (_14491_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_14492_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_14493_, _14492_, _14491_);
  and (_14494_, _14493_, _09527_);
  and (_14496_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_14497_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_14498_, _14497_, _14496_);
  and (_14499_, _14498_, _05352_);
  or (_14500_, _14499_, _14494_);
  or (_14501_, _14500_, _09540_);
  and (_14502_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_14503_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_14504_, _14503_, _14502_);
  and (_14505_, _14504_, _09527_);
  and (_14506_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_14507_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_14508_, _14507_, _14506_);
  and (_14509_, _14508_, _05352_);
  or (_14510_, _14509_, _14505_);
  or (_14511_, _14510_, _05373_);
  and (_14512_, _14511_, _09566_);
  and (_14513_, _14512_, _14501_);
  or (_14514_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_14515_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_14516_, _14515_, _14514_);
  and (_14517_, _14516_, _09527_);
  or (_14518_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_14519_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_14520_, _14519_, _14518_);
  and (_14521_, _14520_, _05352_);
  or (_14522_, _14521_, _14517_);
  or (_14523_, _14522_, _09540_);
  or (_14524_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_14525_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_14526_, _14525_, _14524_);
  and (_14527_, _14526_, _09527_);
  or (_14528_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_14529_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_14530_, _14529_, _14528_);
  and (_14531_, _14530_, _05352_);
  or (_14532_, _14531_, _14527_);
  or (_14533_, _14532_, _05373_);
  and (_14534_, _14533_, _05379_);
  and (_14535_, _14534_, _14523_);
  or (_14536_, _14535_, _14513_);
  and (_14537_, _14536_, _05361_);
  or (_14538_, _14537_, _14490_);
  and (_14539_, _14538_, _09682_);
  or (_14540_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_14541_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_14542_, _14541_, _14540_);
  and (_14543_, _14542_, _09527_);
  or (_14544_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_14545_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_14546_, _14545_, _14544_);
  and (_14547_, _14546_, _05352_);
  or (_14548_, _14547_, _14543_);
  and (_14549_, _14548_, _09540_);
  or (_14550_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_14551_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_14552_, _14551_, _14550_);
  and (_14553_, _14552_, _09527_);
  or (_14554_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_14555_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_14556_, _14555_, _14554_);
  and (_14557_, _14556_, _05352_);
  or (_14558_, _14557_, _14553_);
  and (_14559_, _14558_, _05373_);
  or (_14560_, _14559_, _14549_);
  and (_14561_, _14560_, _05379_);
  and (_14562_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_14563_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_14564_, _14563_, _14562_);
  and (_14565_, _14564_, _09527_);
  and (_14566_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_14567_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_14568_, _14567_, _14566_);
  and (_14569_, _14568_, _05352_);
  or (_14570_, _14569_, _14565_);
  and (_14571_, _14570_, _09540_);
  and (_14572_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_14573_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_14574_, _14573_, _14572_);
  and (_14575_, _14574_, _09527_);
  and (_14576_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_14577_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_14578_, _14577_, _14576_);
  and (_14579_, _14578_, _05352_);
  or (_14580_, _14579_, _14575_);
  and (_14581_, _14580_, _05373_);
  or (_14582_, _14581_, _14571_);
  and (_14583_, _14582_, _09566_);
  or (_14584_, _14583_, _14561_);
  and (_14585_, _14584_, _05361_);
  or (_14586_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_14587_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_14588_, _14587_, _05352_);
  and (_14589_, _14588_, _14586_);
  or (_14590_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_14591_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_14592_, _14591_, _09527_);
  and (_14593_, _14592_, _14590_);
  or (_14594_, _14593_, _14589_);
  and (_14595_, _14594_, _09540_);
  or (_14597_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_14598_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_14599_, _14598_, _05352_);
  and (_14600_, _14599_, _14597_);
  or (_14601_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_14602_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_14603_, _14602_, _09527_);
  and (_14604_, _14603_, _14601_);
  or (_14605_, _14604_, _14600_);
  and (_14606_, _14605_, _05373_);
  or (_14607_, _14606_, _14595_);
  and (_14608_, _14607_, _05379_);
  and (_14609_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_14610_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_14611_, _14610_, _14609_);
  and (_14612_, _14611_, _09527_);
  and (_14613_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_14614_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_14615_, _14614_, _14613_);
  and (_14616_, _14615_, _05352_);
  or (_14617_, _14616_, _14612_);
  and (_14618_, _14617_, _09540_);
  and (_14619_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_14620_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_14621_, _14620_, _14619_);
  and (_14622_, _14621_, _09527_);
  and (_14623_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_14624_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_14625_, _14624_, _14623_);
  and (_14626_, _14625_, _05352_);
  or (_14627_, _14626_, _14622_);
  and (_14628_, _14627_, _05373_);
  or (_14629_, _14628_, _14618_);
  and (_14630_, _14629_, _09566_);
  or (_14631_, _14630_, _14608_);
  and (_14632_, _14631_, _09581_);
  or (_14633_, _14632_, _14585_);
  and (_14634_, _14633_, _05363_);
  or (_14635_, _14634_, _14539_);
  or (_14636_, _14635_, _09739_);
  and (_14637_, _14636_, _14444_);
  or (_14638_, _14637_, _04360_);
  and (_14639_, _14638_, _14252_);
  or (_14640_, _14639_, _05401_);
  or (_14641_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_14642_, _14641_, _22761_);
  and (_04575_, _14642_, _14640_);
  and (_14643_, _24622_, _23676_);
  and (_14644_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_04577_, _14644_, _14643_);
  and (_14646_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  and (_14647_, _13718_, _23982_);
  or (_04581_, _14647_, _14646_);
  and (_14648_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_14649_, _12478_, _23755_);
  or (_04586_, _14649_, _14648_);
  and (_14650_, _24622_, _23791_);
  and (_14651_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_04590_, _14651_, _14650_);
  and (_14652_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and (_14653_, _06040_, _23635_);
  or (_04594_, _14653_, _14652_);
  and (_14654_, _06009_, _23589_);
  and (_14655_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_27098_, _14655_, _14654_);
  and (_14656_, _06041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_14657_, _06040_, _23718_);
  or (_04600_, _14657_, _14656_);
  and (_14658_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and (_14659_, _13718_, _23838_);
  or (_27026_, _14659_, _14658_);
  and (_14660_, _12479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_14661_, _12478_, _23589_);
  or (_04605_, _14661_, _14660_);
  and (_14662_, _02877_, _23718_);
  and (_14663_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_04607_, _14663_, _14662_);
  and (_14664_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and (_14665_, _03641_, _23676_);
  or (_04610_, _14665_, _14664_);
  and (_14666_, _12505_, _23755_);
  and (_14667_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or (_04611_, _14667_, _14666_);
  and (_14668_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and (_14669_, _04599_, _23676_);
  or (_04616_, _14669_, _14668_);
  and (_14670_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_14671_, _09168_, _23982_);
  or (_04618_, _14671_, _14670_);
  and (_14672_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_14673_, _12474_, _23676_);
  or (_04620_, _14673_, _14672_);
  and (_14674_, _13846_, _23791_);
  and (_14675_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or (_27197_, _14675_, _14674_);
  and (_14676_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_14677_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_14678_, _14677_, _14676_);
  and (_14679_, _14678_, _05352_);
  and (_14680_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_14681_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_14682_, _14681_, _14680_);
  and (_14683_, _14682_, _09527_);
  or (_14684_, _14683_, _14679_);
  or (_14685_, _14684_, _09540_);
  and (_14686_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_14687_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_14688_, _14687_, _14686_);
  and (_14689_, _14688_, _05352_);
  and (_14690_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_14691_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_14692_, _14691_, _14690_);
  and (_14693_, _14692_, _09527_);
  or (_14694_, _14693_, _14689_);
  or (_14695_, _14694_, _05373_);
  and (_14696_, _14695_, _09566_);
  and (_14697_, _14696_, _14685_);
  or (_14698_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_14699_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_14700_, _14699_, _09527_);
  and (_14701_, _14700_, _14698_);
  or (_14702_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_14703_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_14704_, _14703_, _05352_);
  and (_14705_, _14704_, _14702_);
  or (_14706_, _14705_, _14701_);
  or (_14707_, _14706_, _09540_);
  or (_14708_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_14709_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_14710_, _14709_, _09527_);
  and (_14711_, _14710_, _14708_);
  or (_14712_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_14713_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_14714_, _14713_, _05352_);
  and (_14715_, _14714_, _14712_);
  or (_14716_, _14715_, _14711_);
  or (_14717_, _14716_, _05373_);
  and (_14718_, _14717_, _05379_);
  and (_14719_, _14718_, _14707_);
  or (_14720_, _14719_, _14697_);
  and (_14721_, _14720_, _09581_);
  and (_14722_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_14723_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_14724_, _14723_, _09527_);
  or (_14725_, _14724_, _14722_);
  and (_14726_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_14727_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_14728_, _14727_, _05352_);
  or (_14729_, _14728_, _14726_);
  and (_14730_, _14729_, _14725_);
  or (_14731_, _14730_, _09540_);
  and (_14732_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_14733_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_14734_, _14733_, _09527_);
  or (_14735_, _14734_, _14732_);
  and (_14736_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_14737_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_14738_, _14737_, _05352_);
  or (_14739_, _14738_, _14736_);
  and (_14740_, _14739_, _14735_);
  or (_14742_, _14740_, _05373_);
  and (_14743_, _14742_, _09566_);
  and (_14744_, _14743_, _14731_);
  or (_14745_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_14746_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_14747_, _14746_, _14745_);
  or (_14748_, _14747_, _05352_);
  or (_14749_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_14750_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_14751_, _14750_, _14749_);
  or (_14752_, _14751_, _09527_);
  and (_14753_, _14752_, _14748_);
  or (_14754_, _14753_, _09540_);
  or (_14755_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_14756_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_14757_, _14756_, _14755_);
  or (_14758_, _14757_, _05352_);
  or (_14759_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_14760_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_14761_, _14760_, _14759_);
  or (_14762_, _14761_, _09527_);
  and (_14763_, _14762_, _14758_);
  or (_14764_, _14763_, _05373_);
  and (_14765_, _14764_, _05379_);
  and (_14766_, _14765_, _14754_);
  or (_14767_, _14766_, _14744_);
  and (_14768_, _14767_, _05361_);
  or (_14769_, _14768_, _14721_);
  and (_14770_, _14769_, _09682_);
  and (_14771_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_14772_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_14773_, _14772_, _14771_);
  and (_14774_, _14773_, _09527_);
  and (_14775_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_14776_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_14777_, _14776_, _14775_);
  and (_14778_, _14777_, _05352_);
  or (_14779_, _14778_, _14774_);
  and (_14780_, _14779_, _05373_);
  and (_14781_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_14782_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_14783_, _14782_, _14781_);
  and (_14784_, _14783_, _09527_);
  and (_14785_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_14786_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_14787_, _14786_, _14785_);
  and (_14788_, _14787_, _05352_);
  or (_14789_, _14788_, _14784_);
  and (_14790_, _14789_, _09540_);
  or (_14791_, _14790_, _05379_);
  or (_14792_, _14791_, _14780_);
  or (_14793_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_14794_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_14795_, _14794_, _14793_);
  and (_14796_, _14795_, _09527_);
  or (_14797_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_14798_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_14799_, _14798_, _14797_);
  and (_14800_, _14799_, _05352_);
  or (_14801_, _14800_, _14796_);
  and (_14802_, _14801_, _05373_);
  or (_14803_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_14804_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_14805_, _14804_, _14803_);
  and (_14806_, _14805_, _09527_);
  or (_14807_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_14808_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_14809_, _14808_, _14807_);
  and (_14810_, _14809_, _05352_);
  or (_14811_, _14810_, _14806_);
  and (_14812_, _14811_, _09540_);
  or (_14813_, _14812_, _09566_);
  or (_14814_, _14813_, _14802_);
  and (_14815_, _14814_, _14792_);
  or (_14816_, _14815_, _09581_);
  and (_14817_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and (_14818_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or (_14819_, _14818_, _14817_);
  and (_14820_, _14819_, _09527_);
  and (_14821_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and (_14822_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or (_14823_, _14822_, _14821_);
  and (_14824_, _14823_, _05352_);
  or (_14825_, _14824_, _14820_);
  and (_14826_, _14825_, _05373_);
  and (_14827_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and (_14828_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or (_14829_, _14828_, _14827_);
  and (_14830_, _14829_, _09527_);
  and (_14831_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and (_14832_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or (_14833_, _14832_, _14831_);
  and (_14834_, _14833_, _05352_);
  or (_14835_, _14834_, _14830_);
  and (_14836_, _14835_, _09540_);
  or (_14837_, _14836_, _05379_);
  or (_14838_, _14837_, _14826_);
  or (_14839_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or (_14840_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  and (_14841_, _14840_, _14839_);
  and (_14842_, _14841_, _09527_);
  or (_14843_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or (_14844_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and (_14845_, _14844_, _14843_);
  and (_14846_, _14845_, _05352_);
  or (_14847_, _14846_, _14842_);
  and (_14848_, _14847_, _05373_);
  or (_14849_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or (_14850_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and (_14851_, _14850_, _14849_);
  and (_14852_, _14851_, _09527_);
  or (_14853_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or (_14854_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and (_14855_, _14854_, _14853_);
  and (_14856_, _14855_, _05352_);
  or (_14857_, _14856_, _14852_);
  and (_14858_, _14857_, _09540_);
  or (_14859_, _14858_, _09566_);
  or (_14860_, _14859_, _14848_);
  and (_14861_, _14860_, _14838_);
  or (_14862_, _14861_, _05361_);
  and (_14863_, _14862_, _05363_);
  and (_14864_, _14863_, _14816_);
  or (_14865_, _14864_, _14770_);
  or (_14866_, _14865_, _05357_);
  and (_14867_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_14868_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_14869_, _14868_, _14867_);
  and (_14870_, _14869_, _09527_);
  and (_14871_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_14872_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_14873_, _14872_, _14871_);
  and (_14874_, _14873_, _05352_);
  or (_14875_, _14874_, _14870_);
  and (_14876_, _14875_, _09540_);
  and (_14877_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_14878_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_14879_, _14878_, _14877_);
  and (_14880_, _14879_, _09527_);
  and (_14881_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_14882_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_14883_, _14882_, _14881_);
  and (_14884_, _14883_, _05352_);
  or (_14885_, _14884_, _14880_);
  and (_14886_, _14885_, _05373_);
  or (_14887_, _14886_, _14876_);
  and (_14888_, _14887_, _09566_);
  or (_14889_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_14890_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_14891_, _14890_, _05352_);
  and (_14892_, _14891_, _14889_);
  or (_14893_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_14894_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_14895_, _14894_, _09527_);
  and (_14896_, _14895_, _14893_);
  or (_14897_, _14896_, _14892_);
  and (_14898_, _14897_, _09540_);
  or (_14899_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_14900_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_14901_, _14900_, _05352_);
  and (_14902_, _14901_, _14899_);
  or (_14903_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_14904_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_14905_, _14904_, _09527_);
  and (_14906_, _14905_, _14903_);
  or (_14907_, _14906_, _14902_);
  and (_14908_, _14907_, _05373_);
  or (_14909_, _14908_, _14898_);
  and (_14910_, _14909_, _05379_);
  or (_14911_, _14910_, _14888_);
  or (_14912_, _14911_, _05361_);
  and (_14913_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_14914_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_14915_, _14914_, _14913_);
  and (_14916_, _14915_, _09527_);
  and (_14917_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_14918_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_14919_, _14918_, _14917_);
  and (_14920_, _14919_, _05352_);
  or (_14921_, _14920_, _14916_);
  and (_14922_, _14921_, _09540_);
  and (_14923_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_14924_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_14925_, _14924_, _14923_);
  and (_14926_, _14925_, _09527_);
  and (_14927_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_14928_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_14929_, _14928_, _14927_);
  and (_14930_, _14929_, _05352_);
  or (_14931_, _14930_, _14926_);
  and (_14932_, _14931_, _05373_);
  or (_14933_, _14932_, _14922_);
  and (_14934_, _14933_, _09566_);
  or (_14935_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_14936_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_14937_, _14936_, _14935_);
  and (_14938_, _14937_, _09527_);
  or (_14939_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_14940_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_14941_, _14940_, _14939_);
  and (_14942_, _14941_, _05352_);
  or (_14943_, _14942_, _14938_);
  and (_14944_, _14943_, _09540_);
  or (_14945_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_14946_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_14947_, _14946_, _14945_);
  and (_14948_, _14947_, _09527_);
  or (_14949_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_14950_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_14951_, _14950_, _14949_);
  and (_14952_, _14951_, _05352_);
  or (_14953_, _14952_, _14948_);
  and (_14954_, _14953_, _05373_);
  or (_14955_, _14954_, _14944_);
  and (_14956_, _14955_, _05379_);
  or (_14957_, _14956_, _14934_);
  or (_14958_, _14957_, _09581_);
  and (_14959_, _14958_, _05363_);
  and (_14960_, _14959_, _14912_);
  and (_14961_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_14962_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_14963_, _14962_, _14961_);
  and (_14964_, _14963_, _09527_);
  and (_14965_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_14966_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_14967_, _14966_, _14965_);
  and (_14968_, _14967_, _05352_);
  or (_14969_, _14968_, _14964_);
  or (_14970_, _14969_, _09540_);
  and (_14971_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_14972_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_14973_, _14972_, _14971_);
  and (_14974_, _14973_, _09527_);
  and (_14975_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_14976_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_14977_, _14976_, _14975_);
  and (_14978_, _14977_, _05352_);
  or (_14979_, _14978_, _14974_);
  or (_14980_, _14979_, _05373_);
  and (_14981_, _14980_, _09566_);
  and (_14982_, _14981_, _14970_);
  or (_14983_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_14984_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_14985_, _14984_, _05352_);
  and (_14986_, _14985_, _14983_);
  or (_14987_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_14988_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_14989_, _14988_, _09527_);
  and (_14990_, _14989_, _14987_);
  or (_14991_, _14990_, _14986_);
  or (_14992_, _14991_, _09540_);
  or (_14993_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_14994_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_14995_, _14994_, _05352_);
  and (_14996_, _14995_, _14993_);
  or (_14997_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_14998_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_14999_, _14998_, _09527_);
  and (_15000_, _14999_, _14997_);
  or (_15001_, _15000_, _14996_);
  or (_15002_, _15001_, _05373_);
  and (_15003_, _15002_, _05379_);
  and (_15004_, _15003_, _14992_);
  or (_15005_, _15004_, _14982_);
  or (_15006_, _15005_, _05361_);
  and (_15007_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_15008_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_15009_, _15008_, _15007_);
  and (_15010_, _15009_, _09527_);
  and (_15011_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_15012_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_15013_, _15012_, _15011_);
  and (_15014_, _15013_, _05352_);
  or (_15015_, _15014_, _15010_);
  or (_15016_, _15015_, _09540_);
  and (_15017_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_15018_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_15019_, _15018_, _15017_);
  and (_15020_, _15019_, _09527_);
  and (_15021_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_15022_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_15023_, _15022_, _15021_);
  and (_15024_, _15023_, _05352_);
  or (_15025_, _15024_, _15020_);
  or (_15026_, _15025_, _05373_);
  and (_15027_, _15026_, _09566_);
  and (_15028_, _15027_, _15016_);
  or (_15029_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_15030_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_15031_, _15030_, _15029_);
  and (_15032_, _15031_, _09527_);
  or (_15033_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_15034_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_15035_, _15034_, _15033_);
  and (_15036_, _15035_, _05352_);
  or (_15037_, _15036_, _15032_);
  or (_15038_, _15037_, _09540_);
  or (_15039_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_15040_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_15041_, _15040_, _15039_);
  and (_15042_, _15041_, _09527_);
  or (_15043_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_15044_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_15045_, _15044_, _15043_);
  and (_15046_, _15045_, _05352_);
  or (_15047_, _15046_, _15042_);
  or (_15048_, _15047_, _05373_);
  and (_15049_, _15048_, _05379_);
  and (_15050_, _15049_, _15038_);
  or (_15051_, _15050_, _15028_);
  or (_15052_, _15051_, _09581_);
  and (_15053_, _15052_, _09682_);
  and (_15054_, _15053_, _15006_);
  or (_15055_, _15054_, _14960_);
  or (_15056_, _15055_, _09739_);
  and (_15057_, _15056_, _26838_);
  and (_15058_, _15057_, _14866_);
  and (_15059_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_15060_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_15061_, _15060_, _15059_);
  and (_15062_, _15061_, _05352_);
  and (_15063_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_15064_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_15065_, _15064_, _15063_);
  and (_15066_, _15065_, _09527_);
  or (_15067_, _15066_, _15062_);
  or (_15068_, _15067_, _09540_);
  and (_15069_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_15070_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_15071_, _15070_, _15069_);
  and (_15072_, _15071_, _05352_);
  and (_15073_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_15074_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_15075_, _15074_, _15073_);
  and (_15076_, _15075_, _09527_);
  or (_15077_, _15076_, _15072_);
  or (_15078_, _15077_, _05373_);
  and (_15079_, _15078_, _09566_);
  and (_15080_, _15079_, _15068_);
  or (_15081_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_15082_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_15083_, _15082_, _09527_);
  and (_15084_, _15083_, _15081_);
  or (_15085_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_15086_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_15087_, _15086_, _05352_);
  and (_15088_, _15087_, _15085_);
  or (_15089_, _15088_, _15084_);
  or (_15090_, _15089_, _09540_);
  or (_15091_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_15092_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and (_15093_, _15092_, _09527_);
  and (_15094_, _15093_, _15091_);
  or (_15095_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_15096_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_15097_, _15096_, _05352_);
  and (_15098_, _15097_, _15095_);
  or (_15099_, _15098_, _15094_);
  or (_15100_, _15099_, _05373_);
  and (_15101_, _15100_, _05379_);
  and (_15102_, _15101_, _15090_);
  or (_15103_, _15102_, _15080_);
  and (_15104_, _15103_, _09581_);
  and (_15105_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_15106_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_15107_, _15106_, _09527_);
  or (_15108_, _15107_, _15105_);
  and (_15109_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_15110_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_15111_, _15110_, _05352_);
  or (_15112_, _15111_, _15109_);
  and (_15113_, _15112_, _15108_);
  or (_15114_, _15113_, _09540_);
  and (_15115_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_15116_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_15117_, _15116_, _09527_);
  or (_15118_, _15117_, _15115_);
  and (_15119_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_15120_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_15121_, _15120_, _05352_);
  or (_15122_, _15121_, _15119_);
  and (_15123_, _15122_, _15118_);
  or (_15124_, _15123_, _05373_);
  and (_15125_, _15124_, _09566_);
  and (_15126_, _15125_, _15114_);
  or (_15127_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_15128_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_15129_, _15128_, _15127_);
  or (_15130_, _15129_, _05352_);
  or (_15131_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_15132_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_15133_, _15132_, _15131_);
  or (_15134_, _15133_, _09527_);
  and (_15135_, _15134_, _15130_);
  or (_15136_, _15135_, _09540_);
  or (_15137_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_15138_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_15139_, _15138_, _15137_);
  or (_15140_, _15139_, _05352_);
  or (_15141_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_15142_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_15143_, _15142_, _15141_);
  or (_15144_, _15143_, _09527_);
  and (_15145_, _15144_, _15140_);
  or (_15146_, _15145_, _05373_);
  and (_15147_, _15146_, _05379_);
  and (_15148_, _15147_, _15136_);
  or (_15149_, _15148_, _15126_);
  and (_15150_, _15149_, _05361_);
  or (_15151_, _15150_, _15104_);
  and (_15152_, _15151_, _09682_);
  or (_15153_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_15154_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_15155_, _15154_, _15153_);
  and (_15156_, _15155_, _09527_);
  or (_15157_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_15158_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and (_15159_, _15158_, _15157_);
  and (_15160_, _15159_, _05352_);
  or (_15161_, _15160_, _15156_);
  and (_15162_, _15161_, _09540_);
  or (_15163_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_15164_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_15165_, _15164_, _15163_);
  and (_15166_, _15165_, _09527_);
  or (_15167_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_15168_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_15169_, _15168_, _15167_);
  and (_15170_, _15169_, _05352_);
  or (_15171_, _15170_, _15166_);
  and (_15172_, _15171_, _05373_);
  or (_15173_, _15172_, _15162_);
  and (_15174_, _15173_, _05379_);
  and (_15175_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_15176_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_15177_, _15176_, _15175_);
  and (_15178_, _15177_, _09527_);
  and (_15179_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_15180_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_15181_, _15180_, _15179_);
  and (_15182_, _15181_, _05352_);
  or (_15183_, _15182_, _15178_);
  and (_15184_, _15183_, _09540_);
  and (_15185_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_15186_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_15187_, _15186_, _15185_);
  and (_15188_, _15187_, _09527_);
  and (_15189_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_15190_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_15191_, _15190_, _15189_);
  and (_15192_, _15191_, _05352_);
  or (_15193_, _15192_, _15188_);
  and (_15194_, _15193_, _05373_);
  or (_15195_, _15194_, _15184_);
  and (_15196_, _15195_, _09566_);
  or (_15197_, _15196_, _15174_);
  and (_15198_, _15197_, _05361_);
  or (_15199_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or (_15200_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and (_15201_, _15200_, _15199_);
  and (_15202_, _15201_, _09527_);
  or (_15203_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_15204_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and (_15205_, _15204_, _15203_);
  and (_15206_, _15205_, _05352_);
  or (_15207_, _15206_, _15202_);
  and (_15208_, _15207_, _09540_);
  or (_15209_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or (_15210_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and (_15211_, _15210_, _15209_);
  and (_15212_, _15211_, _09527_);
  or (_15213_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_15214_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  and (_15215_, _15214_, _15213_);
  and (_15216_, _15215_, _05352_);
  or (_15217_, _15216_, _15212_);
  and (_15218_, _15217_, _05373_);
  or (_15219_, _15218_, _15208_);
  and (_15220_, _15219_, _05379_);
  and (_15221_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and (_15222_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or (_15223_, _15222_, _15221_);
  and (_15224_, _15223_, _09527_);
  and (_15225_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  and (_15226_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_15227_, _15226_, _15225_);
  and (_15228_, _15227_, _05352_);
  or (_15229_, _15228_, _15224_);
  and (_15230_, _15229_, _09540_);
  and (_15231_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and (_15232_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_15233_, _15232_, _15231_);
  and (_15234_, _15233_, _09527_);
  and (_15235_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and (_15236_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or (_15237_, _15236_, _15235_);
  and (_15238_, _15237_, _05352_);
  or (_15239_, _15238_, _15234_);
  and (_15240_, _15239_, _05373_);
  or (_15241_, _15240_, _15230_);
  and (_15242_, _15241_, _09566_);
  or (_15243_, _15242_, _15220_);
  and (_15244_, _15243_, _09581_);
  or (_15245_, _15244_, _15198_);
  and (_15246_, _15245_, _05363_);
  or (_15247_, _15246_, _15152_);
  or (_15248_, _15247_, _09739_);
  or (_15249_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_15250_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_15251_, _15250_, _15249_);
  and (_15252_, _15251_, _09527_);
  or (_15253_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_15254_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_15255_, _15254_, _15253_);
  and (_15256_, _15255_, _05352_);
  or (_15257_, _15256_, _15252_);
  and (_15258_, _15257_, _09540_);
  or (_15259_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_15260_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_15261_, _15260_, _15259_);
  and (_15262_, _15261_, _09527_);
  or (_15263_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_15264_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_15265_, _15264_, _15263_);
  and (_15266_, _15265_, _05352_);
  or (_15267_, _15266_, _15262_);
  and (_15268_, _15267_, _05373_);
  or (_15269_, _15268_, _15258_);
  and (_15270_, _15269_, _05379_);
  and (_15271_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_15272_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_15273_, _15272_, _15271_);
  and (_15274_, _15273_, _09527_);
  and (_15275_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_15276_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_15277_, _15276_, _15275_);
  and (_15278_, _15277_, _05352_);
  or (_15279_, _15278_, _15274_);
  and (_15280_, _15279_, _09540_);
  and (_15281_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_15282_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_15283_, _15282_, _15281_);
  and (_15284_, _15283_, _09527_);
  and (_15285_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and (_15286_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_15287_, _15286_, _15285_);
  and (_15288_, _15287_, _05352_);
  or (_15289_, _15288_, _15284_);
  and (_15290_, _15289_, _05373_);
  or (_15291_, _15290_, _15280_);
  and (_15292_, _15291_, _09566_);
  or (_15293_, _15292_, _15270_);
  and (_15294_, _15293_, _05361_);
  or (_15295_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_15296_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_15297_, _15296_, _05352_);
  and (_15298_, _15297_, _15295_);
  or (_15299_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_15300_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_15301_, _15300_, _09527_);
  and (_15302_, _15301_, _15299_);
  or (_15303_, _15302_, _15298_);
  and (_15304_, _15303_, _09540_);
  or (_15305_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_15306_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_15307_, _15306_, _05352_);
  and (_15308_, _15307_, _15305_);
  or (_15309_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_15310_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_15311_, _15310_, _09527_);
  and (_15312_, _15311_, _15309_);
  or (_15313_, _15312_, _15308_);
  and (_15314_, _15313_, _05373_);
  or (_15315_, _15314_, _15304_);
  and (_15316_, _15315_, _05379_);
  and (_15317_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_15318_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_15319_, _15318_, _15317_);
  and (_15320_, _15319_, _09527_);
  and (_15321_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_15322_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_15323_, _15322_, _15321_);
  and (_15324_, _15323_, _05352_);
  or (_15325_, _15324_, _15320_);
  and (_15326_, _15325_, _09540_);
  and (_15327_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_15328_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_15329_, _15328_, _15327_);
  and (_15330_, _15329_, _09527_);
  and (_15331_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_15332_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_15333_, _15332_, _15331_);
  and (_15334_, _15333_, _05352_);
  or (_15335_, _15334_, _15330_);
  and (_15336_, _15335_, _05373_);
  or (_15337_, _15336_, _15326_);
  and (_15338_, _15337_, _09566_);
  or (_15339_, _15338_, _15316_);
  and (_15340_, _15339_, _09581_);
  or (_15341_, _15340_, _15294_);
  and (_15342_, _15341_, _05363_);
  and (_15343_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_15344_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_15345_, _15344_, _15343_);
  and (_15346_, _15345_, _09527_);
  and (_15347_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_15348_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_15349_, _15348_, _15347_);
  and (_15350_, _15349_, _05352_);
  or (_15351_, _15350_, _15346_);
  or (_15352_, _15351_, _09540_);
  and (_15353_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_15354_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_15355_, _15354_, _15353_);
  and (_15356_, _15355_, _09527_);
  and (_15357_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_15358_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_15359_, _15358_, _15357_);
  and (_15360_, _15359_, _05352_);
  or (_15361_, _15360_, _15356_);
  or (_15362_, _15361_, _05373_);
  and (_15363_, _15362_, _09566_);
  and (_15364_, _15363_, _15352_);
  or (_15365_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_15366_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and (_15367_, _15366_, _05352_);
  and (_15368_, _15367_, _15365_);
  or (_15369_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_15370_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and (_15371_, _15370_, _09527_);
  and (_15372_, _15371_, _15369_);
  or (_15373_, _15372_, _15368_);
  or (_15374_, _15373_, _09540_);
  or (_15375_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_15376_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_15377_, _15376_, _05352_);
  and (_15378_, _15377_, _15375_);
  or (_15379_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_15380_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_15381_, _15380_, _09527_);
  and (_15382_, _15381_, _15379_);
  or (_15383_, _15382_, _15378_);
  or (_15384_, _15383_, _05373_);
  and (_15385_, _15384_, _05379_);
  and (_15386_, _15385_, _15374_);
  or (_15387_, _15386_, _15364_);
  and (_15388_, _15387_, _09581_);
  and (_15389_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_15390_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_15391_, _15390_, _15389_);
  and (_15392_, _15391_, _09527_);
  and (_15393_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_15394_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_15395_, _15394_, _15393_);
  and (_15396_, _15395_, _05352_);
  or (_15397_, _15396_, _15392_);
  or (_15398_, _15397_, _09540_);
  and (_15399_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_15400_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_15401_, _15400_, _15399_);
  and (_15402_, _15401_, _09527_);
  and (_15403_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_15404_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_15405_, _15404_, _15403_);
  and (_15406_, _15405_, _05352_);
  or (_15407_, _15406_, _15402_);
  or (_15408_, _15407_, _05373_);
  and (_15409_, _15408_, _09566_);
  and (_15410_, _15409_, _15398_);
  or (_15411_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_15412_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_15413_, _15412_, _15411_);
  and (_15414_, _15413_, _09527_);
  or (_15415_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_15416_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_15417_, _15416_, _15415_);
  and (_15418_, _15417_, _05352_);
  or (_15419_, _15418_, _15414_);
  or (_15420_, _15419_, _09540_);
  or (_15421_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_15422_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_15423_, _15422_, _15421_);
  and (_15424_, _15423_, _09527_);
  or (_15425_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_15426_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_15427_, _15426_, _15425_);
  and (_15428_, _15427_, _05352_);
  or (_15429_, _15428_, _15424_);
  or (_15430_, _15429_, _05373_);
  and (_15431_, _15430_, _05379_);
  and (_15432_, _15431_, _15420_);
  or (_15433_, _15432_, _15410_);
  and (_15434_, _15433_, _05361_);
  or (_15435_, _15434_, _15388_);
  and (_15436_, _15435_, _09682_);
  or (_15437_, _15436_, _15342_);
  or (_15438_, _15437_, _05357_);
  and (_15439_, _15438_, _04360_);
  and (_15440_, _15439_, _15248_);
  or (_15441_, _15440_, _15058_);
  or (_15442_, _15441_, _05401_);
  or (_15443_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_15444_, _15443_, _22761_);
  and (_04628_, _15444_, _15442_);
  and (_15445_, _12505_, _23635_);
  and (_15446_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or (_27264_, _15446_, _15445_);
  and (_15447_, _13846_, _23676_);
  and (_15448_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or (_04647_, _15448_, _15447_);
  or (_15449_, _23928_, _23709_);
  and (_15450_, _23939_, _23938_);
  nor (_15451_, _15450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_15452_, _15451_, _13543_);
  and (_15453_, _15452_, _13538_);
  and (_15454_, _13539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_15455_, _13580_, _23948_);
  and (_15456_, _15455_, _24148_);
  nand (_15457_, _15456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_15458_, _15457_, _23921_);
  or (_15459_, _15458_, _15454_);
  or (_15460_, _15459_, _15453_);
  or (_15461_, _15460_, _23927_);
  and (_15462_, _15461_, _22761_);
  and (_04648_, _15462_, _15449_);
  and (_15463_, _04733_, _23863_);
  not (_15464_, _15463_);
  and (_15465_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  and (_15466_, _15463_, _23838_);
  or (_04666_, _15466_, _15465_);
  and (_15467_, _13846_, _23635_);
  and (_15468_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or (_04669_, _15468_, _15467_);
  and (_15469_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_15470_, _09168_, _23838_);
  or (_04680_, _15470_, _15469_);
  and (_15471_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  and (_15472_, _15463_, _23718_);
  or (_04685_, _15472_, _15471_);
  and (_15473_, _13846_, _23982_);
  and (_15474_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or (_04691_, _15474_, _15473_);
  and (_15475_, _13846_, _23838_);
  and (_15476_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or (_04694_, _15476_, _15475_);
  and (_15477_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  and (_15478_, _15463_, _23791_);
  or (_04697_, _15478_, _15477_);
  and (_15479_, _24597_, _23791_);
  and (_15480_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or (_04716_, _15480_, _15479_);
  and (_15481_, _23842_, _23028_);
  and (_15482_, _15481_, _23635_);
  not (_15483_, _15481_);
  and (_15484_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or (_04721_, _15484_, _15482_);
  and (_15485_, _24768_, _24583_);
  and (_15486_, _15485_, _23838_);
  not (_15487_, _15485_);
  and (_15488_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or (_04723_, _15488_, _15486_);
  and (_15489_, _15485_, _23718_);
  and (_15490_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or (_04725_, _15490_, _15489_);
  and (_15491_, _15481_, _23982_);
  and (_15492_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or (_04729_, _15492_, _15491_);
  and (_15493_, _24597_, _23676_);
  and (_15494_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or (_04732_, _15494_, _15493_);
  and (_15495_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and (_15496_, _15463_, _23982_);
  or (_04738_, _15496_, _15495_);
  and (_15497_, _15485_, _23791_);
  and (_15498_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or (_04745_, _15498_, _15497_);
  and (_15499_, _15485_, _23676_);
  and (_15500_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or (_04748_, _15500_, _15499_);
  and (_15501_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  and (_15502_, _15463_, _23755_);
  or (_27023_, _15502_, _15501_);
  and (_15503_, _23649_, _23028_);
  and (_15504_, _15503_, _23755_);
  not (_15505_, _15503_);
  and (_15506_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_04755_, _15506_, _15504_);
  and (_15507_, _06264_, _23838_);
  and (_15508_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_04760_, _15508_, _15507_);
  and (_15509_, _15503_, _23635_);
  and (_15510_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_04762_, _15510_, _15509_);
  and (_15511_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and (_15512_, _15463_, _23635_);
  or (_04768_, _15512_, _15511_);
  and (_15513_, _15503_, _23982_);
  and (_15514_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_04770_, _15514_, _15513_);
  and (_15515_, _15485_, _23755_);
  and (_15516_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or (_04782_, _15516_, _15515_);
  and (_15517_, _15485_, _23635_);
  and (_15518_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or (_04784_, _15518_, _15517_);
  and (_15519_, _15485_, _23982_);
  and (_15520_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or (_04788_, _15520_, _15519_);
  and (_15521_, _07101_, _23791_);
  and (_15522_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or (_04791_, _15522_, _15521_);
  and (_15523_, _04733_, _24103_);
  not (_15524_, _15523_);
  and (_15525_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_15526_, _15523_, _23718_);
  or (_04806_, _15526_, _15525_);
  and (_15527_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_15528_, _15523_, _23982_);
  or (_04809_, _15528_, _15527_);
  and (_15529_, _13690_, _23589_);
  and (_15530_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_04821_, _15530_, _15529_);
  and (_15531_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_15532_, _15523_, _23838_);
  or (_27021_, _15532_, _15531_);
  and (_15533_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_15534_, _09168_, _23589_);
  or (_27117_, _15534_, _15533_);
  and (_15535_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_15536_, _09168_, _23755_);
  or (_04862_, _15536_, _15535_);
  and (_15537_, _24583_, _23863_);
  and (_15538_, _15537_, _23838_);
  not (_15539_, _15537_);
  and (_15540_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_04872_, _15540_, _15538_);
  and (_15541_, _15537_, _23718_);
  and (_15542_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_04877_, _15542_, _15541_);
  and (_15543_, _15537_, _23791_);
  and (_15544_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_04885_, _15544_, _15543_);
  and (_15545_, _02779_, _23635_);
  and (_15546_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_04891_, _15546_, _15545_);
  and (_15547_, _06009_, _23755_);
  and (_15548_, _06011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_04900_, _15548_, _15547_);
  and (_15549_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_15550_, _15523_, _23589_);
  or (_04903_, _15550_, _15549_);
  and (_15551_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_15552_, _15523_, _23755_);
  or (_04914_, _15552_, _15551_);
  and (_15553_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_15554_, _15523_, _23635_);
  or (_27022_, _15554_, _15553_);
  and (_15555_, _15537_, _23755_);
  and (_15556_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_04927_, _15556_, _15555_);
  and (_15557_, _15537_, _23635_);
  and (_15558_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_04934_, _15558_, _15557_);
  and (_15559_, _15537_, _23982_);
  and (_15560_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_04941_, _15560_, _15559_);
  and (_15561_, _23791_, _23601_);
  and (_15562_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or (_04943_, _15562_, _15561_);
  and (_15563_, _04733_, _23594_);
  not (_15564_, _15563_);
  and (_15565_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_15566_, _15563_, _23755_);
  or (_04982_, _15566_, _15565_);
  and (_15567_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_15568_, _15563_, _23635_);
  or (_04986_, _15568_, _15567_);
  and (_15569_, _24584_, _23635_);
  and (_15570_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or (_04991_, _15570_, _15569_);
  and (_15571_, _24584_, _23982_);
  and (_15572_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or (_04997_, _15572_, _15571_);
  and (_15573_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and (_15574_, _03205_, _23755_);
  or (_04999_, _15574_, _15573_);
  and (_15575_, _12505_, _23676_);
  and (_15576_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_05003_, _15576_, _15575_);
  and (_15577_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_15578_, _12474_, _23755_);
  or (_05015_, _15578_, _15577_);
  and (_15579_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_15580_, _12474_, _23635_);
  or (_27141_, _15580_, _15579_);
  and (_15581_, _03256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_15582_, _03255_, _23982_);
  or (_05024_, _15582_, _15581_);
  and (_15583_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_15584_, _12474_, _23589_);
  or (_05033_, _15584_, _15583_);
  and (_15585_, _24584_, _23589_);
  and (_15586_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_05036_, _15586_, _15585_);
  and (_15587_, _03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and (_15588_, _03184_, _23755_);
  or (_05041_, _15588_, _15587_);
  and (_15589_, _24584_, _23755_);
  and (_15590_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or (_05053_, _15590_, _15589_);
  and (_15591_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_15592_, _15523_, _23676_);
  or (_05071_, _15592_, _15591_);
  and (_15593_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_15594_, _15563_, _23589_);
  or (_05075_, _15594_, _15593_);
  and (_15595_, _03322_, _23676_);
  and (_15596_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_05086_, _15596_, _15595_);
  and (_15597_, _03322_, _23718_);
  and (_15598_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_05089_, _15598_, _15597_);
  and (_15599_, _13864_, _23718_);
  and (_15600_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_05094_, _15600_, _15599_);
  and (_15601_, _13864_, _23791_);
  and (_15602_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_05098_, _15602_, _15601_);
  and (_15603_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  and (_15604_, _03205_, _23791_);
  or (_05107_, _15604_, _15603_);
  and (_15605_, _13864_, _23676_);
  and (_15606_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_27150_, _15606_, _15605_);
  and (_15607_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and (_15608_, _04557_, _23676_);
  or (_05112_, _15608_, _15607_);
  and (_15609_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and (_15610_, _03205_, _23676_);
  or (_05114_, _15610_, _15609_);
  and (_15611_, _04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  and (_15612_, _04557_, _23982_);
  or (_05116_, _15612_, _15611_);
  and (_15613_, _03206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  and (_15614_, _03205_, _23718_);
  or (_05118_, _15614_, _15613_);
  and (_15615_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_15616_, _03314_, _23755_);
  or (_05121_, _15616_, _15615_);
  and (_15617_, _04733_, _23962_);
  not (_15618_, _15617_);
  and (_15619_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  and (_15620_, _15617_, _23589_);
  or (_05132_, _15620_, _15619_);
  and (_15621_, _15503_, _23589_);
  and (_15622_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_05136_, _15622_, _15621_);
  and (_15623_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  and (_15624_, _09509_, _23718_);
  or (_05139_, _15624_, _15623_);
  and (_15625_, _13864_, _23982_);
  and (_15626_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_05150_, _15626_, _15625_);
  and (_15627_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  and (_15628_, _15617_, _23755_);
  or (_27017_, _15628_, _15627_);
  and (_15629_, _13864_, _23838_);
  and (_15630_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_27151_, _15630_, _15629_);
  and (_15631_, _03322_, _23755_);
  and (_15632_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_05174_, _15632_, _15631_);
  and (_15633_, _13864_, _23589_);
  and (_15634_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_05192_, _15634_, _15633_);
  and (_15635_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_15636_, _15563_, _23718_);
  or (_05209_, _15636_, _15635_);
  and (_15637_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_15638_, _12474_, _23982_);
  or (_05224_, _15638_, _15637_);
  and (_15639_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and (_15640_, _04595_, _23589_);
  or (_05231_, _15640_, _15639_);
  nor (_15641_, _13566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_15642_, _15641_, _15450_);
  and (_15643_, _15642_, _13538_);
  and (_15644_, _13539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_15645_, _15644_, _15643_);
  nand (_15646_, _24165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_15647_, _15646_, _23921_);
  or (_15648_, _15647_, _23927_);
  or (_15649_, _15648_, _15645_);
  nand (_15650_, _23927_, _23784_);
  and (_15651_, _15650_, _22761_);
  and (_05233_, _15651_, _15649_);
  and (_15652_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  and (_15653_, _04599_, _23755_);
  or (_27122_, _15653_, _15652_);
  and (_15654_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_15655_, _12474_, _23718_);
  or (_27140_, _15655_, _15654_);
  and (_15656_, _04601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  and (_15657_, _04599_, _23838_);
  or (_05243_, _15657_, _15656_);
  and (_15658_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_15659_, _15563_, _23791_);
  or (_27018_, _15659_, _15658_);
  and (_15660_, _04596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_15661_, _04595_, _23982_);
  or (_05275_, _15661_, _15660_);
  and (_15662_, _12475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_15663_, _12474_, _23838_);
  or (_05277_, _15663_, _15662_);
  and (_15664_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and (_15665_, _13838_, _23589_);
  or (_05279_, _15665_, _15664_);
  and (_15666_, _02877_, _23982_);
  and (_15667_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_05285_, _15667_, _15666_);
  and (_15668_, _03322_, _23838_);
  and (_15669_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_05310_, _15669_, _15668_);
  and (_15670_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  and (_15671_, _13838_, _23755_);
  or (_05337_, _15671_, _15670_);
  and (_15672_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_15673_, _10517_, _23589_);
  or (_05340_, _15673_, _15672_);
  and (_15674_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_15675_, _10517_, _23982_);
  or (_27059_, _15675_, _15674_);
  and (_15676_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_15677_, _10517_, _23676_);
  or (_05366_, _15677_, _15676_);
  and (_15678_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  and (_15679_, _09523_, _23589_);
  or (_05370_, _15679_, _15678_);
  and (_15680_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and (_15681_, _09523_, _23635_);
  or (_05383_, _15681_, _15680_);
  and (_15682_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_15683_, _09481_, _23982_);
  or (_05406_, _15683_, _15682_);
  and (_15684_, _00301_, _25117_);
  and (_15685_, _15684_, _24713_);
  not (_15686_, _15685_);
  or (_15687_, _15686_, _00874_);
  or (_15688_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_15689_, _15688_, _23880_);
  and (_15690_, _15689_, _15687_);
  and (_15691_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_15692_, _15684_, _24671_);
  nand (_15693_, _15692_, _23522_);
  or (_15694_, _15692_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_15695_, _15694_, _24629_);
  and (_15696_, _15695_, _15693_);
  or (_15697_, _15696_, _15691_);
  or (_15698_, _15697_, _15690_);
  and (_05419_, _15698_, _22761_);
  and (_15699_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_15700_, _09481_, _23676_);
  or (_05422_, _15700_, _15699_);
  and (_15701_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_15702_, _08427_, _23635_);
  or (_05429_, _15702_, _15701_);
  and (_15703_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_15704_, _08427_, _23718_);
  or (_05432_, _15704_, _15703_);
  and (_15705_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and (_15706_, _06296_, _23589_);
  or (_27047_, _15706_, _15705_);
  and (_15707_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and (_15708_, _06296_, _23838_);
  or (_27044_, _15708_, _15707_);
  and (_15709_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_15710_, _06296_, _23676_);
  or (_05467_, _15710_, _15709_);
  and (_15711_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and (_15712_, _05439_, _23589_);
  or (_05472_, _15712_, _15711_);
  and (_15713_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and (_15714_, _05439_, _23635_);
  or (_05476_, _15714_, _15713_);
  and (_15715_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and (_15716_, _05439_, _23676_);
  or (_05491_, _15716_, _15715_);
  and (_15717_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_15718_, _05420_, _23755_);
  or (_05494_, _15718_, _15717_);
  and (_15719_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_15720_, _05420_, _23791_);
  or (_05506_, _15720_, _15719_);
  and (_15721_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and (_15722_, _05407_, _23755_);
  or (_05512_, _15722_, _15721_);
  and (_15723_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and (_15724_, _05407_, _23791_);
  or (_05516_, _15724_, _15723_);
  and (_15725_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  and (_15726_, _04810_, _23755_);
  or (_05520_, _15726_, _15725_);
  and (_15727_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  and (_15728_, _04810_, _23982_);
  or (_27036_, _15728_, _15727_);
  and (_15729_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and (_15730_, _04810_, _23676_);
  or (_05527_, _15730_, _15729_);
  and (_15731_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_15732_, _04792_, _23589_);
  or (_05531_, _15732_, _15731_);
  and (_15733_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_15734_, _04792_, _23635_);
  or (_05535_, _15734_, _15733_);
  and (_15735_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_15736_, _04792_, _23791_);
  or (_05540_, _15736_, _15735_);
  and (_15737_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_15738_, _04776_, _23755_);
  or (_05572_, _15738_, _15737_);
  and (_15739_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_15740_, _04756_, _23635_);
  or (_05579_, _15740_, _15739_);
  and (_15741_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_15742_, _04756_, _23718_);
  or (_05581_, _15742_, _15741_);
  and (_15743_, _03302_, _23838_);
  and (_15744_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  or (_05587_, _15744_, _15743_);
  and (_15745_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  and (_15746_, _09523_, _23791_);
  or (_27055_, _15746_, _15745_);
  and (_15747_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_15748_, _09481_, _23755_);
  or (_27054_, _15748_, _15747_);
  and (_15749_, _09482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_15750_, _09481_, _23718_);
  or (_27052_, _15750_, _15749_);
  and (_15751_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_15752_, _08427_, _23589_);
  or (_05629_, _15752_, _15751_);
  and (_15753_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  and (_15754_, _05439_, _23718_);
  or (_05652_, _15754_, _15753_);
  and (_15755_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_15756_, _05420_, _23838_);
  or (_05658_, _15756_, _15755_);
  and (_15757_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and (_15758_, _05407_, _23838_);
  or (_05664_, _15758_, _15757_);
  and (_15759_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and (_15760_, _15617_, _23791_);
  or (_05667_, _15760_, _15759_);
  and (_15761_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  and (_15762_, _15617_, _23676_);
  or (_05672_, _15762_, _15761_);
  and (_15763_, _05322_, _24078_);
  and (_15764_, _15763_, _23982_);
  not (_15765_, _15763_);
  and (_15766_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_05702_, _15766_, _15764_);
  and (_15767_, _10518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_15768_, _10517_, _23791_);
  or (_05711_, _15768_, _15767_);
  and (_15769_, _15763_, _23791_);
  and (_15770_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_05713_, _15770_, _15769_);
  and (_15771_, _23982_, _23644_);
  and (_15772_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_05716_, _15772_, _15771_);
  and (_15773_, _08428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_15774_, _08427_, _23838_);
  or (_27050_, _15774_, _15773_);
  and (_15775_, _06298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and (_15776_, _06296_, _23982_);
  or (_05722_, _15776_, _15775_);
  and (_15777_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and (_15778_, _15617_, _23982_);
  or (_05725_, _15778_, _15777_);
  and (_15779_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_15780_, _05420_, _23589_);
  or (_05729_, _15780_, _15779_);
  and (_15781_, _24573_, _23838_);
  and (_15782_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or (_05731_, _15782_, _15781_);
  and (_15783_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  and (_15784_, _15617_, _23838_);
  or (_05734_, _15784_, _15783_);
  and (_15785_, _05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and (_15786_, _05407_, _23589_);
  or (_05737_, _15786_, _15785_);
  and (_15787_, _04811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  and (_15788_, _04810_, _23791_);
  or (_05742_, _15788_, _15787_);
  and (_15789_, _04793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_15790_, _04792_, _23718_);
  or (_05745_, _15790_, _15789_);
  and (_15791_, _04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_15792_, _04756_, _23755_);
  or (_05748_, _15792_, _15791_);
  and (_15793_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and (_15794_, _09523_, _23718_);
  or (_27056_, _15794_, _15793_);
  and (_15795_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and (_15796_, _04734_, _23589_);
  or (_27032_, _15796_, _15795_);
  and (_15797_, _04733_, _24078_);
  not (_15798_, _15797_);
  and (_15799_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  and (_15800_, _15797_, _23838_);
  or (_27015_, _15800_, _15799_);
  and (_15801_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  and (_15802_, _15797_, _23718_);
  or (_05812_, _15802_, _15801_);
  and (_15803_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  and (_15804_, _10557_, _23982_);
  or (_05818_, _15804_, _15803_);
  and (_15805_, _12469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_15806_, _12468_, _23676_);
  or (_05828_, _15806_, _15805_);
  and (_15807_, _12600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_15808_, _12599_, _23718_);
  or (_05830_, _15808_, _15807_);
  and (_15809_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  and (_15810_, _13718_, _23635_);
  or (_05837_, _15810_, _15809_);
  and (_15811_, _03326_, _23718_);
  and (_15812_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_05841_, _15812_, _15811_);
  and (_15813_, _03326_, _23982_);
  and (_15814_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_05844_, _15814_, _15813_);
  and (_15815_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_15816_, _15563_, _23838_);
  or (_27019_, _15816_, _15815_);
  and (_15817_, _03326_, _23838_);
  and (_15818_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_27194_, _15818_, _15817_);
  and (_15819_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  and (_15820_, _15797_, _23791_);
  or (_05859_, _15820_, _15819_);
  and (_15821_, _04733_, _23649_);
  not (_15822_, _15821_);
  and (_15823_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_15824_, _15821_, _23838_);
  or (_05863_, _15824_, _15823_);
  and (_15825_, _03233_, _23017_);
  and (_15826_, _15825_, _23589_);
  not (_15827_, _15825_);
  and (_15828_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or (_05868_, _15828_, _15826_);
  and (_15829_, _03233_, _23849_);
  and (_15830_, _15829_, _23589_);
  not (_15831_, _15829_);
  and (_15832_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_05873_, _15832_, _15830_);
  and (_15833_, _15829_, _23676_);
  and (_15834_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_05878_, _15834_, _15833_);
  and (_15835_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  and (_15836_, _15797_, _23635_);
  or (_05880_, _15836_, _15835_);
  and (_15837_, _03233_, _23803_);
  and (_15838_, _15837_, _23676_);
  not (_15839_, _15837_);
  and (_15840_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_05883_, _15840_, _15838_);
  and (_15841_, _03233_, _23842_);
  and (_15842_, _15841_, _23718_);
  not (_15843_, _15841_);
  and (_15844_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or (_27006_, _15844_, _15842_);
  and (_15845_, _03233_, _23854_);
  and (_15846_, _15845_, _23718_);
  not (_15847_, _15845_);
  and (_15848_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or (_27005_, _15848_, _15846_);
  and (_15849_, _03233_, _23797_);
  and (_15850_, _15849_, _23982_);
  not (_15851_, _15849_);
  and (_15852_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_27004_, _15852_, _15850_);
  and (_15853_, _03233_, _24768_);
  and (_15854_, _15853_, _23755_);
  not (_15855_, _15853_);
  and (_15856_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_05897_, _15856_, _15854_);
  and (_15857_, _03233_, _24541_);
  and (_15858_, _15857_, _23791_);
  not (_15859_, _15857_);
  and (_15860_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or (_05902_, _15860_, _15858_);
  and (_15861_, _25407_, _23925_);
  nand (_15862_, _15861_, _23522_);
  or (_15863_, _15861_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_15864_, _15863_, _24629_);
  and (_15865_, _15864_, _15862_);
  nand (_15866_, _25413_, _23832_);
  or (_15867_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_15868_, _15867_, _23880_);
  and (_15869_, _15868_, _15866_);
  and (_15870_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_15871_, _15870_, rst);
  or (_15872_, _15871_, _15869_);
  or (_05905_, _15872_, _15865_);
  and (_15873_, _03233_, _23641_);
  and (_15874_, _15873_, _23791_);
  not (_15875_, _15873_);
  and (_15876_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or (_05910_, _15876_, _15874_);
  and (_15877_, _03233_, _24103_);
  and (_15878_, _15877_, _23755_);
  not (_15879_, _15877_);
  and (_15880_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_05915_, _15880_, _15878_);
  and (_15881_, _03234_, _23982_);
  and (_15882_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or (_05927_, _15882_, _15881_);
  and (_15883_, _25309_, _23986_);
  nand (_15884_, _15883_, _23522_);
  or (_15885_, _15883_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_15886_, _15885_, _24629_);
  and (_15887_, _15886_, _15884_);
  nand (_15888_, _25317_, _23914_);
  or (_15889_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_15890_, _15889_, _23880_);
  and (_15891_, _15890_, _15888_);
  and (_15892_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_15893_, _15892_, rst);
  or (_15894_, _15893_, _15891_);
  or (_05929_, _15894_, _15887_);
  and (_15895_, _05322_, _23017_);
  and (_15896_, _15895_, _23982_);
  not (_15897_, _15895_);
  and (_15898_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_05937_, _15898_, _15896_);
  nor (_26870_[2], _26830_, rst);
  and (_15899_, _05322_, _23803_);
  and (_15900_, _15899_, _23589_);
  not (_15901_, _15899_);
  and (_15902_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or (_05942_, _15902_, _15900_);
  and (_15903_, _03326_, _23755_);
  and (_15904_, _03328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_27195_, _15904_, _15903_);
  and (_15905_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_15906_, _15821_, _23589_);
  or (_05949_, _15906_, _15905_);
  and (_15907_, _15899_, _23838_);
  and (_15908_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or (_05969_, _15908_, _15907_);
  and (_15909_, _05322_, _23842_);
  and (_15910_, _15909_, _23838_);
  not (_15911_, _15909_);
  and (_15912_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_05982_, _15912_, _15910_);
  and (_15913_, _06264_, _23635_);
  and (_15914_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_05984_, _15914_, _15913_);
  and (_15915_, _06264_, _23791_);
  and (_15916_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_05987_, _15916_, _15915_);
  and (_15917_, _12516_, _23982_);
  and (_15918_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or (_05989_, _15918_, _15917_);
  and (_15919_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_15920_, _15821_, _23755_);
  or (_05992_, _15920_, _15919_);
  and (_15921_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_15922_, _15821_, _23635_);
  or (_05995_, _15922_, _15921_);
  and (_15923_, _25209_, _24688_);
  nand (_15924_, _15923_, _23522_);
  or (_15925_, _15923_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_15926_, _15925_, _24629_);
  and (_15927_, _15926_, _15924_);
  nand (_15928_, _25216_, _23748_);
  or (_15929_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_15930_, _15929_, _23880_);
  and (_15931_, _15930_, _15928_);
  and (_15932_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_15933_, _15932_, rst);
  or (_15934_, _15933_, _15931_);
  or (_05998_, _15934_, _15927_);
  and (_15935_, _05323_, _23791_);
  and (_15936_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or (_26972_, _15936_, _15935_);
  and (_15937_, _25118_, _23986_);
  nand (_15938_, _15937_, _23522_);
  or (_15939_, _15937_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_15940_, _15939_, _24629_);
  and (_15941_, _15940_, _15938_);
  nand (_15942_, _25124_, _23914_);
  or (_15943_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_15944_, _15943_, _23880_);
  and (_15945_, _15944_, _15942_);
  and (_15946_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_15947_, _15946_, rst);
  or (_15948_, _15947_, _15945_);
  or (_06005_, _15948_, _15941_);
  and (_15949_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  and (_15950_, _15797_, _23676_);
  or (_27014_, _15950_, _15949_);
  and (_15951_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  and (_15952_, _13434_, _23982_);
  or (_06024_, _15952_, _15951_);
  and (_15953_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  and (_15954_, _15463_, _23676_);
  or (_06028_, _15954_, _15953_);
  and (_15955_, _03241_, _23635_);
  and (_15956_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or (_06032_, _15956_, _15955_);
  and (_15957_, _03241_, _23982_);
  and (_15958_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or (_06034_, _15958_, _15957_);
  and (_15959_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and (_15960_, _15797_, _23589_);
  or (_06039_, _15960_, _15959_);
  and (_15961_, _03241_, _23838_);
  and (_15962_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or (_06048_, _15962_, _15961_);
  and (_15963_, _15873_, _23589_);
  and (_15964_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or (_06050_, _15964_, _15963_);
  and (_15965_, _15763_, _23718_);
  and (_15966_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_26949_, _15966_, _15965_);
  and (_15967_, _03233_, _23649_);
  and (_15968_, _15967_, _23791_);
  not (_15969_, _15967_);
  and (_15970_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_26984_, _15970_, _15968_);
  and (_15971_, _15763_, _23755_);
  and (_15972_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_26950_, _15972_, _15971_);
  nand (_15973_, _23921_, _23784_);
  and (_15974_, _24155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_15975_, _15974_, _24146_);
  nor (_15976_, _15975_, _24147_);
  and (_15977_, _13564_, _23938_);
  nor (_15978_, _15977_, _24182_);
  nor (_15979_, _15978_, _15976_);
  not (_15980_, _15979_);
  nor (_15981_, _15980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_15982_, _15980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_15983_, _15982_, _15981_);
  or (_15984_, _15983_, _23921_);
  and (_15985_, _15984_, _23928_);
  and (_15986_, _15985_, _15973_);
  and (_15987_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_15988_, _15987_, _15986_);
  and (_06060_, _15988_, _22761_);
  and (_15989_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_15990_, _15821_, _23676_);
  or (_06068_, _15990_, _15989_);
  and (_15991_, _05323_, _23635_);
  and (_15992_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or (_06072_, _15992_, _15991_);
  and (_15993_, _07861_, _23838_);
  and (_15994_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_06087_, _15994_, _15993_);
  and (_15995_, _03233_, _23962_);
  and (_15996_, _15995_, _23982_);
  not (_15997_, _15995_);
  and (_15998_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or (_06091_, _15998_, _15996_);
  and (_15999_, _13719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  and (_16000_, _13718_, _23755_);
  or (_06096_, _16000_, _15999_);
  and (_16001_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_16002_, _15563_, _23982_);
  or (_06102_, _16002_, _16001_);
  and (_16003_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_16004_, _15821_, _23982_);
  or (_06105_, _16004_, _16003_);
  and (_16005_, _15837_, _23791_);
  and (_16006_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_06109_, _16006_, _16005_);
  nand (_16007_, _23927_, _23914_);
  and (_16008_, _13539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_16009_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_16010_, _16009_, _13580_);
  and (_16011_, _16010_, _13538_);
  and (_16012_, _24148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_16013_, _16012_, _23948_);
  and (_16014_, _16013_, _23938_);
  nand (_16015_, _16014_, _23942_);
  nor (_16016_, _16015_, _23921_);
  or (_16017_, _16016_, _16011_);
  or (_16018_, _16017_, _16008_);
  or (_16019_, _16018_, _23927_);
  and (_16020_, _16019_, _22761_);
  and (_06116_, _16020_, _16007_);
  and (_16021_, _03234_, _23635_);
  and (_16022_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or (_06119_, _16022_, _16021_);
  and (_16023_, _15895_, _23676_);
  and (_16024_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_06122_, _16024_, _16023_);
  and (_16025_, _15763_, _23589_);
  and (_16026_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_06128_, _16026_, _16025_);
  and (_16027_, _03241_, _23589_);
  and (_16028_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or (_06134_, _16028_, _16027_);
  and (_16029_, _03241_, _23755_);
  and (_16030_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  or (_06135_, _16030_, _16029_);
  and (_16031_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_16032_, _15821_, _23718_);
  or (_06141_, _16032_, _16031_);
  and (_16033_, _15877_, _23676_);
  and (_16034_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_06145_, _16034_, _16033_);
  and (_26893_, _26838_, _22761_);
  and (_16035_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_16036_, _15821_, _23791_);
  or (_06153_, _16036_, _16035_);
  and (_16037_, _05322_, _23962_);
  and (_16038_, _16037_, _23676_);
  not (_16039_, _16037_);
  and (_16040_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_26951_, _16040_, _16038_);
  and (_16041_, _15995_, _23676_);
  and (_16042_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or (_06160_, _16042_, _16041_);
  and (_16043_, _16037_, _23718_);
  and (_16044_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_26953_, _16044_, _16043_);
  and (_16045_, _15995_, _23838_);
  and (_16046_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or (_06163_, _16046_, _16045_);
  and (_16047_, _15995_, _23589_);
  and (_16048_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or (_06167_, _16048_, _16047_);
  and (_16049_, _15995_, _23635_);
  and (_16050_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  or (_06170_, _16050_, _16049_);
  and (_16051_, _07861_, _23718_);
  and (_16052_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_06173_, _16052_, _16051_);
  and (_16053_, _03250_, _23635_);
  and (_16054_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  or (_06180_, _16054_, _16053_);
  and (_16055_, _03250_, _23589_);
  and (_16056_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  or (_06182_, _16056_, _16055_);
  and (_16057_, _05323_, _23676_);
  and (_16058_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or (_06199_, _16058_, _16057_);
  and (_16059_, _05323_, _23982_);
  and (_16060_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or (_26973_, _16060_, _16059_);
  and (_16061_, _05323_, _23838_);
  and (_16062_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or (_06206_, _16062_, _16061_);
  nor (_26894_[4], _25915_, rst);
  and (_26895_[7], _26816_, _22761_);
  and (_16063_, _15825_, _23676_);
  and (_16064_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  or (_27013_, _16064_, _16063_);
  and (_16065_, _12516_, _23676_);
  and (_16066_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or (_06213_, _16066_, _16065_);
  and (_16067_, _12516_, _23718_);
  and (_16068_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or (_06219_, _16068_, _16067_);
  and (_16069_, _03250_, _23755_);
  and (_16070_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or (_06221_, _16070_, _16069_);
  and (_16071_, _15825_, _23718_);
  and (_16072_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or (_06226_, _16072_, _16071_);
  and (_16073_, _15825_, _23791_);
  and (_16074_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or (_06232_, _16074_, _16073_);
  and (_16075_, _15909_, _23676_);
  and (_16076_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_06237_, _16076_, _16075_);
  and (_16077_, _15909_, _23589_);
  and (_16078_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_26977_, _16078_, _16077_);
  and (_16079_, _15899_, _23635_);
  and (_16080_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or (_06249_, _16080_, _16079_);
  and (_16081_, _05322_, _23849_);
  and (_16082_, _16081_, _23838_);
  not (_16083_, _16081_);
  and (_16084_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or (_06252_, _16084_, _16082_);
  and (_16085_, _15895_, _23718_);
  and (_16086_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_26980_, _16086_, _16085_);
  and (_16087_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  and (_16088_, _09509_, _23791_);
  or (_27107_, _16088_, _16087_);
  and (_16089_, _15967_, _23676_);
  and (_16090_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_06263_, _16090_, _16089_);
  and (_16091_, _15825_, _23982_);
  and (_16092_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or (_06266_, _16092_, _16091_);
  and (_16093_, _15825_, _23755_);
  and (_16094_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or (_06272_, _16094_, _16093_);
  and (_16095_, _15967_, _23982_);
  and (_16096_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_06278_, _16096_, _16095_);
  and (_16097_, _03234_, _23791_);
  and (_16098_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or (_06287_, _16098_, _16097_);
  and (_16099_, _03233_, _23863_);
  and (_16100_, _16099_, _23982_);
  not (_16101_, _16099_);
  and (_16102_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or (_06291_, _16102_, _16100_);
  and (_16103_, _15825_, _23635_);
  and (_16104_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  or (_06295_, _16104_, _16103_);
  and (_16105_, _03241_, _23791_);
  and (_16106_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or (_27193_, _16106_, _16105_);
  and (_16107_, _16099_, _23589_);
  and (_16108_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or (_06297_, _16108_, _16107_);
  and (_16109_, _15873_, _23755_);
  and (_16110_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or (_27002_, _16110_, _16109_);
  and (_16111_, _03233_, _24117_);
  and (_16112_, _16111_, _23982_);
  not (_16113_, _16111_);
  and (_16114_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_06314_, _16114_, _16112_);
  and (_16115_, _16111_, _23791_);
  and (_16116_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_06319_, _16116_, _16115_);
  and (_16117_, _03241_, _23676_);
  and (_16118_, _03244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or (_06321_, _16118_, _16117_);
  and (_16119_, _16111_, _23589_);
  and (_16120_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_06324_, _16120_, _16119_);
  and (_16121_, _15857_, _23635_);
  and (_16122_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or (_06333_, _16122_, _16121_);
  nor (_16123_, _26608_, rst);
  and (_26897_, _16123_, _00320_);
  and (_16124_, _15845_, _23755_);
  and (_16125_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or (_06349_, _16125_, _16124_);
  and (_16126_, _15829_, _23838_);
  and (_16127_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_06354_, _16127_, _16126_);
  and (_26898_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _22761_);
  and (_16128_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_16129_, _22770_, _22824_);
  or (_16130_, _16129_, _16128_);
  and (_26891_[8], _16130_, _22761_);
  and (_16131_, _15841_, _23982_);
  and (_16132_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or (_27007_, _16132_, _16131_);
  or (_16133_, _01387_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_16134_, _01388_, _01329_);
  or (_16135_, _16134_, _00907_);
  and (_16136_, _16135_, _16133_);
  nand (_16137_, _16136_, _03836_);
  or (_16138_, _16136_, _03836_);
  and (_16139_, _16138_, _16137_);
  and (_16140_, _16139_, _00323_);
  and (_16141_, _00874_, _26608_);
  and (_16142_, _03869_, _26574_);
  and (_16143_, _26604_, _26833_);
  not (_16144_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_16145_, _01323_, _16144_);
  and (_16146_, _01323_, _16144_);
  or (_16147_, _16146_, _16145_);
  and (_16148_, _16147_, _00349_);
  and (_16149_, _26630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_16150_, _16149_, _16148_);
  or (_16151_, _16150_, _16143_);
  nor (_16152_, _16151_, _16142_);
  nand (_16153_, _16152_, _00320_);
  or (_16154_, _16153_, _16141_);
  or (_16155_, _16154_, _16140_);
  and (_16156_, _01398_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_16157_, _01398_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_16158_, _16157_, _16156_);
  or (_16159_, _16158_, _00320_);
  and (_16160_, _16159_, _22761_);
  and (_26899_[15], _16160_, _16155_);
  and (_16161_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _22761_);
  and (_16162_, _16161_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_16163_, _01788_, _16144_);
  and (_16164_, _01788_, _16144_);
  nor (_16165_, _16164_, _16163_);
  and (_16166_, _16165_, _01791_);
  nor (_16167_, _16165_, _01791_);
  or (_16168_, _16167_, _16166_);
  or (_16169_, _16168_, _25562_);
  or (_16170_, _25561_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_16171_, _16170_, _01834_);
  and (_16172_, _16171_, _16169_);
  or (_26900_[15], _16172_, _16162_);
  and (_16173_, _15829_, _23718_);
  and (_16174_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_06365_, _16174_, _16173_);
  and (_16175_, _15825_, _23838_);
  and (_16176_, _15827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or (_06372_, _16176_, _16175_);
  and (_16177_, _15829_, _23791_);
  and (_16178_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_06374_, _16178_, _16177_);
  and (_16179_, _02322_, _23635_);
  and (_16180_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_06378_, _16180_, _16179_);
  and (_16181_, _23849_, _23806_);
  and (_16182_, _16181_, _23676_);
  not (_16183_, _16181_);
  and (_16184_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_06382_, _16184_, _16182_);
  nand (_16185_, _23994_, _23585_);
  and (_16186_, _23997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_16187_, _24053_, _13606_);
  nor (_16188_, _16187_, _16186_);
  nand (_16189_, _16188_, _24054_);
  or (_16190_, _16189_, _23988_);
  and (_16191_, _16190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_16192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand (_16193_, _16192_, _24050_);
  or (_16194_, _16193_, _16188_);
  nor (_16195_, _16194_, _23988_);
  or (_16196_, _16195_, _16191_);
  or (_16197_, _16196_, _23994_);
  and (_16198_, _16197_, _22761_);
  and (_06385_, _16198_, _16185_);
  and (_16199_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  and (_16200_, _15797_, _23755_);
  or (_06389_, _16200_, _16199_);
  and (_16201_, _15798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  and (_16202_, _15797_, _23982_);
  or (_06392_, _16202_, _16201_);
  and (_16203_, _03250_, _23676_);
  and (_16204_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  or (_06394_, _16204_, _16203_);
  and (_16205_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and (_16206_, _15617_, _23635_);
  or (_27016_, _16206_, _16205_);
  and (_16207_, _15618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and (_16208_, _15617_, _23718_);
  or (_06400_, _16208_, _16207_);
  and (_16209_, _15564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_16210_, _15563_, _23676_);
  or (_06405_, _16210_, _16209_);
  and (_16211_, _15524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_16212_, _15523_, _23791_);
  or (_27020_, _16212_, _16211_);
  or (_16213_, _15686_, _26568_);
  or (_16214_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_16215_, _16214_, _23880_);
  and (_16216_, _16215_, _16213_);
  and (_16217_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_16218_, _15685_, _23522_);
  and (_16219_, _16214_, _24629_);
  and (_16220_, _16219_, _16218_);
  or (_16221_, _16220_, _16217_);
  or (_16222_, _16221_, _16216_);
  and (_06433_, _16222_, _22761_);
  or (_16223_, _15686_, _00484_);
  or (_16224_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_16225_, _16224_, _23880_);
  and (_16226_, _16225_, _16223_);
  and (_16227_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_16228_, _15684_, _23992_);
  nand (_16229_, _16228_, _23522_);
  or (_16230_, _16228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_16231_, _16230_, _24629_);
  and (_16232_, _16231_, _16229_);
  or (_16233_, _16232_, _16227_);
  or (_16234_, _16233_, _16226_);
  and (_06435_, _16234_, _22761_);
  or (_16235_, _15686_, _00408_);
  or (_16236_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_16237_, _16236_, _23880_);
  and (_16238_, _16237_, _16235_);
  and (_16239_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_16240_, _15684_, _23878_);
  nand (_16241_, _16240_, _23522_);
  or (_16242_, _16240_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_16243_, _16242_, _24629_);
  and (_16244_, _16243_, _16241_);
  or (_16245_, _16244_, _16239_);
  or (_16246_, _16245_, _16238_);
  and (_06437_, _16246_, _22761_);
  and (_16247_, _15829_, _23982_);
  and (_16248_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_06440_, _16248_, _16247_);
  and (_16249_, _15829_, _23755_);
  and (_16250_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_06442_, _16250_, _16249_);
  and (_16251_, _15829_, _23635_);
  and (_16252_, _15831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_06447_, _16252_, _16251_);
  nor (_16253_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_26901_, _16253_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  or (_16254_, _15686_, _00580_);
  or (_16255_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_16256_, _16255_, _23880_);
  and (_16257_, _16256_, _16254_);
  and (_16258_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_16259_, _15684_, _23925_);
  nand (_16260_, _16259_, _23522_);
  or (_16261_, _16259_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_16262_, _16261_, _24629_);
  and (_16263_, _16262_, _16260_);
  or (_16264_, _16263_, _16258_);
  or (_16265_, _16264_, _16257_);
  and (_06450_, _16265_, _22761_);
  and (_16266_, _15464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  and (_16267_, _15463_, _23589_);
  or (_06453_, _16267_, _16266_);
  or (_16268_, _15686_, _00708_);
  or (_16269_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_16270_, _16269_, _23880_);
  and (_16271_, _16270_, _16268_);
  and (_16272_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_16273_, _15684_, _23919_);
  nand (_16274_, _16273_, _23522_);
  or (_16275_, _16273_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_16276_, _16275_, _24629_);
  and (_16277_, _16276_, _16274_);
  or (_16278_, _16277_, _16272_);
  or (_16279_, _16278_, _16271_);
  and (_06456_, _16279_, _22761_);
  or (_16280_, _15686_, _00647_);
  or (_16281_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_16282_, _16281_, _23880_);
  and (_16283_, _16282_, _16280_);
  and (_16284_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_16285_, _15684_);
  or (_16286_, _16285_, _24728_);
  and (_16287_, _16286_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_16288_, _23012_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_16289_, _16288_, _24732_);
  and (_16290_, _16289_, _15684_);
  or (_16291_, _16290_, _16287_);
  and (_16292_, _16291_, _24629_);
  or (_16293_, _16292_, _16284_);
  or (_16294_, _16293_, _16283_);
  and (_06459_, _16294_, _22761_);
  and (_16295_, _03335_, _23589_);
  and (_16296_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_06461_, _16296_, _16295_);
  and (_16297_, _13525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_16298_, _13524_, _23982_);
  or (_06463_, _16298_, _16297_);
  nand (_16299_, _15685_, _00791_);
  or (_16300_, _15685_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_16301_, _16300_, _23880_);
  and (_16302_, _16301_, _16299_);
  and (_16303_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_16304_, _15684_, _24688_);
  nand (_16305_, _16304_, _23522_);
  or (_16306_, _16304_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_16307_, _16306_, _24629_);
  and (_16308_, _16307_, _16305_);
  or (_16309_, _16308_, _16303_);
  or (_16310_, _16309_, _16302_);
  and (_06465_, _16310_, _22761_);
  and (_16311_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  and (_16312_, _13434_, _23838_);
  or (_06468_, _16312_, _16311_);
  and (_16313_, _13435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  and (_16314_, _13434_, _23589_);
  or (_06473_, _16314_, _16313_);
  and (_26902_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _22761_);
  nand (_16315_, _22768_, _01573_);
  nand (_16316_, _16315_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_16317_, _16316_, _01815_);
  and (_26903_, _16317_, _22761_);
  and (_16318_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  and (_16319_, _10557_, _23791_);
  or (_27030_, _16319_, _16318_);
  and (_16320_, _04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and (_16321_, _04734_, _23791_);
  or (_06498_, _16321_, _16320_);
  and (_16322_, _15837_, _23982_);
  and (_16323_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_27010_, _16323_, _16322_);
  and (_16324_, _10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  and (_16325_, _10557_, _23589_);
  or (_27031_, _16325_, _16324_);
  and (_16326_, _15837_, _23838_);
  and (_16327_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_06518_, _16327_, _16326_);
  and (_16328_, _03250_, _23718_);
  and (_16329_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or (_06520_, _16329_, _16328_);
  and (_16330_, _15837_, _23718_);
  and (_16331_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_06523_, _16331_, _16330_);
  and (_16332_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _22761_);
  and (_16333_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _22761_);
  and (_16334_, _16333_, _01815_);
  or (_26904_[7], _16334_, _16332_);
  nor (_16335_, _25781_, _25566_);
  nor (_16336_, _01841_, _01838_);
  nor (_16337_, _16336_, _25566_);
  and (_16338_, _16337_, _24237_);
  nor (_16339_, _16337_, _24237_);
  nor (_16340_, _16339_, _16338_);
  nor (_16341_, _16340_, _16335_);
  and (_16342_, _24248_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_16343_, _16342_, _16335_);
  nor (_16344_, _16343_, _01560_);
  or (_16345_, _16344_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_16346_, _16345_, _16341_);
  and (_26905_[2], _16346_, _22761_);
  or (_16347_, _24039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_16348_, _24038_, _22761_);
  and (_16349_, _16348_, _16347_);
  not (_16350_, _24039_);
  or (_16351_, _16350_, _24006_);
  nand (_16352_, _16351_, _16349_);
  nor (_16353_, _16352_, _23994_);
  and (_06553_, _16353_, _13625_);
  and (_16354_, _13706_, _23791_);
  and (_16355_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or (_06556_, _16355_, _16354_);
  and (_16356_, _03250_, _23791_);
  and (_16357_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  or (_06559_, _16357_, _16356_);
  and (_16358_, _15837_, _23589_);
  and (_16359_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_06584_, _16359_, _16358_);
  and (_16360_, _07101_, _23982_);
  and (_16361_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or (_06592_, _16361_, _16360_);
  and (_16362_, _15837_, _23755_);
  and (_16363_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_27012_, _16363_, _16362_);
  and (_16364_, _15837_, _23635_);
  and (_16365_, _15839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_27011_, _16365_, _16364_);
  and (_06619_, _26842_, _22761_);
  and (_06641_, _26794_, _22761_);
  and (_16366_, _03335_, _23718_);
  and (_16367_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_06643_, _16367_, _16366_);
  and (_16368_, _02342_, _23635_);
  and (_16369_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_06650_, _16369_, _16368_);
  and (_16370_, _15841_, _23838_);
  and (_16371_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or (_06657_, _16371_, _16370_);
  and (_16372_, _03335_, _23635_);
  and (_16373_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_06689_, _16373_, _16372_);
  and (_16374_, _13706_, _23838_);
  and (_16375_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or (_06698_, _16375_, _16374_);
  and (_16376_, _15841_, _23589_);
  and (_16377_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or (_06700_, _16377_, _16376_);
  and (_16378_, _15841_, _23755_);
  and (_16379_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or (_27009_, _16379_, _16378_);
  and (_16380_, _03335_, _23982_);
  and (_16381_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_06713_, _16381_, _16380_);
  and (_16382_, _15841_, _23635_);
  and (_16383_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  or (_27008_, _16383_, _16382_);
  and (_16384_, _07101_, _23838_);
  and (_16385_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or (_06722_, _16385_, _16384_);
  and (_16386_, _13706_, _23718_);
  and (_16387_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or (_06741_, _16387_, _16386_);
  and (_16388_, _23599_, _23017_);
  and (_16389_, _16388_, _23589_);
  not (_16390_, _16388_);
  and (_16391_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_06744_, _16391_, _16389_);
  and (_16392_, _15845_, _23838_);
  and (_16393_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  or (_06750_, _16393_, _16392_);
  and (_16394_, _15845_, _23635_);
  and (_16395_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or (_06756_, _16395_, _16394_);
  and (_16396_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  and (_16397_, _09509_, _23635_);
  or (_06762_, _16397_, _16396_);
  and (_16398_, _15845_, _23982_);
  and (_16399_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or (_06771_, _16399_, _16398_);
  and (_16400_, _06373_, _23635_);
  and (_16401_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_06785_, _16401_, _16400_);
  and (_16402_, _06373_, _23982_);
  and (_16403_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_06808_, _16403_, _16402_);
  and (_16404_, _15845_, _23589_);
  and (_16405_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or (_06819_, _16405_, _16404_);
  and (_16406_, _15841_, _23791_);
  and (_16407_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or (_06825_, _16407_, _16406_);
  and (_16408_, _15841_, _23676_);
  and (_16409_, _15843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  or (_06830_, _16409_, _16408_);
  and (_16410_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_16411_, _25845_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_16412_, _16411_, _16410_);
  and (_26912_[31], _16412_, _22761_);
  or (_16413_, _25781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_16414_, _25845_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_16415_, _16414_, _22761_);
  and (_26913_[31], _16415_, _16413_);
  and (_16416_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _01853_);
  and (_16417_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_16418_, _16417_, _16416_);
  and (_26908_[7], _16418_, _22761_);
  and (_26909_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _22761_);
  not (_16419_, _01883_);
  and (_16420_, _01886_, _16419_);
  and (_16421_, _26911_[3], _01891_);
  and (_26910_, _16421_, _16420_);
  and (_16422_, _06373_, _23589_);
  and (_16423_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_06888_, _16423_, _16422_);
  and (_16424_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_16425_, _04776_, _23838_);
  or (_06890_, _16425_, _16424_);
  and (_16426_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_16427_, _04776_, _23791_);
  or (_06892_, _16427_, _16426_);
  nand (_06894_, _00169_, _22761_);
  and (_16428_, _15849_, _23755_);
  and (_16429_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_06897_, _16429_, _16428_);
  nand (_06900_, _00187_, _22761_);
  and (_16430_, _15849_, _23635_);
  and (_16431_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_06904_, _16431_, _16430_);
  and (_06908_, _00099_, _22761_);
  nor (_06909_, _00116_, rst);
  nand (_06911_, _00210_, _22761_);
  and (_16432_, _04777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_16433_, _04776_, _23676_);
  or (_06914_, _16433_, _16432_);
  nor (_06916_, _00041_, rst);
  nor (_06918_, _00001_, rst);
  and (_16434_, _09510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  and (_16435_, _09509_, _23982_);
  or (_06923_, _16435_, _16434_);
  and (_16436_, _02237_, _23635_);
  and (_16437_, _02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_06925_, _16437_, _16436_);
  and (_16438_, _13485_, _23838_);
  and (_16439_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_26969_, _16439_, _16438_);
  and (_16440_, _13485_, _23791_);
  and (_16441_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_06928_, _16441_, _16440_);
  and (_26916_, _02054_, _22761_);
  and (_16442_, _26909_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_26915_, _16442_, _26916_);
  and (_16443_, _05322_, _24117_);
  and (_16444_, _16443_, _23718_);
  not (_16445_, _16443_);
  and (_16446_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or (_06956_, _16446_, _16444_);
  and (_16447_, _05322_, _23641_);
  and (_16448_, _16447_, _23755_);
  not (_16449_, _16447_);
  and (_16450_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_06962_, _16450_, _16448_);
  and (_16451_, _15845_, _23791_);
  and (_16452_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or (_06966_, _16452_, _16451_);
  and (_16453_, _16447_, _23791_);
  and (_16454_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_06970_, _16454_, _16453_);
  and (_16455_, _05322_, _23863_);
  and (_16456_, _16455_, _23755_);
  not (_16457_, _16455_);
  and (_16458_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_06973_, _16458_, _16456_);
  and (_16459_, _15845_, _23676_);
  and (_16460_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or (_06975_, _16460_, _16459_);
  and (_16461_, _16455_, _23791_);
  and (_16462_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_06982_, _16462_, _16461_);
  and (_16463_, _05322_, _24103_);
  and (_16464_, _16463_, _23589_);
  not (_16465_, _16463_);
  and (_16466_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or (_26956_, _16466_, _16464_);
  and (_16467_, _06373_, _23676_);
  and (_16468_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_06986_, _16468_, _16467_);
  and (_16469_, _15849_, _23589_);
  and (_16470_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_06988_, _16470_, _16469_);
  and (_16471_, _16463_, _23718_);
  and (_16472_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or (_06994_, _16472_, _16471_);
  and (_16473_, _16463_, _23676_);
  and (_16474_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or (_06999_, _16474_, _16473_);
  and (_16475_, _05322_, _23594_);
  and (_16476_, _16475_, _23755_);
  not (_16477_, _16475_);
  and (_16478_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or (_07004_, _16478_, _16476_);
  and (_16479_, _16475_, _23718_);
  and (_16480_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or (_07009_, _16480_, _16479_);
  and (_16481_, _16037_, _23589_);
  and (_16482_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_07013_, _16482_, _16481_);
  and (_16483_, _05322_, _23649_);
  and (_16484_, _16483_, _23755_);
  not (_16485_, _16483_);
  and (_16486_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or (_07017_, _16486_, _16484_);
  and (_16487_, _16483_, _23982_);
  and (_16488_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or (_26948_, _16488_, _16487_);
  and (_16489_, _15853_, _23589_);
  and (_16490_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_07020_, _16490_, _16489_);
  and (_16491_, _24577_, _23755_);
  and (_16492_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or (_07023_, _16492_, _16491_);
  and (_16493_, _15849_, _23791_);
  and (_16494_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_07027_, _16494_, _16493_);
  and (_16495_, _15849_, _23676_);
  and (_16496_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_07042_, _16496_, _16495_);
  and (_16497_, _23806_, _23017_);
  and (_16498_, _16497_, _23589_);
  not (_16499_, _16497_);
  and (_16500_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or (_07046_, _16500_, _16498_);
  and (_16501_, _16497_, _23838_);
  and (_16502_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or (_07067_, _16502_, _16501_);
  and (_16503_, _16181_, _23838_);
  and (_16504_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_07078_, _16504_, _16503_);
  and (_16505_, _02069_, _23982_);
  and (_16506_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_07080_, _16506_, _16505_);
  and (_16507_, _24577_, _23635_);
  and (_16508_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or (_07082_, _16508_, _16507_);
  and (_16509_, _16037_, _23791_);
  and (_16510_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_26952_, _16510_, _16509_);
  and (_16511_, _06373_, _23718_);
  and (_16512_, _06376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_07089_, _16512_, _16511_);
  and (_16513_, _23641_, _23599_);
  and (_16514_, _16513_, _23982_);
  not (_16515_, _16513_);
  and (_16516_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_27246_, _16516_, _16514_);
  and (_16517_, _15763_, _23838_);
  and (_16518_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_07098_, _16518_, _16517_);
  and (_16519_, _15849_, _23838_);
  and (_16520_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_07100_, _16520_, _16519_);
  and (_16521_, _15763_, _23635_);
  and (_16522_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_07106_, _16522_, _16521_);
  and (_16523_, _15849_, _23718_);
  and (_16524_, _15851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_07114_, _16524_, _16523_);
  and (_16525_, _16443_, _23982_);
  and (_16526_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or (_07117_, _16526_, _16525_);
  and (_16527_, _16447_, _23838_);
  and (_16528_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_07121_, _16528_, _16527_);
  and (_16529_, _16455_, _23838_);
  and (_16530_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_07125_, _16530_, _16529_);
  and (_16531_, _16463_, _23982_);
  and (_16532_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or (_07131_, _16532_, _16531_);
  and (_16533_, _16483_, _23791_);
  and (_16534_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or (_07141_, _16534_, _16533_);
  and (_16535_, _02069_, _23718_);
  and (_16536_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_27252_, _16536_, _16535_);
  and (_16537_, _15853_, _23718_);
  and (_16538_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_07148_, _16538_, _16537_);
  and (_16539_, _16497_, _23676_);
  and (_16540_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or (_07169_, _16540_, _16539_);
  and (_16541_, _16181_, _23635_);
  and (_16542_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_07173_, _16542_, _16541_);
  and (_16543_, _03260_, _23755_);
  and (_16544_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_07175_, _16544_, _16543_);
  and (_16545_, _15853_, _23791_);
  and (_16546_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_07178_, _16546_, _16545_);
  and (_16547_, _16037_, _23838_);
  and (_16548_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_07184_, _16548_, _16547_);
  and (_16549_, _15853_, _23676_);
  and (_16550_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_07187_, _16550_, _16549_);
  and (_16551_, _03260_, _23635_);
  and (_16552_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_07189_, _16552_, _16551_);
  and (_16553_, _16513_, _23838_);
  and (_16554_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_27245_, _16554_, _16553_);
  and (_16555_, _16447_, _23589_);
  and (_16556_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_07195_, _16556_, _16555_);
  and (_16557_, _16455_, _23589_);
  and (_16558_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_07197_, _16558_, _16557_);
  and (_16559_, _16475_, _23838_);
  and (_16560_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or (_26954_, _16560_, _16559_);
  and (_16561_, _15763_, _23676_);
  and (_16562_, _15765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_07202_, _16562_, _16561_);
  not (_16563_, _06202_);
  and (_16564_, _06195_, _24713_);
  or (_16565_, _16564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_16566_, _16565_, _16563_);
  nand (_16567_, _16564_, _23522_);
  and (_16568_, _16567_, _16566_);
  and (_16569_, _06202_, _24763_);
  or (_16570_, _16569_, _16568_);
  and (_07206_, _16570_, _22761_);
  and (_16571_, _06195_, _23919_);
  or (_16572_, _16571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_16573_, _16572_, _16563_);
  nand (_16574_, _16571_, _23522_);
  and (_16575_, _16574_, _16573_);
  nor (_16576_, _16563_, _23628_);
  or (_16577_, _16576_, _16575_);
  and (_07208_, _16577_, _22761_);
  not (_16578_, _06195_);
  or (_16579_, _16578_, _24728_);
  and (_16580_, _16579_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_16581_, _16580_, _06202_);
  and (_16582_, _23012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_16583_, _16582_, _24732_);
  and (_16584_, _16583_, _06195_);
  or (_16585_, _16584_, _16581_);
  nand (_16586_, _06202_, _23914_);
  and (_16587_, _16586_, _22761_);
  and (_07211_, _16587_, _16585_);
  and (_16588_, _06195_, _23925_);
  or (_16589_, _16588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_16590_, _16589_, _16563_);
  nand (_16591_, _16588_, _23522_);
  and (_16592_, _16591_, _16590_);
  nor (_16593_, _16563_, _23832_);
  or (_16594_, _16593_, _16592_);
  and (_07213_, _16594_, _22761_);
  and (_16595_, _06195_, _23992_);
  or (_16596_, _16595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_16597_, _16596_, _16563_);
  nand (_16598_, _16595_, _23522_);
  and (_16599_, _16598_, _16597_);
  and (_16600_, _06202_, _23709_);
  or (_16601_, _16600_, _16599_);
  and (_07217_, _16601_, _22761_);
  and (_16602_, _06195_, _23878_);
  and (_16603_, _16602_, _23522_);
  nor (_16604_, _16602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_16605_, _16604_, _16603_);
  nand (_16606_, _16605_, _16563_);
  nand (_16607_, _06202_, _23784_);
  and (_16608_, _16607_, _22761_);
  and (_07219_, _16608_, _16606_);
  and (_16609_, _16497_, _23982_);
  and (_16610_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or (_07221_, _16610_, _16609_);
  and (_16611_, _16181_, _23791_);
  and (_16612_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_26947_, _16612_, _16611_);
  and (_16613_, _15853_, _23635_);
  and (_16614_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_07232_, _16614_, _16613_);
  and (_16615_, _16037_, _23982_);
  and (_16616_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_07239_, _16616_, _16615_);
  and (_16617_, _02342_, _23838_);
  and (_16618_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_27159_, _16618_, _16617_);
  and (_16619_, _15853_, _23982_);
  and (_16620_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_07247_, _16620_, _16619_);
  or (_16621_, _25674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_16622_, _25682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_16623_, _25683_, _25674_);
  and (_16624_, _16623_, _16622_);
  and (_16625_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_16626_, _16625_, _25701_);
  or (_16627_, _16626_, _16624_);
  and (_16628_, _16627_, _16621_);
  or (_16629_, _16628_, _25699_);
  nor (_16630_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_16631_, _16630_, _25667_);
  and (_16632_, _16631_, _16629_);
  and (_16633_, _25667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_16634_, _16633_, _25711_);
  or (_16635_, _16634_, _16632_);
  nand (_16636_, _25711_, _23669_);
  and (_16637_, _16636_, _22761_);
  and (_07249_, _16637_, _16635_);
  and (_16638_, _15853_, _23838_);
  and (_16639_, _15855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_07252_, _16639_, _16638_);
  nor (_16640_, _10470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_16641_, _16640_, _10471_);
  or (_16642_, _16641_, _25699_);
  and (_16643_, _10475_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_16644_, _16643_, _25701_);
  or (_16645_, _16644_, _16642_);
  or (_16646_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_16647_, _16646_, _25712_);
  and (_16648_, _16647_, _16645_);
  and (_16649_, _25667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_16650_, _16649_, _16648_);
  nor (_16651_, _25716_, _23914_);
  or (_16652_, _16651_, _16650_);
  and (_07255_, _16652_, _22761_);
  nand (_16653_, _25711_, _23832_);
  and (_16654_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_16655_, _16654_, _25674_);
  and (_16656_, _16655_, _25701_);
  not (_16657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_16658_, _25687_, _25674_);
  and (_16659_, _16658_, _16657_);
  nor (_16660_, _16659_, _10470_);
  or (_16661_, _16660_, _25699_);
  or (_16662_, _16661_, _16656_);
  nor (_16663_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_16664_, _16663_, _25667_);
  and (_16665_, _16664_, _16662_);
  and (_16666_, _25667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_16667_, _16666_, _25711_);
  or (_16668_, _16667_, _16665_);
  and (_16669_, _16668_, _22761_);
  and (_07273_, _16669_, _16653_);
  or (_16670_, _25716_, _23709_);
  and (_16671_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_16672_, _16671_, _25674_);
  and (_16673_, _16672_, _25701_);
  and (_16674_, _25685_, _25674_);
  or (_16675_, _16674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_16676_, _16675_, _16658_);
  or (_16677_, _16676_, _25699_);
  or (_16678_, _16677_, _16673_);
  nor (_16679_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_16680_, _16679_, _25667_);
  and (_16681_, _16680_, _16678_);
  and (_16682_, _25667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_16683_, _16682_, _25711_);
  or (_16684_, _16683_, _16681_);
  and (_16685_, _16684_, _22761_);
  and (_07275_, _16685_, _16670_);
  nand (_16686_, _25711_, _23784_);
  and (_16687_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_16688_, _16687_, _25674_);
  and (_16689_, _16688_, _25701_);
  and (_16690_, _16623_, _13439_);
  nor (_16691_, _16690_, _16674_);
  or (_16692_, _16691_, _25699_);
  or (_16693_, _16692_, _16689_);
  nor (_16694_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_16695_, _16694_, _25667_);
  and (_16696_, _16695_, _16693_);
  and (_16697_, _25667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_16698_, _16697_, _25711_);
  or (_16699_, _16698_, _16696_);
  and (_16700_, _16699_, _22761_);
  and (_07277_, _16700_, _16686_);
  and (_16701_, _15481_, _23838_);
  and (_16702_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_07283_, _16702_, _16701_);
  and (_16703_, _23854_, _23028_);
  and (_16704_, _16703_, _23635_);
  not (_16705_, _16703_);
  and (_16706_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or (_27280_, _16706_, _16704_);
  and (_16707_, _23797_, _23028_);
  and (_16708_, _16707_, _23791_);
  not (_16709_, _16707_);
  and (_16710_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_07291_, _16710_, _16708_);
  and (_16711_, _02785_, _23791_);
  and (_16712_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  or (_07294_, _16712_, _16711_);
  and (_16713_, _24542_, _23635_);
  and (_16714_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_07298_, _16714_, _16713_);
  and (_16715_, _02785_, _23676_);
  and (_16716_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or (_07300_, _16716_, _16715_);
  and (_16717_, _02862_, _23589_);
  and (_16718_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_07304_, _16718_, _16717_);
  and (_16719_, _02326_, _23676_);
  and (_16720_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or (_07311_, _16720_, _16719_);
  nor (_16721_, _06164_, _23748_);
  and (_16722_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_16723_, _16722_, _25674_);
  and (_16724_, _16723_, _25701_);
  and (_16725_, _25680_, _25674_);
  or (_16726_, _16725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_16727_, _16726_, _06171_);
  or (_16728_, _16727_, _25699_);
  or (_16729_, _16728_, _16724_);
  nor (_16730_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_16731_, _16730_, _25667_);
  and (_16732_, _16731_, _16729_);
  or (_16733_, _16732_, _25711_);
  or (_16734_, _16733_, _16721_);
  or (_16735_, _25716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_16736_, _16735_, _22761_);
  and (_07314_, _16736_, _16734_);
  nor (_16737_, _06164_, _23628_);
  and (_16738_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_16739_, _16738_, _25674_);
  and (_16740_, _16739_, _25701_);
  and (_16741_, _25679_, _25674_);
  nor (_16742_, _16741_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_16743_, _16742_, _16725_);
  or (_16744_, _16743_, _25699_);
  or (_16745_, _16744_, _16740_);
  nor (_16746_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_16747_, _16746_, _25667_);
  and (_16748_, _16747_, _16745_);
  or (_16749_, _16748_, _25711_);
  or (_16750_, _16749_, _16737_);
  or (_16751_, _25716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_16752_, _16751_, _22761_);
  and (_07316_, _16752_, _16750_);
  and (_16753_, _25742_, _23791_);
  and (_16754_, _25744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_07318_, _16754_, _16753_);
  nor (_16755_, _06164_, _23914_);
  and (_16756_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_16757_, _16756_, _25674_);
  and (_16758_, _16757_, _25701_);
  and (_16759_, _25678_, _25674_);
  nor (_16760_, _16759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_16761_, _16760_, _16741_);
  or (_16762_, _16761_, _25699_);
  or (_16763_, _16762_, _16758_);
  nor (_16764_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_16765_, _16764_, _25667_);
  and (_16766_, _16765_, _16763_);
  or (_16767_, _16766_, _25711_);
  or (_16768_, _16767_, _16755_);
  or (_16769_, _25716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_16770_, _16769_, _22761_);
  and (_07320_, _16770_, _16768_);
  or (_16771_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_16772_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_16773_, _16772_, _25674_);
  and (_16774_, _16773_, _25701_);
  and (_16775_, _25677_, _25674_);
  nor (_16776_, _16775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_16777_, _16776_, _16759_);
  or (_16778_, _16777_, _25699_);
  or (_16779_, _16778_, _16774_);
  nand (_16780_, _16779_, _16771_);
  nand (_16781_, _16780_, _06164_);
  nand (_16782_, _25667_, _23832_);
  and (_16783_, _16782_, _16781_);
  or (_16784_, _16783_, _25711_);
  or (_16785_, _25716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_16786_, _16785_, _22761_);
  and (_07323_, _16786_, _16784_);
  and (_16787_, _25667_, _23709_);
  and (_16788_, _25703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_16789_, _16788_, _25674_);
  and (_16790_, _16789_, _25701_);
  not (_16791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand (_16792_, _25676_, _25674_);
  and (_16793_, _16792_, _16791_);
  nor (_16794_, _16793_, _16775_);
  or (_16795_, _16794_, _25699_);
  or (_16796_, _16795_, _16790_);
  nor (_16797_, _25709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor (_16798_, _16797_, _25667_);
  and (_16799_, _16798_, _16796_);
  or (_16800_, _16799_, _25711_);
  or (_16801_, _16800_, _16787_);
  nand (_16802_, _25711_, _16791_);
  and (_16803_, _16802_, _22761_);
  and (_07325_, _16803_, _16801_);
  or (_16804_, _10450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_16805_, _16804_, _16792_);
  and (_16806_, _10475_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_16807_, _16806_, _25701_);
  or (_16808_, _16807_, _16805_);
  and (_16809_, _16808_, _25709_);
  and (_16810_, _25699_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nor (_16811_, _16810_, _16809_);
  nand (_16812_, _16811_, _06164_);
  nand (_16813_, _25667_, _23784_);
  and (_16814_, _16813_, _16812_);
  or (_16815_, _16814_, _25711_);
  or (_16816_, _25716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_16817_, _16816_, _22761_);
  and (_07327_, _16817_, _16815_);
  and (_16818_, _15857_, _23982_);
  and (_16819_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or (_07330_, _16819_, _16818_);
  and (_16820_, _16181_, _23718_);
  and (_16821_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_07333_, _16821_, _16820_);
  and (_16822_, _15503_, _23791_);
  and (_16823_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_07335_, _16823_, _16822_);
  and (_16824_, _16181_, _23982_);
  and (_16825_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_07338_, _16825_, _16824_);
  nand (_16826_, _02073_, _23832_);
  or (_16827_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nand (_16828_, _02078_, _16657_);
  and (_16829_, _16828_, _16827_);
  or (_16830_, _16829_, _02073_);
  and (_16831_, _16830_, _22761_);
  and (_07339_, _16831_, _16826_);
  and (_16832_, _16388_, _23676_);
  and (_16833_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_07342_, _16833_, _16832_);
  and (_16834_, _15857_, _23838_);
  and (_16835_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  or (_07345_, _16835_, _16834_);
  nand (_16836_, _02073_, _23748_);
  and (_16837_, _09498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_16838_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_16839_, _16838_, _16837_);
  or (_16840_, _16839_, _02073_);
  and (_16841_, _16840_, _22761_);
  and (_07347_, _16841_, _16836_);
  and (_16842_, _15857_, _23718_);
  and (_16843_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or (_07350_, _16843_, _16842_);
  nand (_16844_, _02073_, _23628_);
  or (_16845_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand (_16846_, _02078_, _10468_);
  and (_16847_, _16846_, _16845_);
  or (_16848_, _16847_, _02073_);
  and (_16849_, _16848_, _22761_);
  and (_07352_, _16849_, _16844_);
  and (_16850_, _23803_, _23599_);
  and (_16851_, _16850_, _23838_);
  not (_16852_, _16850_);
  and (_16853_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or (_07355_, _16853_, _16851_);
  nand (_16854_, _02073_, _23914_);
  and (_16855_, _09498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_16856_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_16857_, _16856_, _16855_);
  or (_16858_, _16857_, _02073_);
  and (_16859_, _16858_, _22761_);
  and (_07358_, _16859_, _16854_);
  or (_16860_, _04740_, _23709_);
  and (_16861_, _09498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_16862_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_16863_, _16862_, _16861_);
  or (_16864_, _16863_, _02073_);
  and (_16865_, _16864_, _22761_);
  and (_07360_, _16865_, _16860_);
  and (_16866_, _02069_, _23635_);
  and (_16867_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_07362_, _16867_, _16866_);
  and (_16868_, _23798_, _23589_);
  and (_16869_, _23800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or (_07364_, _16869_, _16868_);
  and (_16870_, _03001_, _23589_);
  and (_16871_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or (_07367_, _16871_, _16870_);
  and (_16872_, _05287_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_16873_, _24472_, _24392_);
  or (_16874_, _16873_, _24514_);
  or (_16875_, _16874_, _24457_);
  or (_16876_, _26720_, _26596_);
  and (_16877_, _26692_, _24418_);
  or (_16878_, _16877_, _02243_);
  or (_16879_, _16878_, _16876_);
  or (_16880_, _16879_, _00272_);
  or (_16881_, _16880_, _05309_);
  or (_16882_, _16881_, _16875_);
  or (_16883_, _16882_, _05304_);
  and (_16884_, _16883_, _25615_);
  or (_26881_[0], _16884_, _16872_);
  and (_16885_, _03264_, _23589_);
  and (_16886_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_07395_, _16886_, _16885_);
  and (_16887_, _15857_, _23589_);
  and (_16888_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or (_27003_, _16888_, _16887_);
  and (_16889_, _23863_, _23599_);
  and (_16890_, _16889_, _23635_);
  not (_16891_, _16889_);
  and (_16892_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_07401_, _16892_, _16890_);
  and (_16893_, _03260_, _23676_);
  and (_16894_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_07404_, _16894_, _16893_);
  nand (_16895_, _02077_, _23748_);
  and (_16896_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_16897_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_16898_, _16897_, _16896_);
  or (_16899_, _16898_, _02077_);
  and (_16900_, _16899_, _04740_);
  and (_16901_, _16900_, _16895_);
  and (_16902_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_16903_, _16902_, _16901_);
  and (_07409_, _16903_, _22761_);
  nand (_16904_, _02077_, _23628_);
  and (_16905_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_16906_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_16907_, _16906_, _16905_);
  or (_16908_, _16907_, _02077_);
  and (_16910_, _16908_, _04740_);
  and (_16911_, _16910_, _16904_);
  and (_16912_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_16913_, _16912_, _16911_);
  and (_07411_, _16913_, _22761_);
  and (_16914_, _07861_, _23791_);
  and (_16915_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_07414_, _16915_, _16914_);
  and (_16916_, _05323_, _23589_);
  and (_16917_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or (_07416_, _16917_, _16916_);
  and (_16918_, _15857_, _23755_);
  and (_16919_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or (_07418_, _16919_, _16918_);
  and (_16920_, _06044_, _23635_);
  and (_16921_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_07420_, _16921_, _16920_);
  or (_16922_, _24288_, _02363_);
  or (_16923_, _22767_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_16924_, _16923_, _22761_);
  and (_26873_[2], _16924_, _16922_);
  and (_16925_, _02877_, _23635_);
  and (_16926_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_07423_, _16926_, _16925_);
  and (_16927_, _16181_, _23755_);
  and (_16928_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_07430_, _16928_, _16927_);
  and (_16929_, _02322_, _23755_);
  and (_16930_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_07432_, _16930_, _16929_);
  and (_16931_, _02322_, _23718_);
  and (_16932_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_07434_, _16932_, _16931_);
  and (_16933_, _02459_, _23635_);
  and (_16934_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or (_07437_, _16934_, _16933_);
  and (_16935_, _24104_, _23718_);
  and (_16936_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or (_27243_, _16936_, _16935_);
  and (_16937_, _23601_, _23589_);
  and (_16938_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or (_07442_, _16938_, _16937_);
  and (_16939_, _03260_, _23791_);
  and (_16940_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_07445_, _16940_, _16939_);
  and (_16941_, _16181_, _23589_);
  and (_16942_, _16183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_07448_, _16942_, _16941_);
  and (_16943_, _16111_, _23755_);
  and (_16944_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_07451_, _16944_, _16943_);
  and (_16945_, _25536_, _23676_);
  and (_16946_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_07452_, _16946_, _16945_);
  and (_16947_, _03260_, _23838_);
  and (_16948_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_07454_, _16948_, _16947_);
  and (_16949_, _16111_, _23635_);
  and (_16950_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_07460_, _16950_, _16949_);
  and (_16951_, _16497_, _23791_);
  and (_16952_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or (_07463_, _16952_, _16951_);
  not (_16953_, _02077_);
  or (_16954_, _16953_, _23709_);
  and (_16955_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_16956_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_16957_, _16956_, _16955_);
  or (_16958_, _16957_, _02077_);
  and (_16959_, _16958_, _04740_);
  and (_16960_, _16959_, _16954_);
  and (_16961_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_16962_, _16961_, _16960_);
  and (_07465_, _16962_, _22761_);
  nand (_16963_, _02077_, _23784_);
  and (_16964_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_16965_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_16966_, _16965_, _16964_);
  or (_16967_, _16966_, _02077_);
  and (_16968_, _16967_, _04740_);
  and (_16969_, _16968_, _16963_);
  and (_16970_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_16971_, _16970_, _16969_);
  and (_07467_, _16971_, _22761_);
  or (_16972_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_16973_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_16974_, _16973_, _16972_);
  or (_16975_, _16974_, _02077_);
  nand (_16976_, _02077_, _23669_);
  and (_16977_, _16976_, _16975_);
  or (_16978_, _16977_, _02073_);
  or (_16979_, _04740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_16980_, _16979_, _22761_);
  and (_07470_, _16980_, _16978_);
  and (_16981_, _24209_, _23791_);
  and (_16982_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_07471_, _16982_, _16981_);
  and (_16983_, _03260_, _23718_);
  and (_16984_, _03262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_07489_, _16984_, _16983_);
  and (_16985_, _03046_, _23982_);
  and (_16986_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_07495_, _16986_, _16985_);
  and (_16987_, _16497_, _23718_);
  and (_16988_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or (_07499_, _16988_, _16987_);
  and (_16989_, _15857_, _23676_);
  and (_16990_, _15859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  or (_07514_, _16990_, _16989_);
  and (_16991_, _02436_, _23755_);
  and (_16992_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or (_07526_, _16992_, _16991_);
  and (_16993_, _03264_, _23718_);
  and (_16994_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_07544_, _16994_, _16993_);
  and (_16995_, _06044_, _23982_);
  and (_16996_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_27235_, _16996_, _16995_);
  and (_16997_, _02877_, _23791_);
  and (_16998_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_07547_, _16998_, _16997_);
  and (_16999_, _03264_, _23791_);
  and (_17000_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_07552_, _17000_, _16999_);
  and (_17001_, _24118_, _23854_);
  and (_17002_, _17001_, _23676_);
  not (_17003_, _17001_);
  and (_17004_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or (_07783_, _17004_, _17002_);
  and (_17005_, _16111_, _23676_);
  and (_17006_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_07787_, _17006_, _17005_);
  and (_17007_, _16497_, _23635_);
  and (_17008_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or (_07789_, _17008_, _17007_);
  and (_17009_, _24769_, _23676_);
  and (_17010_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or (_07791_, _17010_, _17009_);
  and (_17011_, _03264_, _23635_);
  and (_17012_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_07805_, _17012_, _17011_);
  and (_17013_, _02862_, _23676_);
  and (_17014_, _02864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_07809_, _17014_, _17013_);
  and (_17015_, _03264_, _23982_);
  and (_17016_, _03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_27183_, _17016_, _17015_);
  and (_17017_, _15503_, _23718_);
  and (_17018_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_27261_, _17018_, _17017_);
  and (_17019_, _16850_, _23982_);
  and (_17020_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or (_07816_, _17020_, _17019_);
  and (_17021_, _16111_, _23838_);
  and (_17022_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_07819_, _17022_, _17021_);
  and (_17023_, _16111_, _23718_);
  and (_17024_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_07823_, _17024_, _17023_);
  and (_17025_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  and (_17027_, _13838_, _23635_);
  or (_07862_, _17027_, _17025_);
  and (_17028_, _24577_, _23676_);
  and (_17029_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or (_07864_, _17029_, _17028_);
  and (_17030_, _24104_, _23838_);
  and (_17031_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or (_07867_, _17031_, _17030_);
  and (_17032_, _25536_, _23755_);
  and (_17033_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_07868_, _17033_, _17032_);
  and (_17034_, _24209_, _23718_);
  and (_17035_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_07874_, _17035_, _17034_);
  and (_17036_, _15503_, _23838_);
  and (_17037_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_27262_, _17037_, _17036_);
  and (_17038_, _23803_, _23651_);
  and (_17039_, _17038_, _23718_);
  not (_17040_, _17038_);
  and (_17041_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or (_07882_, _17041_, _17039_);
  and (_17042_, _23842_, _23651_);
  and (_17043_, _17042_, _23755_);
  not (_17044_, _17042_);
  and (_17045_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_07887_, _17045_, _17043_);
  and (_17046_, _17042_, _23718_);
  and (_17047_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_07890_, _17047_, _17046_);
  and (_17048_, _17042_, _23676_);
  and (_17049_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_07892_, _17049_, _17048_);
  and (_17050_, _23854_, _23651_);
  and (_17051_, _17050_, _23589_);
  not (_17052_, _17050_);
  and (_17053_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_07896_, _17053_, _17051_);
  and (_17054_, _17050_, _23838_);
  and (_17055_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_07899_, _17055_, _17054_);
  and (_17056_, _17050_, _23791_);
  and (_17057_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_07902_, _17057_, _17056_);
  and (_17058_, _23797_, _23651_);
  and (_17059_, _17058_, _23838_);
  not (_17060_, _17058_);
  and (_17061_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or (_07907_, _17061_, _17059_);
  and (_17062_, _17058_, _23791_);
  and (_17063_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or (_07909_, _17063_, _17062_);
  and (_17064_, _24768_, _23651_);
  and (_17065_, _17064_, _23982_);
  not (_17066_, _17064_);
  and (_17067_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or (_07914_, _17067_, _17065_);
  and (_17068_, _17064_, _23718_);
  and (_17069_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or (_07916_, _17069_, _17068_);
  and (_17070_, _24541_, _23651_);
  and (_17071_, _17070_, _23635_);
  not (_17072_, _17070_);
  and (_17073_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_07920_, _17073_, _17071_);
  and (_17074_, _16497_, _23755_);
  and (_17075_, _16499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or (_07923_, _17075_, _17074_);
  and (_17076_, _17070_, _23791_);
  and (_17077_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_07925_, _17077_, _17076_);
  and (_17078_, _23863_, _23651_);
  and (_17079_, _17078_, _23589_);
  not (_17080_, _17078_);
  and (_17081_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_07934_, _17081_, _17079_);
  and (_17082_, _17078_, _23635_);
  and (_17083_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_07936_, _17083_, _17082_);
  and (_17084_, _03277_, _23635_);
  and (_17085_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or (_08160_, _17085_, _17084_);
  and (_17086_, _24103_, _23651_);
  and (_17087_, _17086_, _23635_);
  not (_17088_, _17086_);
  and (_17089_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_08161_, _17089_, _17087_);
  and (_17090_, _03277_, _23982_);
  and (_17091_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or (_08163_, _17091_, _17090_);
  and (_17092_, _15873_, _23838_);
  and (_17093_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  or (_27001_, _17093_, _17092_);
  and (_17094_, _17086_, _23838_);
  and (_17095_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or (_08167_, _17095_, _17094_);
  and (_17096_, _15873_, _23718_);
  and (_17097_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or (_08170_, _17097_, _17096_);
  and (_17098_, _23811_, _23755_);
  and (_17099_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or (_08172_, _17099_, _17098_);
  and (_17100_, _16388_, _23755_);
  and (_17101_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_08175_, _17101_, _17100_);
  and (_17102_, _03277_, _23838_);
  and (_17103_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or (_08177_, _17103_, _17102_);
  and (_17104_, _24117_, _23651_);
  and (_17105_, _17104_, _23838_);
  not (_17106_, _17104_);
  and (_17107_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or (_08184_, _17107_, _17105_);
  and (_17108_, _15873_, _23635_);
  and (_17109_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  or (_08189_, _17109_, _17108_);
  and (_17110_, _15873_, _23982_);
  and (_17111_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or (_08196_, _17111_, _17110_);
  and (_17112_, _23651_, _23641_);
  and (_17113_, _17112_, _23982_);
  not (_17114_, _17112_);
  and (_17115_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_08201_, _17115_, _17113_);
  and (_17116_, _17112_, _23589_);
  and (_17117_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_08203_, _17117_, _17116_);
  and (_17118_, _02300_, _24184_);
  and (_17119_, _24194_, _24191_);
  or (_17120_, _17119_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_17121_, _17120_, _17118_);
  nor (_17122_, _02306_, _23921_);
  and (_17123_, _17122_, _17121_);
  nor (_17124_, _23922_, _23914_);
  or (_17125_, _17124_, _17123_);
  and (_17126_, _17125_, _23928_);
  and (_17127_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_17128_, _17127_, _17126_);
  and (_08256_, _17128_, _22761_);
  or (_17129_, _24538_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_17130_, _26621_, _24418_);
  and (_17131_, _26577_, _26584_);
  and (_17132_, _26580_, _24443_);
  or (_17133_, _17132_, _17131_);
  or (_17134_, _17133_, _17130_);
  and (_17135_, _17134_, _26575_);
  and (_17136_, _17133_, _26571_);
  or (_17137_, _17136_, _17135_);
  or (_17138_, _17137_, _17129_);
  or (_17139_, _22765_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17140_, _17139_, _22761_);
  and (_26878_[2], _17140_, _17138_);
  or (_17141_, _24497_, _24449_);
  or (_17142_, _02038_, _01992_);
  or (_17143_, _17142_, _17141_);
  and (_17144_, _17143_, _22768_);
  nor (_17145_, _26826_, _24529_);
  and (_17146_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17147_, _17146_, _17145_);
  or (_17148_, _17147_, _17144_);
  and (_26875_[1], _17148_, _22761_);
  and (_17149_, _05287_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_17150_, _01997_, _26617_);
  or (_17151_, _02041_, _17150_);
  or (_17152_, _17151_, _17141_);
  and (_17153_, _26595_, _24486_);
  or (_17154_, _17153_, _05307_);
  or (_17155_, _17154_, _17152_);
  not (_17156_, _26659_);
  or (_17157_, _02026_, _17156_);
  or (_17158_, _17157_, _17155_);
  and (_17159_, _17158_, _25615_);
  or (_26876_[1], _17159_, _17149_);
  or (_17160_, _16877_, _26693_);
  and (_17161_, _24517_, _24416_);
  or (_17162_, _17161_, _26619_);
  or (_17163_, _17162_, _17160_);
  or (_17164_, _17130_, _02023_);
  or (_17165_, _26622_, _26592_);
  or (_17166_, _17165_, _17164_);
  or (_17167_, _17166_, _26590_);
  or (_17168_, _17167_, _17163_);
  and (_17169_, _17168_, _25615_);
  and (_17170_, _05287_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_26874_, _17170_, _17169_);
  and (_17171_, _05287_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_17172_, _01990_, _04057_);
  or (_17173_, _17172_, _24420_);
  or (_17174_, _26658_, _24456_);
  or (_17175_, _17174_, _17173_);
  not (_17176_, _26688_);
  nand (_17177_, _26708_, _17176_);
  or (_17178_, _17177_, _17175_);
  or (_17179_, _26697_, _26680_);
  or (_17180_, _02038_, _17150_);
  or (_17181_, _17180_, _17179_);
  or (_17182_, _17181_, _02026_);
  or (_17183_, _17182_, _17178_);
  or (_17184_, _04071_, _02035_);
  or (_17185_, _17184_, _02250_);
  or (_17186_, _17185_, _02263_);
  or (_17187_, _17186_, _17183_);
  and (_17188_, _17187_, _25615_);
  or (_26880_[3], _17188_, _17171_);
  and (_17189_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_17190_, _26732_, _22768_);
  or (_17191_, _17190_, _17189_);
  or (_17192_, _17191_, _17145_);
  and (_26877_[2], _17192_, _22761_);
  and (_17193_, _05287_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_17194_, _05293_, _24449_);
  and (_17195_, _26577_, _24447_);
  or (_17196_, _17195_, _17161_);
  or (_17197_, _17196_, _17194_);
  or (_17198_, _26711_, _05289_);
  or (_17199_, _17198_, _17197_);
  or (_17200_, _02031_, _05306_);
  or (_17201_, _17200_, _17199_);
  and (_17202_, _17201_, _25615_);
  or (_26879_[1], _17202_, _17193_);
  and (_17203_, _02937_, _23982_);
  and (_17204_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or (_08295_, _17204_, _17203_);
  and (_17205_, _02322_, _23838_);
  and (_17206_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_08301_, _17206_, _17205_);
  and (_17207_, _02379_, _23589_);
  and (_17208_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_08464_, _17208_, _17207_);
  nor (_26906_[0], _00341_, rst);
  and (_17210_, _25301_, _23635_);
  and (_17211_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_27091_, _17211_, _17210_);
  and (_17212_, _25301_, _23755_);
  and (_17213_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_08500_, _17213_, _17212_);
  and (_17214_, _02379_, _23982_);
  and (_17215_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_08507_, _17215_, _17214_);
  and (_17216_, _02379_, _23635_);
  and (_17217_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_08510_, _17217_, _17216_);
  and (_17218_, _25301_, _23982_);
  and (_17219_, _25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_08517_, _17219_, _17218_);
  and (_17220_, _02459_, _23676_);
  and (_17221_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or (_08529_, _17221_, _17220_);
  and (_17222_, _24475_, _24443_);
  and (_17223_, _17222_, _24489_);
  or (_17224_, _02002_, _17131_);
  or (_17225_, _17224_, _17223_);
  not (_17226_, _26716_);
  nand (_17227_, _17226_, _26708_);
  or (_17228_, _26732_, _02261_);
  or (_17229_, _17228_, _17227_);
  nand (_17230_, _26715_, _26696_);
  or (_17231_, _17230_, _17229_);
  or (_17232_, _17231_, _17225_);
  and (_17233_, _24470_, _24474_);
  or (_17234_, _17233_, _26728_);
  or (_17235_, _17234_, _17132_);
  or (_17236_, _17235_, _26650_);
  and (_17237_, _26656_, _24475_);
  or (_17238_, _17237_, _26658_);
  or (_17239_, _17238_, _26740_);
  and (_17240_, _24458_, _24475_);
  or (_17241_, _17240_, _26718_);
  or (_17242_, _17241_, _17150_);
  or (_17243_, _17242_, _01992_);
  or (_17244_, _17243_, _17239_);
  or (_17245_, _17244_, _17236_);
  or (_17246_, _17245_, _17232_);
  and (_17247_, _17246_, _22768_);
  and (_17248_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_17249_, _26585_, _26571_);
  or (_17250_, _17136_, _17145_);
  or (_17251_, _17250_, _17249_);
  or (_17252_, _17251_, _17248_);
  or (_17253_, _17252_, _17247_);
  and (_26882_, _17253_, _22761_);
  and (_17254_, _24104_, _23791_);
  and (_17255_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or (_08539_, _17255_, _17254_);
  and (_17256_, _02444_, _23755_);
  and (_17257_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_08543_, _17257_, _17256_);
  and (_17258_, _02444_, _23589_);
  and (_17259_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_08552_, _17259_, _17258_);
  and (_17260_, _02436_, _23676_);
  and (_17261_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or (_08570_, _17261_, _17260_);
  and (_17262_, _24542_, _23676_);
  and (_17263_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_08574_, _17263_, _17262_);
  nor (_26906_[2], _00504_, rst);
  and (_17264_, _23850_, _23676_);
  and (_17265_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or (_08593_, _17265_, _17264_);
  and (_17266_, _17042_, _23982_);
  and (_17267_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_08607_, _17267_, _17266_);
  and (_17268_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  and (_17269_, _13838_, _23982_);
  or (_08609_, _17269_, _17268_);
  and (_17270_, _17001_, _23791_);
  and (_17271_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or (_08627_, _17271_, _17270_);
  and (_17272_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  and (_17273_, _13764_, _23982_);
  or (_08682_, _17273_, _17272_);
  and (_17274_, _07861_, _23676_);
  and (_17275_, _07865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_08696_, _17275_, _17274_);
  and (_17276_, _17050_, _23635_);
  and (_17277_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_08701_, _17277_, _17276_);
  and (_17278_, _17058_, _23635_);
  and (_17279_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or (_08705_, _17279_, _17278_);
  and (_17280_, _17064_, _23755_);
  and (_17281_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or (_27305_, _17281_, _17280_);
  and (_17282_, _17112_, _23676_);
  and (_17283_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_08717_, _17283_, _17282_);
  and (_17284_, _16483_, _23676_);
  and (_17285_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or (_08718_, _17285_, _17284_);
  and (_17286_, _17078_, _23718_);
  and (_17287_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_08721_, _17287_, _17286_);
  and (_17288_, _17086_, _23589_);
  and (_17289_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or (_08723_, _17289_, _17288_);
  and (_17290_, _03277_, _23589_);
  and (_17291_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or (_08726_, _17291_, _17290_);
  and (_17292_, _03277_, _23755_);
  and (_17293_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  or (_08730_, _17293_, _17292_);
  and (_17294_, _17104_, _23635_);
  and (_17295_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_08733_, _17295_, _17294_);
  and (_17296_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  and (_17297_, _13764_, _23838_);
  or (_27105_, _17297_, _17296_);
  and (_17298_, _16513_, _23755_);
  and (_17299_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_08741_, _17299_, _17298_);
  and (_17300_, _16483_, _23718_);
  and (_17301_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or (_08761_, _17301_, _17300_);
  and (_17302_, _17038_, _23838_);
  and (_17303_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or (_27308_, _17303_, _17302_);
  and (_17304_, _16099_, _23755_);
  and (_17305_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or (_08772_, _17305_, _17304_);
  and (_17306_, _16099_, _23635_);
  and (_17307_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or (_08777_, _17307_, _17306_);
  and (_17308_, _16889_, _23589_);
  and (_17309_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_08787_, _17309_, _17308_);
  and (_17310_, _17058_, _23755_);
  and (_17311_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or (_08790_, _17311_, _17310_);
  and (_17312_, _23806_, _23797_);
  and (_17313_, _17312_, _23838_);
  not (_17314_, _17312_);
  and (_17315_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_08800_, _17315_, _17313_);
  and (_17316_, _24768_, _23806_);
  and (_17317_, _17316_, _23589_);
  not (_17318_, _17316_);
  and (_17319_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_26937_, _17319_, _17317_);
  and (_17320_, _17316_, _23635_);
  and (_17321_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_08806_, _17321_, _17320_);
  and (_17322_, _06290_, _23755_);
  and (_17323_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or (_08812_, _17323_, _17322_);
  and (_17324_, _17316_, _23676_);
  and (_17325_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_08815_, _17325_, _17324_);
  and (_17326_, _24541_, _23806_);
  and (_17327_, _17326_, _23755_);
  not (_17328_, _17326_);
  and (_17329_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or (_26935_, _17329_, _17327_);
  and (_17330_, _06290_, _23635_);
  and (_17331_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or (_08819_, _17331_, _17330_);
  and (_17332_, _06290_, _23982_);
  and (_17333_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  or (_08821_, _17333_, _17332_);
  and (_17334_, _24117_, _23806_);
  and (_17335_, _17334_, _23635_);
  not (_17336_, _17334_);
  and (_17337_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_08842_, _17337_, _17335_);
  and (_17338_, _17334_, _23718_);
  and (_17339_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_08844_, _17339_, _17338_);
  and (_17340_, _02444_, _23982_);
  and (_17341_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_08849_, _17341_, _17340_);
  and (_17342_, _02937_, _23718_);
  and (_17343_, _02939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or (_08878_, _17343_, _17342_);
  and (_17344_, _13706_, _23755_);
  and (_17345_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or (_08884_, _17345_, _17344_);
  and (_17346_, _16889_, _23755_);
  and (_17347_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_08888_, _17347_, _17346_);
  and (_17348_, _23806_, _23641_);
  and (_17349_, _17348_, _23589_);
  not (_17350_, _17348_);
  and (_17351_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or (_08904_, _17351_, _17349_);
  and (_17352_, _17348_, _23838_);
  and (_17353_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or (_08907_, _17353_, _17352_);
  and (_17354_, _23863_, _23806_);
  and (_17355_, _17354_, _23982_);
  not (_17356_, _17354_);
  and (_17357_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or (_08914_, _17357_, _17355_);
  and (_17358_, _24103_, _23806_);
  and (_17359_, _17358_, _23635_);
  not (_17360_, _17358_);
  and (_17361_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_08917_, _17361_, _17359_);
  and (_17362_, _17358_, _23676_);
  and (_17363_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_08921_, _17363_, _17362_);
  and (_17364_, _15873_, _23676_);
  and (_17365_, _15875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or (_08923_, _17365_, _17364_);
  and (_17366_, _23962_, _23806_);
  and (_17367_, _17366_, _23838_);
  not (_17368_, _17366_);
  and (_17369_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or (_08927_, _17369_, _17367_);
  not (_17370_, _24017_);
  and (_17371_, _17370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  or (_17372_, _17371_, _24055_);
  and (_17373_, _17372_, _24053_);
  not (_17374_, _17371_);
  nand (_17375_, _17374_, _24027_);
  and (_17376_, _17375_, _23998_);
  or (_17377_, _17371_, _24026_);
  and (_17378_, _17377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_17379_, _17378_, _17376_);
  or (_17380_, _17379_, _17373_);
  and (_17381_, _17380_, _22761_);
  nor (_17382_, _23994_, _23988_);
  and (_08935_, _17382_, _17381_);
  and (_17383_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  and (_17384_, _13764_, _23589_);
  or (_08937_, _17384_, _17383_);
  and (_17385_, _24567_, _23718_);
  and (_17386_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or (_08939_, _17386_, _17385_);
  and (_17387_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  and (_17388_, _13764_, _23755_);
  or (_08941_, _17388_, _17387_);
  and (_17389_, _24078_, _23806_);
  and (_17390_, _17389_, _23755_);
  not (_17391_, _17389_);
  and (_17392_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or (_08951_, _17392_, _17390_);
  and (_17393_, _17389_, _23838_);
  and (_17394_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or (_08954_, _17394_, _17393_);
  and (_17395_, _17389_, _23676_);
  and (_17396_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or (_08956_, _17396_, _17395_);
  and (_17397_, _23806_, _23649_);
  and (_17398_, _17397_, _23589_);
  not (_17399_, _17397_);
  and (_17400_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_08959_, _17400_, _17398_);
  and (_17401_, _17397_, _23635_);
  and (_17402_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_08961_, _17402_, _17401_);
  and (_17403_, _17397_, _23718_);
  and (_17404_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_08965_, _17404_, _17403_);
  and (_17405_, _24547_, _23589_);
  and (_17406_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_08968_, _17406_, _17405_);
  and (_17407_, _23806_, _23594_);
  and (_17408_, _17407_, _23982_);
  not (_17409_, _17407_);
  and (_17410_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_08973_, _17410_, _17408_);
  and (_17411_, _17407_, _23718_);
  and (_17412_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_08976_, _17412_, _17411_);
  and (_17413_, _03277_, _23791_);
  and (_17414_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  or (_08985_, _17414_, _17413_);
  and (_17415_, _16099_, _23676_);
  and (_17416_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  or (_08989_, _17416_, _17415_);
  and (_17417_, _24769_, _23718_);
  and (_17418_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or (_09018_, _17418_, _17417_);
  nor (_26896_[6], _00061_, rst);
  and (_17419_, _02225_, _23982_);
  and (_17420_, _02227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_09027_, _17420_, _17419_);
  and (_17421_, _17366_, _23589_);
  and (_17422_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or (_09051_, _17422_, _17421_);
  and (_17423_, _16483_, _23838_);
  and (_17424_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or (_09053_, _17424_, _17423_);
  and (_17425_, _17312_, _23676_);
  and (_17426_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_09056_, _17426_, _17425_);
  and (_17427_, _17316_, _23718_);
  and (_17428_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_26936_, _17428_, _17427_);
  and (_17429_, _17326_, _23791_);
  and (_17430_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or (_09062_, _17430_, _17429_);
  and (_17431_, _17348_, _23676_);
  and (_17432_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or (_26929_, _17432_, _17431_);
  and (_17433_, _17354_, _23791_);
  and (_17434_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or (_09067_, _17434_, _17433_);
  and (_17435_, _15877_, _23589_);
  and (_17436_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_09069_, _17436_, _17435_);
  and (_17437_, _03277_, _23676_);
  and (_17438_, _03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  or (_09071_, _17438_, _17437_);
  and (_17439_, _17358_, _23718_);
  and (_17440_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_09076_, _17440_, _17439_);
  and (_17441_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_17442_, _17441_, _26153_);
  and (_17443_, _17441_, _26153_);
  or (_17444_, _17443_, _17442_);
  and (_09083_, _17444_, _22761_);
  and (_09091_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _22761_);
  and (_09094_, _00843_, _22761_);
  and (_09097_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _22761_);
  or (_17445_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_17446_, _17441_, rst);
  and (_09101_, _17446_, _17445_);
  and (_17447_, _16513_, _23791_);
  and (_17448_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_09106_, _17448_, _17447_);
  and (_17449_, _16513_, _23676_);
  and (_17450_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_09109_, _17450_, _17449_);
  and (_17451_, _17407_, _23755_);
  and (_17452_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_09112_, _17452_, _17451_);
  and (_17453_, _17312_, _23982_);
  and (_17454_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_09115_, _17454_, _17453_);
  and (_17455_, _17326_, _23589_);
  and (_17456_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_09118_, _17456_, _17455_);
  and (_17457_, _17334_, _23838_);
  and (_17458_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_26931_, _17458_, _17457_);
  and (_17459_, _17348_, _23982_);
  and (_17460_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or (_09122_, _17460_, _17459_);
  and (_17461_, _17358_, _23755_);
  and (_17462_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_09126_, _17462_, _17461_);
  and (_17463_, _17389_, _23791_);
  and (_17464_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or (_09130_, _17464_, _17463_);
  and (_17465_, _17354_, _23635_);
  and (_17466_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or (_09137_, _17466_, _17465_);
  and (_17467_, _16483_, _23635_);
  and (_17468_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or (_09140_, _17468_, _17467_);
  and (_17469_, _17407_, _23589_);
  and (_17470_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_09142_, _17470_, _17469_);
  and (_17471_, _16483_, _23589_);
  and (_17472_, _16485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or (_09148_, _17472_, _17471_);
  and (_17473_, _25536_, _23635_);
  and (_17474_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_09150_, _17474_, _17473_);
  and (_17475_, _06290_, _23676_);
  and (_17476_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or (_09152_, _17476_, _17475_);
  and (_17477_, _16099_, _23838_);
  and (_17478_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or (_09155_, _17478_, _17477_);
  and (_17479_, _17366_, _23755_);
  and (_17480_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or (_27316_, _17480_, _17479_);
  and (_17481_, _16099_, _23718_);
  and (_17482_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or (_09159_, _17482_, _17481_);
  and (_17483_, _16099_, _23791_);
  and (_17484_, _16101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or (_27000_, _17484_, _17483_);
  and (_17485_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_17486_, _09515_, _23589_);
  or (_09194_, _17486_, _17485_);
  and (_17487_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_17488_, _09515_, _23755_);
  or (_09198_, _17488_, _17487_);
  and (_17489_, _16889_, _23791_);
  and (_17490_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_09202_, _17490_, _17489_);
  and (_17491_, _16889_, _23676_);
  and (_17492_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_09205_, _17492_, _17491_);
  and (_17493_, _25536_, _23791_);
  and (_17494_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_09233_, _17494_, _17493_);
  and (_17495_, _02845_, _23589_);
  and (_17496_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_09235_, _17496_, _17495_);
  and (_17497_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  and (_17498_, _13764_, _23791_);
  or (_27104_, _17498_, _17497_);
  and (_17499_, _16889_, _23982_);
  and (_17500_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_09251_, _17500_, _17499_);
  and (_17501_, _13765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and (_17502_, _13764_, _23676_);
  or (_09271_, _17502_, _17501_);
  and (_17503_, _16889_, _23838_);
  and (_17504_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_09281_, _17504_, _17503_);
  and (_17505_, _24577_, _23589_);
  and (_17506_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_09283_, _17506_, _17505_);
  and (_17507_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_17508_, _09515_, _23791_);
  or (_09329_, _17508_, _17507_);
  and (_17509_, _24104_, _23635_);
  and (_17510_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or (_09341_, _17510_, _17509_);
  and (_17511_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and (_17512_, _09515_, _23676_);
  or (_09362_, _17512_, _17511_);
  and (_17513_, _24104_, _23982_);
  and (_17514_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or (_09366_, _17514_, _17513_);
  and (_17515_, _02779_, _23589_);
  and (_17516_, _02781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_09392_, _17516_, _17515_);
  and (_17517_, _13706_, _23635_);
  and (_17518_, _13708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or (_09406_, _17518_, _17517_);
  and (_17519_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_17520_, _09519_, _23589_);
  or (_09421_, _17520_, _17519_);
  and (_17521_, _15503_, _23676_);
  and (_17522_, _15505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_09439_, _17522_, _17521_);
  and (_17523_, _24542_, _23589_);
  and (_17524_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or (_09529_, _17524_, _17523_);
  and (_17525_, _24104_, _23589_);
  and (_17526_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_09546_, _17526_, _17525_);
  and (_17527_, _24597_, _23635_);
  and (_17528_, _24599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or (_09562_, _17528_, _17527_);
  and (_17529_, _24542_, _23755_);
  and (_17530_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or (_09565_, _17530_, _17529_);
  and (_17531_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  and (_17532_, _03641_, _23635_);
  or (_09583_, _17532_, _17531_);
  and (_17533_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_17534_, _09168_, _23791_);
  or (_09616_, _17534_, _17533_);
  and (_17535_, _09169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_17536_, _09168_, _23676_);
  or (_09632_, _17536_, _17535_);
  and (_17537_, _16388_, _23838_);
  and (_17538_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_09668_, _17538_, _17537_);
  and (_17539_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_17540_, _09515_, _23982_);
  or (_09701_, _17540_, _17539_);
  and (_17541_, _16388_, _23718_);
  and (_17542_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_09706_, _17542_, _17541_);
  and (_17543_, _23838_, _23644_);
  and (_17544_, _23646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_09719_, _17544_, _17543_);
  and (_17545_, _17112_, _23755_);
  and (_17546_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_09725_, _17546_, _17545_);
  and (_17547_, _25536_, _23838_);
  and (_17548_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_09729_, _17548_, _17547_);
  and (_17549_, _17366_, _23982_);
  and (_17550_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or (_09731_, _17550_, _17549_);
  and (_17551_, _24670_, _23875_);
  nand (_17552_, _17551_, _23925_);
  and (_17553_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_17554_, _15861_, _23879_);
  and (_17555_, _17554_, _22856_);
  and (_17556_, _17555_, _00708_);
  or (_17557_, _17556_, _17553_);
  or (_17558_, _17557_, _04353_);
  not (_17559_, _04353_);
  or (_17560_, _17559_, _01300_);
  and (_17561_, _17560_, _22761_);
  and (_09740_, _17561_, _17558_);
  and (_17562_, _25400_, _23635_);
  and (_17563_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_09746_, _17563_, _17562_);
  and (_17564_, _17112_, _23838_);
  and (_17565_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_09752_, _17565_, _17564_);
  and (_17566_, _25400_, _23838_);
  and (_17567_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_09754_, _17567_, _17566_);
  and (_17568_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_17569_, _17555_, _00874_);
  or (_17570_, _17569_, _17568_);
  or (_17571_, _17570_, _04353_);
  or (_17572_, _17559_, _03869_);
  and (_17573_, _17572_, _22761_);
  and (_09762_, _17573_, _17571_);
  and (_17574_, _17366_, _23635_);
  and (_17575_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or (_27315_, _17575_, _17574_);
  and (_17576_, _17112_, _23635_);
  and (_17577_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_09767_, _17577_, _17576_);
  and (_17578_, _17551_, _23992_);
  nor (_17579_, _17578_, _04353_);
  or (_17580_, _17579_, _26568_);
  not (_17581_, _17579_);
  or (_17582_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_17583_, _17582_, _22761_);
  and (_09776_, _17583_, _17580_);
  and (_17584_, _16388_, _23791_);
  and (_17585_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_09781_, _17585_, _17584_);
  and (_17586_, _06290_, _23791_);
  and (_17587_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or (_09788_, _17587_, _17586_);
  and (_17588_, _16037_, _23635_);
  and (_17589_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_09791_, _17589_, _17588_);
  and (_17590_, _17407_, _23676_);
  and (_17591_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_09798_, _17591_, _17590_);
  or (_17592_, _17579_, _00580_);
  or (_17593_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_17594_, _17593_, _22761_);
  and (_09806_, _17594_, _17592_);
  and (_17595_, _17104_, _23676_);
  and (_17596_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or (_09811_, _17596_, _17595_);
  and (_17597_, _16037_, _23755_);
  and (_17598_, _16039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_09816_, _17598_, _17597_);
  and (_17599_, _16475_, _23676_);
  and (_17600_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or (_09818_, _17600_, _17599_);
  and (_17601_, _25536_, _23589_);
  and (_17602_, _25538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_09821_, _17602_, _17601_);
  and (_17603_, _03354_, _23676_);
  and (_17604_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_09823_, _17604_, _17603_);
  and (_17605_, _17104_, _23791_);
  and (_17606_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or (_09835_, _17606_, _17605_);
  and (_17607_, _23982_, _23601_);
  and (_17608_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or (_09838_, _17608_, _17607_);
  and (_17609_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_17610_, _17609_, _03826_);
  and (_17611_, _17610_, _00310_);
  or (_17612_, _00311_, _00310_);
  nor (_17613_, _17612_, _23522_);
  and (_17614_, _00313_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_17615_, _17614_, _25771_);
  or (_17616_, _17615_, _17613_);
  or (_17617_, _17616_, _17611_);
  nand (_17618_, _25775_, _23585_);
  and (_17619_, _17618_, _22761_);
  and (_09841_, _17619_, _17617_);
  and (_17620_, _17407_, _23791_);
  and (_17621_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_09847_, _17621_, _17620_);
  nand (_17622_, _17581_, _00791_);
  or (_17623_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_17624_, _17623_, _22761_);
  and (_09852_, _17624_, _17622_);
  or (_17625_, _17579_, _00484_);
  or (_17626_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_17627_, _17626_, _22761_);
  and (_09854_, _17627_, _17625_);
  and (_17628_, _16475_, _23791_);
  and (_17629_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or (_09861_, _17629_, _17628_);
  and (_17630_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_17631_, _17555_, _00647_);
  or (_17632_, _17631_, _17630_);
  or (_17633_, _17632_, _04353_);
  or (_17634_, _17559_, _01228_);
  and (_17635_, _17634_, _22761_);
  and (_09879_, _17635_, _17633_);
  and (_17636_, _17407_, _23838_);
  and (_17637_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_09889_, _17637_, _17636_);
  and (_17638_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_17639_, _17555_, _00580_);
  or (_17640_, _17639_, _17638_);
  or (_17641_, _17640_, _04353_);
  nand (_17642_, _04353_, _01138_);
  and (_17643_, _17642_, _22761_);
  and (_09892_, _17643_, _17641_);
  and (_17644_, _17104_, _23718_);
  and (_17645_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or (_09894_, _17645_, _17644_);
  and (_17646_, _23755_, _23601_);
  and (_17647_, _23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or (_09897_, _17647_, _17646_);
  and (_17648_, _17407_, _23635_);
  and (_17649_, _17409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_09900_, _17649_, _17648_);
  and (_17650_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_17651_, _17555_, _00484_);
  or (_17652_, _17651_, _17650_);
  or (_17653_, _17652_, _04353_);
  nand (_17654_, _04353_, _01071_);
  and (_17655_, _17654_, _22761_);
  and (_09907_, _17655_, _17653_);
  and (_17656_, _17104_, _23982_);
  and (_17657_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or (_09912_, _17657_, _17656_);
  and (_17658_, _23982_, _23811_);
  and (_17659_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or (_09920_, _17659_, _17658_);
  and (_17660_, _02459_, _23791_);
  and (_17661_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or (_09922_, _17661_, _17660_);
  and (_17662_, _24547_, _23755_);
  and (_17663_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_09925_, _17663_, _17662_);
  or (_17664_, _17579_, _00408_);
  or (_17665_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_17666_, _17665_, _22761_);
  and (_09932_, _17666_, _17664_);
  or (_17667_, _17579_, _00708_);
  or (_17668_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_17669_, _17668_, _22761_);
  and (_09935_, _17669_, _17667_);
  or (_17670_, _17579_, _00647_);
  or (_17671_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_17672_, _17671_, _22761_);
  and (_09937_, _17672_, _17670_);
  and (_17673_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_17674_, _17555_, _00408_);
  or (_17675_, _17674_, _17673_);
  or (_17676_, _17675_, _04353_);
  nand (_17677_, _04353_, _01011_);
  and (_17678_, _17677_, _22761_);
  and (_09939_, _17678_, _17676_);
  and (_17679_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_17680_, _17555_, _26568_);
  or (_17681_, _17680_, _17679_);
  or (_17682_, _17681_, _04353_);
  nand (_17683_, _04353_, _00950_);
  and (_17684_, _17683_, _22761_);
  and (_09941_, _17684_, _17682_);
  and (_17685_, _15877_, _23718_);
  and (_17686_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_09947_, _17686_, _17685_);
  or (_17687_, _17579_, _00874_);
  or (_17688_, _17581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_17689_, _17688_, _22761_);
  and (_09950_, _17689_, _17687_);
  and (_17690_, _23811_, _23635_);
  and (_17691_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or (_09959_, _17691_, _17690_);
  and (_17692_, _15877_, _23791_);
  and (_17693_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_26997_, _17693_, _17692_);
  and (_17694_, _02459_, _23838_);
  and (_17695_, _02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or (_09963_, _17695_, _17694_);
  and (_17696_, _23811_, _23589_);
  and (_17697_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_09969_, _17697_, _17696_);
  and (_17698_, _17397_, _23676_);
  and (_17699_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_27312_, _17699_, _17698_);
  and (_17700_, _17086_, _23676_);
  and (_17701_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or (_09978_, _17701_, _17700_);
  nor (_17702_, _17552_, _00791_);
  and (_17703_, _17552_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_17704_, _17703_, _04353_);
  or (_17705_, _17704_, _17702_);
  nand (_17706_, _04353_, _01377_);
  and (_17707_, _17706_, _22761_);
  and (_09981_, _17707_, _17705_);
  and (_17709_, _17397_, _23791_);
  and (_17710_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_09983_, _17710_, _17709_);
  and (_17711_, _24104_, _23755_);
  and (_17712_, _24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or (_27244_, _17712_, _17711_);
  and (_17713_, _06290_, _23718_);
  and (_17714_, _06293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or (_09988_, _17714_, _17713_);
  and (_17715_, _17397_, _23838_);
  and (_17716_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_27313_, _17716_, _17715_);
  and (_17717_, _17086_, _23791_);
  and (_17718_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or (_09995_, _17718_, _17717_);
  and (_17719_, _02379_, _23791_);
  and (_17720_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_09997_, _17720_, _17719_);
  nand (_17721_, _23927_, _23748_);
  nor (_17722_, _24156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_17723_, _17722_, _24158_);
  and (_17724_, _17723_, _24150_);
  and (_17725_, _24152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_17726_, _15456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_17727_, _17726_, _23921_);
  or (_17728_, _17727_, _17725_);
  or (_17729_, _17728_, _17724_);
  or (_17730_, _17729_, _23927_);
  and (_17731_, _17730_, _22761_);
  and (_10001_, _17731_, _17721_);
  and (_17732_, _15877_, _23838_);
  and (_17733_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_10008_, _17733_, _17732_);
  and (_17734_, _17397_, _23982_);
  and (_17735_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_10019_, _17735_, _17734_);
  and (_17736_, _15877_, _23635_);
  and (_17737_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_26999_, _17737_, _17736_);
  and (_17738_, _17086_, _23718_);
  and (_17739_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or (_27297_, _17739_, _17738_);
  and (_17740_, _02379_, _23755_);
  and (_17741_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_10025_, _17741_, _17740_);
  and (_17742_, _17001_, _23838_);
  and (_17743_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or (_10030_, _17743_, _17742_);
  and (_17744_, _17397_, _23755_);
  and (_17745_, _17399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_10034_, _17745_, _17744_);
  and (_17746_, _17086_, _23982_);
  and (_17747_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or (_10036_, _17747_, _17746_);
  and (_17748_, _17001_, _23718_);
  and (_17749_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or (_10038_, _17749_, _17748_);
  and (_17750_, _17086_, _23755_);
  and (_17751_, _17088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or (_27298_, _17751_, _17750_);
  and (_17752_, _17001_, _23589_);
  and (_17753_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or (_10046_, _17753_, _17752_);
  and (_17754_, _15877_, _23982_);
  and (_17755_, _15879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_26998_, _17755_, _17754_);
  and (_17756_, _17078_, _23676_);
  and (_17757_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_10066_, _17757_, _17756_);
  and (_17758_, _24577_, _23982_);
  and (_17759_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or (_10070_, _17759_, _17758_);
  and (_17760_, _17389_, _23718_);
  and (_17761_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or (_10073_, _17761_, _17760_);
  and (_17762_, _17389_, _23982_);
  and (_17763_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or (_10080_, _17763_, _17762_);
  and (_17764_, _02877_, _23676_);
  and (_17765_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_10089_, _17765_, _17764_);
  and (_17766_, _17078_, _23791_);
  and (_17767_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_10092_, _17767_, _17766_);
  and (_17768_, _17078_, _23838_);
  and (_17769_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_27299_, _17769_, _17768_);
  and (_17770_, _17389_, _23635_);
  and (_17771_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or (_27314_, _17771_, _17770_);
  and (_17772_, _02877_, _23838_);
  and (_17773_, _02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_10105_, _17773_, _17772_);
  and (_17774_, _17389_, _23589_);
  and (_17775_, _17391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_10110_, _17775_, _17774_);
  and (_17776_, _06044_, _23838_);
  and (_17777_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_27234_, _17777_, _17776_);
  and (_17778_, _17078_, _23982_);
  and (_17779_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_27300_, _17779_, _17778_);
  and (_17780_, _06044_, _23676_);
  and (_17781_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_10120_, _17781_, _17780_);
  and (_17782_, _00310_, _23986_);
  nand (_17783_, _17782_, _23522_);
  or (_17784_, _17782_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_17785_, _17784_, _25776_);
  and (_17786_, _17785_, _17783_);
  or (_17787_, _17786_, _25914_);
  and (_10124_, _17787_, _22761_);
  and (_17788_, _24777_, _23791_);
  and (_17789_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or (_10127_, _17789_, _17788_);
  and (_17790_, _17078_, _23755_);
  and (_17791_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_10136_, _17791_, _17790_);
  and (_17792_, _06044_, _23589_);
  and (_17793_, _06046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_10138_, _17793_, _17792_);
  and (_17794_, _03281_, _23982_);
  and (_17795_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_10141_, _17795_, _17794_);
  and (_17796_, _00310_, _23925_);
  nand (_17797_, _17796_, _23522_);
  or (_17798_, _17796_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_17799_, _17798_, _25772_);
  and (_17800_, _17799_, _17797_);
  or (_17801_, _17800_, _25777_);
  and (_10143_, _17801_, _22761_);
  and (_17802_, _00310_, _23919_);
  and (_17803_, _17802_, _23522_);
  nor (_17804_, _17802_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_17805_, _17804_, _17803_);
  nand (_17806_, _17805_, _25776_);
  nand (_17807_, _25775_, _23628_);
  and (_17808_, _17807_, _22761_);
  and (_10145_, _17808_, _17806_);
  and (_17809_, _15967_, _23589_);
  and (_17810_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_10150_, _17810_, _17809_);
  or (_17811_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_17812_, _00378_, _26546_);
  or (_17813_, _17812_, _00461_);
  or (_17814_, _17813_, _00553_);
  or (_17815_, _17814_, _00625_);
  or (_17816_, _17815_, _00682_);
  and (_17817_, _17816_, _23531_);
  and (_17818_, _23455_, _23402_);
  not (_17819_, _23455_);
  and (_17820_, _23457_, _17819_);
  or (_17821_, _17820_, _17818_);
  and (_17822_, _17821_, _23398_);
  nand (_17823_, _23386_, _23092_);
  or (_17824_, _23387_, _23386_);
  and (_17825_, _17824_, _23037_);
  and (_17826_, _17825_, _17823_);
  and (_17827_, _23528_, _23404_);
  and (_17828_, _17827_, _23278_);
  and (_17829_, _01121_, _26151_);
  and (_17830_, _17829_, _01278_);
  nand (_17831_, _17830_, _17828_);
  nand (_17832_, _17831_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_17833_, _17832_, _17826_);
  nor (_17834_, _17833_, _17822_);
  nand (_17835_, _17834_, _00767_);
  or (_17836_, _17835_, _17817_);
  or (_17837_, _17836_, _00850_);
  and (_17838_, _17837_, _17811_);
  or (_17839_, _17838_, _00310_);
  not (_17840_, _00310_);
  and (_17841_, _02508_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_17842_, _17841_, _02509_);
  or (_17843_, _17842_, _17840_);
  and (_17844_, _17843_, _17839_);
  or (_17845_, _17844_, _25775_);
  or (_17846_, _25776_, _23709_);
  and (_17847_, _17846_, _22761_);
  and (_10155_, _17847_, _17845_);
  or (_17848_, _24688_, _00569_);
  nand (_17849_, _17848_, _00310_);
  or (_17850_, _17849_, _03810_);
  and (_17851_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_17852_, _17851_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_17853_, _23451_, _23398_);
  and (_17854_, _23345_, _23037_);
  nand (_17855_, _23494_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_17856_, _17855_, _17851_);
  or (_17857_, _17856_, _17854_);
  or (_17858_, _17857_, _17853_);
  and (_17859_, _17858_, _17852_);
  or (_17860_, _17859_, _00310_);
  and (_17861_, _17860_, _17850_);
  or (_17862_, _17861_, _25775_);
  nand (_17863_, _25775_, _23748_);
  and (_17864_, _17863_, _22761_);
  and (_10158_, _17864_, _17862_);
  and (_17865_, _24777_, _23589_);
  and (_17866_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_10160_, _17866_, _17865_);
  and (_17867_, _17366_, _23676_);
  and (_17868_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or (_10162_, _17868_, _17867_);
  and (_17869_, _17112_, _23791_);
  and (_17870_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_10168_, _17870_, _17869_);
  and (_17871_, _17366_, _23791_);
  and (_17872_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or (_10172_, _17872_, _17871_);
  and (_17873_, _03234_, _23676_);
  and (_17874_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  or (_10175_, _17874_, _17873_);
  and (_10177_, _03872_, _22761_);
  and (_17875_, _00310_, _23878_);
  and (_17876_, _17875_, _23522_);
  nor (_17877_, _17875_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_17878_, _17877_, _17876_);
  nand (_17879_, _17878_, _25776_);
  nand (_17880_, _25775_, _23784_);
  and (_17881_, _17880_, _22761_);
  and (_10185_, _17881_, _17879_);
  and (_17882_, _17112_, _23718_);
  and (_17883_, _17114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_27301_, _17883_, _17882_);
  and (_17884_, _17366_, _23718_);
  and (_17885_, _17368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or (_10193_, _17885_, _17884_);
  and (_17886_, _17104_, _23755_);
  and (_17887_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or (_27302_, _17887_, _17886_);
  and (_17888_, _17358_, _23791_);
  and (_17889_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_10203_, _17889_, _17888_);
  and (_17890_, _17104_, _23589_);
  and (_17891_, _17106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or (_10209_, _17891_, _17890_);
  and (_17892_, _16889_, _23718_);
  and (_17893_, _16891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_10213_, _17893_, _17892_);
  and (_17894_, _17358_, _23838_);
  and (_17895_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_10216_, _17895_, _17894_);
  and (_17896_, _16513_, _23718_);
  and (_17897_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_10219_, _17897_, _17896_);
  and (_17898_, _17070_, _23676_);
  and (_17899_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_10223_, _17899_, _17898_);
  and (_17900_, _17070_, _23718_);
  and (_17901_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_10226_, _17901_, _17900_);
  and (_17902_, _03234_, _23838_);
  and (_17903_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  or (_10231_, _17903_, _17902_);
  and (_17904_, _03281_, _23755_);
  and (_17905_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_10233_, _17905_, _17904_);
  and (_17906_, _16513_, _23589_);
  and (_17907_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_27248_, _17907_, _17906_);
  and (_17908_, _17358_, _23982_);
  and (_17909_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_26925_, _17909_, _17908_);
  and (_17910_, _16513_, _23635_);
  and (_17911_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_27247_, _17911_, _17910_);
  and (_17912_, _17358_, _23589_);
  and (_17913_, _17360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_26926_, _17913_, _17912_);
  and (_17914_, _03234_, _23718_);
  and (_17915_, _03236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or (_26987_, _17915_, _17914_);
  and (_17916_, _17070_, _23838_);
  and (_17917_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_27303_, _17917_, _17916_);
  nor (_10263_, _03823_, rst);
  and (_17918_, _07101_, _23635_);
  and (_17919_, _07103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or (_10268_, _17919_, _17918_);
  and (_17920_, _17354_, _23676_);
  and (_17921_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or (_10302_, _17921_, _17920_);
  nor (_10307_, _03759_, rst);
  and (_17922_, _04692_, _23838_);
  and (_17923_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_10328_, _17923_, _17922_);
  and (_17924_, _17070_, _23982_);
  and (_17925_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_10332_, _17925_, _17924_);
  and (_17926_, _04692_, _23676_);
  and (_17927_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_10348_, _17927_, _17926_);
  and (_10355_, _03773_, _22761_);
  and (_17928_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  and (_17929_, _13826_, _23589_);
  or (_10368_, _17929_, _17928_);
  nor (_26906_[6], _00812_, rst);
  and (_17930_, _17354_, _23718_);
  and (_17931_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or (_10374_, _17931_, _17930_);
  and (_10380_, _03803_, _22761_);
  and (_17932_, _17070_, _23755_);
  and (_17933_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_10391_, _17933_, _17932_);
  and (_10414_, _03792_, _22761_);
  and (_17934_, _03015_, _23755_);
  and (_17935_, _03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_10418_, _17935_, _17934_);
  and (_17936_, _04692_, _23589_);
  and (_17937_, _04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_10437_, _17937_, _17936_);
  and (_17938_, _16388_, _23982_);
  and (_17939_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_10442_, _17939_, _17938_);
  and (_17940_, _16475_, _23982_);
  and (_17941_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or (_10451_, _17941_, _17940_);
  and (_17942_, _17070_, _23589_);
  and (_17943_, _17072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_10453_, _17943_, _17942_);
  and (_17944_, _17354_, _23838_);
  and (_17945_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or (_10460_, _17945_, _17944_);
  and (_17946_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_17947_, _09515_, _23838_);
  or (_27103_, _17947_, _17946_);
  and (_17948_, _03001_, _23838_);
  and (_17949_, _03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or (_10490_, _17949_, _17948_);
  and (_17950_, _15967_, _23718_);
  and (_17951_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_26985_, _17951_, _17950_);
  and (_17952_, _17354_, _23755_);
  and (_17953_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or (_26927_, _17953_, _17952_);
  and (_10500_, _03743_, _22761_);
  and (_17954_, _17064_, _23676_);
  and (_17955_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or (_10504_, _17955_, _17954_);
  and (_17956_, _15967_, _23838_);
  and (_17957_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_10507_, _17957_, _17956_);
  and (_10511_, _03730_, _22761_);
  and (_17958_, _02322_, _23791_);
  and (_17959_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_10523_, _17959_, _17958_);
  and (_17960_, _09516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_17961_, _09515_, _23718_);
  or (_10528_, _17961_, _17960_);
  and (_17962_, _17354_, _23589_);
  and (_17963_, _17356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_26928_, _17963_, _17962_);
  and (_17964_, _17064_, _23791_);
  and (_17965_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or (_27304_, _17965_, _17964_);
  and (_17966_, _24769_, _23589_);
  and (_17967_, _24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or (_10536_, _17967_, _17966_);
  and (_17968_, _03281_, _23676_);
  and (_17969_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_27179_, _17969_, _17968_);
  and (_17970_, _17348_, _23791_);
  and (_17971_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or (_10546_, _17971_, _17970_);
  and (_17972_, _23842_, _23599_);
  and (_17973_, _17972_, _23982_);
  not (_17974_, _17972_);
  and (_17975_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_10554_, _17975_, _17973_);
  and (_17976_, _17064_, _23838_);
  and (_17977_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or (_10561_, _17977_, _17976_);
  and (_17978_, _23649_, _23599_);
  not (_17979_, _17978_);
  and (_17980_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_17981_, _17978_, _23755_);
  or (_10567_, _17981_, _17980_);
  and (_17982_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  and (_17983_, _13838_, _23791_);
  or (_10569_, _17983_, _17982_);
  and (_17984_, _17064_, _23635_);
  and (_17985_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or (_10576_, _17985_, _17984_);
  and (_17986_, _17348_, _23718_);
  and (_17987_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or (_10579_, _17987_, _17986_);
  and (_17988_, _17348_, _23635_);
  and (_17989_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or (_10586_, _17989_, _17988_);
  and (_17990_, _23849_, _23599_);
  and (_17991_, _17990_, _23982_);
  not (_17992_, _17990_);
  and (_17993_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or (_10592_, _17993_, _17991_);
  and (_17994_, _17990_, _23838_);
  and (_17995_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or (_27258_, _17995_, _17994_);
  and (_17996_, _17990_, _23635_);
  and (_17997_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or (_27259_, _17997_, _17996_);
  and (_17998_, _13839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  and (_17999_, _13838_, _23718_);
  or (_10607_, _17999_, _17998_);
  and (_18000_, _17064_, _23589_);
  and (_18001_, _17066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or (_10609_, _18001_, _18000_);
  and (_18002_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_18003_, _17978_, _23635_);
  or (_10611_, _18003_, _18002_);
  and (_18004_, _03643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  and (_18005_, _03641_, _23982_);
  or (_10616_, _18005_, _18004_);
  and (_18006_, _17348_, _23755_);
  and (_18007_, _17350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or (_10622_, _18007_, _18006_);
  and (_18008_, _17058_, _23676_);
  and (_18009_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or (_10628_, _18009_, _18008_);
  and (_18010_, _17990_, _23755_);
  and (_18011_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or (_10630_, _18011_, _18010_);
  and (_18012_, _17334_, _23676_);
  and (_18013_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_26930_, _18013_, _18012_);
  and (_18014_, _16388_, _23635_);
  and (_18015_, _16390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_10639_, _18015_, _18014_);
  and (_18016_, _17058_, _23718_);
  and (_18017_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or (_27306_, _18017_, _18016_);
  and (_18018_, _16475_, _23635_);
  and (_18019_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or (_10650_, _18019_, _18018_);
  and (_18020_, _17058_, _23982_);
  and (_18021_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or (_10653_, _18021_, _18020_);
  and (_18022_, _16475_, _23589_);
  and (_18023_, _16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or (_10656_, _18023_, _18022_);
  and (_18024_, _17334_, _23791_);
  and (_18025_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_10669_, _18025_, _18024_);
  and (_18026_, _12505_, _23791_);
  and (_18027_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_10673_, _18027_, _18026_);
  and (_18028_, _17334_, _23982_);
  and (_18029_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_10676_, _18029_, _18028_);
  and (_18031_, _17058_, _23589_);
  and (_18032_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or (_10679_, _18032_, _18031_);
  and (_18033_, _17334_, _23755_);
  and (_18034_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_26932_, _18034_, _18033_);
  and (_18035_, _12505_, _23589_);
  and (_18036_, _12508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or (_10688_, _18036_, _18035_);
  and (_18037_, _17050_, _23676_);
  and (_18038_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_27307_, _18038_, _18037_);
  and (_18039_, _17990_, _23589_);
  and (_18040_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or (_27260_, _18040_, _18039_);
  and (_18041_, _06081_, _23635_);
  and (_18042_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or (_10710_, _18042_, _18041_);
  and (_18043_, _17334_, _23589_);
  and (_18044_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_10713_, _18044_, _18043_);
  and (_18045_, _17050_, _23718_);
  and (_18046_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_10716_, _18046_, _18045_);
  and (_18047_, _06081_, _23718_);
  and (_18048_, _06083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or (_10718_, _18048_, _18047_);
  and (_18049_, _17050_, _23982_);
  and (_18050_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_10721_, _18050_, _18049_);
  and (_18051_, _03046_, _23838_);
  and (_18052_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_10724_, _18052_, _18051_);
  and (_18053_, _17326_, _23676_);
  and (_18054_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or (_10727_, _18054_, _18053_);
  and (_18055_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_18056_, _17978_, _23982_);
  or (_10729_, _18056_, _18055_);
  and (_18057_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  and (_18058_, _13826_, _23838_);
  or (_27113_, _18058_, _18057_);
  and (_18059_, _03046_, _23676_);
  and (_18060_, _03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_27266_, _18060_, _18059_);
  and (_18061_, _17326_, _23718_);
  and (_18062_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or (_10737_, _18062_, _18061_);
  and (_18063_, _12516_, _23791_);
  and (_18064_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or (_10742_, _18064_, _18063_);
  and (_18065_, _25517_, _23838_);
  and (_18066_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_10745_, _18066_, _18065_);
  and (_18067_, _16463_, _23791_);
  and (_18068_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or (_10751_, _18068_, _18067_);
  and (_18069_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  and (_18070_, _13826_, _23718_);
  or (_10754_, _18070_, _18069_);
  and (_18071_, _17050_, _23755_);
  and (_18072_, _17052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_10756_, _18072_, _18071_);
  and (_18073_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  and (_18074_, _13826_, _23791_);
  or (_10758_, _18074_, _18073_);
  and (_18075_, _16463_, _23838_);
  and (_18076_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or (_10762_, _18076_, _18075_);
  and (_18077_, _17326_, _23838_);
  and (_18078_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or (_26933_, _18078_, _18077_);
  and (_18079_, _16463_, _23635_);
  and (_18080_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or (_26955_, _18080_, _18079_);
  and (_18081_, _15967_, _23635_);
  and (_18082_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_26986_, _18082_, _18081_);
  and (_18083_, _25517_, _23755_);
  and (_18084_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_10780_, _18084_, _18083_);
  and (_18085_, _03354_, _23791_);
  and (_18086_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_10782_, _18086_, _18085_);
  and (_18087_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_18088_, _09519_, _23838_);
  or (_10787_, _18088_, _18087_);
  and (_18089_, _17326_, _23982_);
  and (_18090_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or (_10792_, _18090_, _18089_);
  and (_18091_, _25209_, _24671_);
  nand (_18092_, _18091_, _23522_);
  or (_18093_, _18091_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_18094_, _18093_, _24629_);
  and (_18095_, _18094_, _18092_);
  nand (_18096_, _25216_, _23585_);
  or (_18097_, _25216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_18098_, _18097_, _23880_);
  and (_18099_, _18098_, _18096_);
  and (_18100_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_18101_, _18100_, rst);
  or (_18102_, _18101_, _18099_);
  or (_10802_, _18102_, _18095_);
  and (_18103_, _17042_, _23791_);
  and (_18104_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_10807_, _18104_, _18103_);
  and (_18105_, _16463_, _23755_);
  and (_18106_, _16465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or (_10809_, _18106_, _18105_);
  and (_18107_, _17042_, _23838_);
  and (_18108_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_10811_, _18108_, _18107_);
  and (_18109_, _15967_, _23755_);
  and (_18110_, _15969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_10813_, _18110_, _18109_);
  and (_18111_, _16850_, _23635_);
  and (_18112_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or (_10815_, _18112_, _18111_);
  and (_18113_, _02326_, _23589_);
  and (_18114_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or (_10818_, _18114_, _18113_);
  and (_18115_, _17326_, _23635_);
  and (_18116_, _17328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or (_26934_, _18116_, _18115_);
  and (_18117_, _16455_, _23676_);
  and (_18118_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_26957_, _18118_, _18117_);
  and (_18119_, _16455_, _23718_);
  and (_18120_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_10823_, _18120_, _18119_);
  and (_18121_, _17042_, _23635_);
  and (_18122_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_10828_, _18122_, _18121_);
  and (_18123_, _17316_, _23791_);
  and (_18124_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_10830_, _18124_, _18123_);
  and (_18125_, _17042_, _23589_);
  and (_18126_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_10832_, _18126_, _18125_);
  and (_18127_, _16850_, _23589_);
  and (_18128_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or (_10835_, _18128_, _18127_);
  and (_18129_, _24542_, _23718_);
  and (_18130_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or (_10838_, _18130_, _18129_);
  and (_18131_, _17316_, _23838_);
  and (_18132_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_10840_, _18132_, _18131_);
  and (_18133_, _17038_, _23676_);
  and (_18134_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or (_10843_, _18134_, _18133_);
  and (_18135_, _02845_, _23718_);
  and (_18136_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_10845_, _18136_, _18135_);
  and (_18137_, _16455_, _23982_);
  and (_18138_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_26958_, _18138_, _18137_);
  and (_18139_, _03281_, _23718_);
  and (_18140_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_10849_, _18140_, _18139_);
  and (_18141_, _16455_, _23635_);
  and (_18142_, _16457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_26959_, _18142_, _18141_);
  and (_18143_, _17316_, _23982_);
  and (_18144_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_10861_, _18144_, _18143_);
  and (_18145_, _02379_, _23838_);
  and (_18146_, _02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_10866_, _18146_, _18145_);
  and (_18147_, _17038_, _23791_);
  and (_18148_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or (_10869_, _18148_, _18147_);
  and (_18149_, _16850_, _23755_);
  and (_18150_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or (_10872_, _18150_, _18149_);
  and (_18151_, _16447_, _23676_);
  and (_18152_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_10874_, _18152_, _18151_);
  and (_18153_, _17038_, _23982_);
  and (_18154_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or (_10876_, _18154_, _18153_);
  and (_18155_, _16707_, _23589_);
  and (_18156_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_10878_, _18156_, _18155_);
  and (_18157_, _17316_, _23755_);
  and (_18158_, _17318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_10880_, _18158_, _18157_);
  and (_18159_, _16447_, _23718_);
  and (_18160_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_10882_, _18160_, _18159_);
  or (_18161_, _16875_, _05308_);
  and (_18162_, _18161_, _22768_);
  nand (_18163_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_18164_, _18163_, _26823_);
  or (_18165_, _18164_, _18162_);
  and (_26881_[1], _18165_, _22761_);
  and (_18166_, _16447_, _23982_);
  and (_18167_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_10888_, _18167_, _18166_);
  and (_18168_, _17038_, _23635_);
  and (_18169_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_10890_, _18169_, _18168_);
  and (_18170_, _17312_, _23791_);
  and (_18171_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_10895_, _18171_, _18170_);
  and (_18172_, _17038_, _23755_);
  and (_18173_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or (_10897_, _18173_, _18172_);
  and (_18174_, _16447_, _23635_);
  and (_18175_, _16449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_10899_, _18175_, _18174_);
  and (_18176_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_18177_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_18178_, _18177_, _18176_);
  and (_18179_, _18178_, _09527_);
  and (_18180_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_18181_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_18182_, _18181_, _18180_);
  and (_18183_, _18182_, _05352_);
  or (_18184_, _18183_, _18179_);
  or (_18185_, _18184_, _09540_);
  and (_18186_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and (_18187_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_18188_, _18187_, _18186_);
  and (_18189_, _18188_, _09527_);
  and (_18190_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_18191_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_18192_, _18191_, _18190_);
  and (_18193_, _18192_, _05352_);
  or (_18194_, _18193_, _18189_);
  or (_18195_, _18194_, _05373_);
  and (_18196_, _18195_, _09566_);
  and (_18197_, _18196_, _18185_);
  or (_18198_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_18199_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_18200_, _18199_, _18198_);
  and (_18201_, _18200_, _09527_);
  or (_18202_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_18203_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_18204_, _18203_, _18202_);
  and (_18205_, _18204_, _05352_);
  or (_18206_, _18205_, _18201_);
  or (_18207_, _18206_, _09540_);
  or (_18208_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_18209_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_18210_, _18209_, _18208_);
  and (_18211_, _18210_, _09527_);
  or (_18212_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_18213_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and (_18214_, _18213_, _18212_);
  and (_18215_, _18214_, _05352_);
  or (_18216_, _18215_, _18211_);
  or (_18217_, _18216_, _05373_);
  and (_18218_, _18217_, _05379_);
  and (_18219_, _18218_, _18207_);
  or (_18220_, _18219_, _18197_);
  and (_18221_, _18220_, _05361_);
  and (_18222_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_18223_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_18224_, _18223_, _18222_);
  and (_18225_, _18224_, _09527_);
  and (_18226_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_18227_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_18228_, _18227_, _18226_);
  and (_18229_, _18228_, _05352_);
  or (_18230_, _18229_, _18225_);
  or (_18231_, _18230_, _09540_);
  and (_18232_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_18233_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_18234_, _18233_, _18232_);
  and (_18235_, _18234_, _09527_);
  and (_18236_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_18237_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_18238_, _18237_, _18236_);
  and (_18239_, _18238_, _05352_);
  or (_18240_, _18239_, _18235_);
  or (_18241_, _18240_, _05373_);
  and (_18242_, _18241_, _09566_);
  and (_18243_, _18242_, _18231_);
  or (_18244_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_18245_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_18246_, _18245_, _05352_);
  and (_18247_, _18246_, _18244_);
  or (_18248_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_18249_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_18250_, _18249_, _09527_);
  and (_18251_, _18250_, _18248_);
  or (_18252_, _18251_, _18247_);
  or (_18253_, _18252_, _09540_);
  or (_18254_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_18255_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and (_18256_, _18255_, _05352_);
  and (_18257_, _18256_, _18254_);
  or (_18258_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_18259_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and (_18260_, _18259_, _09527_);
  and (_18261_, _18260_, _18258_);
  or (_18262_, _18261_, _18257_);
  or (_18263_, _18262_, _05373_);
  and (_18264_, _18263_, _05379_);
  and (_18265_, _18264_, _18253_);
  or (_18266_, _18265_, _18243_);
  and (_18267_, _18266_, _09581_);
  or (_18268_, _18267_, _18221_);
  and (_18269_, _18268_, _09682_);
  and (_18270_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_18271_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_18272_, _18271_, _18270_);
  and (_18273_, _18272_, _09527_);
  and (_18274_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_18275_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_18276_, _18275_, _18274_);
  and (_18277_, _18276_, _05352_);
  or (_18278_, _18277_, _18273_);
  and (_18279_, _18278_, _05373_);
  and (_18280_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_18281_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_18282_, _18281_, _18280_);
  and (_18283_, _18282_, _09527_);
  and (_18284_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_18285_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_18286_, _18285_, _18284_);
  and (_18287_, _18286_, _05352_);
  or (_18288_, _18287_, _18283_);
  and (_18289_, _18288_, _09540_);
  or (_18290_, _18289_, _18279_);
  and (_18291_, _18290_, _09566_);
  or (_18292_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_18293_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_18294_, _18293_, _05352_);
  and (_18295_, _18294_, _18292_);
  or (_18296_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_18297_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_18298_, _18297_, _09527_);
  and (_18299_, _18298_, _18296_);
  or (_18300_, _18299_, _18295_);
  and (_18301_, _18300_, _05373_);
  or (_18302_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_18303_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_18304_, _18303_, _05352_);
  and (_18305_, _18304_, _18302_);
  or (_18306_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_18307_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_18308_, _18307_, _09527_);
  and (_18309_, _18308_, _18306_);
  or (_18310_, _18309_, _18305_);
  and (_18311_, _18310_, _09540_);
  or (_18312_, _18311_, _18301_);
  and (_18313_, _18312_, _05379_);
  or (_18314_, _18313_, _18291_);
  and (_18315_, _18314_, _09581_);
  and (_18316_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_18317_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_18318_, _18317_, _18316_);
  and (_18319_, _18318_, _09527_);
  and (_18320_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_18321_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_18322_, _18321_, _18320_);
  and (_18323_, _18322_, _05352_);
  or (_18324_, _18323_, _18319_);
  and (_18325_, _18324_, _05373_);
  and (_18326_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and (_18327_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_18328_, _18327_, _18326_);
  and (_18329_, _18328_, _09527_);
  and (_18330_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_18331_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_18332_, _18331_, _18330_);
  and (_18333_, _18332_, _05352_);
  or (_18334_, _18333_, _18329_);
  and (_18335_, _18334_, _09540_);
  or (_18336_, _18335_, _18325_);
  and (_18337_, _18336_, _09566_);
  or (_18338_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_18339_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_18340_, _18339_, _18338_);
  and (_18341_, _18340_, _09527_);
  or (_18342_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_18343_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_18344_, _18343_, _18342_);
  and (_18345_, _18344_, _05352_);
  or (_18346_, _18345_, _18341_);
  and (_18347_, _18346_, _05373_);
  or (_18348_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_18349_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_18350_, _18349_, _18348_);
  and (_18351_, _18350_, _09527_);
  or (_18352_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_18353_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_18354_, _18353_, _18352_);
  and (_18355_, _18354_, _05352_);
  or (_18356_, _18355_, _18351_);
  and (_18357_, _18356_, _09540_);
  or (_18358_, _18357_, _18347_);
  and (_18359_, _18358_, _05379_);
  or (_18360_, _18359_, _18337_);
  and (_18361_, _18360_, _05361_);
  or (_18362_, _18361_, _18315_);
  and (_18363_, _18362_, _05363_);
  or (_18364_, _18363_, _18269_);
  or (_18365_, _18364_, _05357_);
  and (_18366_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and (_18367_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_18368_, _18367_, _18366_);
  and (_18369_, _18368_, _09527_);
  and (_18370_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_18371_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_18372_, _18371_, _18370_);
  and (_18373_, _18372_, _05352_);
  or (_18374_, _18373_, _18369_);
  or (_18375_, _18374_, _09540_);
  and (_18376_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and (_18377_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_18378_, _18377_, _18376_);
  and (_18379_, _18378_, _09527_);
  and (_18380_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_18381_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_18382_, _18381_, _18380_);
  and (_18383_, _18382_, _05352_);
  or (_18384_, _18383_, _18379_);
  or (_18385_, _18384_, _05373_);
  and (_18386_, _18385_, _09566_);
  and (_18387_, _18386_, _18375_);
  or (_18388_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_18389_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_18390_, _18389_, _05352_);
  and (_18391_, _18390_, _18388_);
  or (_18392_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_18393_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and (_18394_, _18393_, _09527_);
  and (_18395_, _18394_, _18392_);
  or (_18396_, _18395_, _18391_);
  or (_18397_, _18396_, _09540_);
  or (_18398_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_18399_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_18400_, _18399_, _05352_);
  and (_18401_, _18400_, _18398_);
  or (_18402_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_18403_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and (_18404_, _18403_, _09527_);
  and (_18405_, _18404_, _18402_);
  or (_18406_, _18405_, _18401_);
  or (_18407_, _18406_, _05373_);
  and (_18408_, _18407_, _05379_);
  and (_18409_, _18408_, _18397_);
  or (_18410_, _18409_, _18387_);
  and (_18411_, _18410_, _09581_);
  and (_18412_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_18413_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_18414_, _18413_, _18412_);
  and (_18415_, _18414_, _09527_);
  and (_18416_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_18417_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_18418_, _18417_, _18416_);
  and (_18419_, _18418_, _05352_);
  or (_18420_, _18419_, _18415_);
  or (_18421_, _18420_, _09540_);
  and (_18422_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_18423_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_18424_, _18423_, _18422_);
  and (_18425_, _18424_, _09527_);
  and (_18426_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_18427_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_18428_, _18427_, _18426_);
  and (_18429_, _18428_, _05352_);
  or (_18430_, _18429_, _18425_);
  or (_18431_, _18430_, _05373_);
  and (_18432_, _18431_, _09566_);
  and (_18433_, _18432_, _18421_);
  or (_18434_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_18435_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_18436_, _18435_, _18434_);
  and (_18437_, _18436_, _09527_);
  or (_18438_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_18439_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_18440_, _18439_, _18438_);
  and (_18441_, _18440_, _05352_);
  or (_18442_, _18441_, _18437_);
  or (_18443_, _18442_, _09540_);
  or (_18444_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_18445_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_18446_, _18445_, _18444_);
  and (_18447_, _18446_, _09527_);
  or (_18448_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_18449_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_18450_, _18449_, _18448_);
  and (_18451_, _18450_, _05352_);
  or (_18452_, _18451_, _18447_);
  or (_18453_, _18452_, _05373_);
  and (_18454_, _18453_, _05379_);
  and (_18455_, _18454_, _18443_);
  or (_18456_, _18455_, _18433_);
  and (_18457_, _18456_, _05361_);
  or (_18458_, _18457_, _18411_);
  and (_18459_, _18458_, _09682_);
  or (_18460_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_18461_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_18462_, _18461_, _18460_);
  and (_18463_, _18462_, _09527_);
  or (_18464_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_18465_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and (_18466_, _18465_, _18464_);
  and (_18467_, _18466_, _05352_);
  or (_18468_, _18467_, _18463_);
  and (_18469_, _18468_, _09540_);
  or (_18470_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_18471_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_18472_, _18471_, _18470_);
  and (_18473_, _18472_, _09527_);
  or (_18474_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_18476_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_18477_, _18476_, _18474_);
  and (_18478_, _18477_, _05352_);
  or (_18479_, _18478_, _18473_);
  and (_18480_, _18479_, _05373_);
  or (_18481_, _18480_, _18469_);
  and (_18482_, _18481_, _05379_);
  and (_18483_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_18484_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_18485_, _18484_, _18483_);
  and (_18486_, _18485_, _09527_);
  and (_18487_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_18488_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_18489_, _18488_, _18487_);
  and (_18490_, _18489_, _05352_);
  or (_18491_, _18490_, _18486_);
  and (_18492_, _18491_, _09540_);
  and (_18493_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and (_18494_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_18495_, _18494_, _18493_);
  and (_18496_, _18495_, _09527_);
  and (_18497_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and (_18498_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_18499_, _18498_, _18497_);
  and (_18500_, _18499_, _05352_);
  or (_18501_, _18500_, _18496_);
  and (_18502_, _18501_, _05373_);
  or (_18503_, _18502_, _18492_);
  and (_18504_, _18503_, _09566_);
  or (_18505_, _18504_, _18482_);
  and (_18506_, _18505_, _05361_);
  or (_18507_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_18508_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_18509_, _18508_, _05352_);
  and (_18510_, _18509_, _18507_);
  or (_18511_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_18512_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_18513_, _18512_, _09527_);
  and (_18514_, _18513_, _18511_);
  or (_18515_, _18514_, _18510_);
  and (_18516_, _18515_, _09540_);
  or (_18517_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_18518_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and (_18519_, _18518_, _05352_);
  and (_18520_, _18519_, _18517_);
  or (_18521_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_18522_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_18523_, _18522_, _09527_);
  and (_18524_, _18523_, _18521_);
  or (_18525_, _18524_, _18520_);
  and (_18526_, _18525_, _05373_);
  or (_18527_, _18526_, _18516_);
  and (_18528_, _18527_, _05379_);
  and (_18529_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and (_18530_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_18531_, _18530_, _18529_);
  and (_18532_, _18531_, _09527_);
  and (_18533_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_18534_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_18535_, _18534_, _18533_);
  and (_18536_, _18535_, _05352_);
  or (_18537_, _18536_, _18532_);
  and (_18538_, _18537_, _09540_);
  and (_18539_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_18540_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_18541_, _18540_, _18539_);
  and (_18542_, _18541_, _09527_);
  and (_18543_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_18544_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_18545_, _18544_, _18543_);
  and (_18546_, _18545_, _05352_);
  or (_18547_, _18546_, _18542_);
  and (_18548_, _18547_, _05373_);
  or (_18549_, _18548_, _18538_);
  and (_18550_, _18549_, _09566_);
  or (_18551_, _18550_, _18528_);
  and (_18552_, _18551_, _09581_);
  or (_18553_, _18552_, _18506_);
  and (_18554_, _18553_, _05363_);
  or (_18555_, _18554_, _18459_);
  or (_18557_, _18555_, _09739_);
  and (_18558_, _18557_, _18365_);
  or (_18559_, _18558_, _26838_);
  and (_18560_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_18561_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_18562_, _18561_, _18560_);
  and (_18563_, _18562_, _09527_);
  and (_18564_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_18565_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_18566_, _18565_, _18564_);
  and (_18567_, _18566_, _05352_);
  or (_18568_, _18567_, _18563_);
  or (_18569_, _18568_, _09540_);
  and (_18570_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_18571_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_18572_, _18571_, _18570_);
  and (_18573_, _18572_, _09527_);
  and (_18574_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_18575_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_18576_, _18575_, _18574_);
  and (_18577_, _18576_, _05352_);
  or (_18578_, _18577_, _18573_);
  or (_18579_, _18578_, _05373_);
  and (_18580_, _18579_, _09566_);
  and (_18581_, _18580_, _18569_);
  or (_18582_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_18583_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_18584_, _18583_, _18582_);
  and (_18585_, _18584_, _09527_);
  or (_18586_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_18588_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_18589_, _18588_, _18586_);
  and (_18590_, _18589_, _05352_);
  or (_18591_, _18590_, _18585_);
  or (_18592_, _18591_, _09540_);
  or (_18593_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_18594_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_18595_, _18594_, _18593_);
  and (_18596_, _18595_, _09527_);
  or (_18597_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_18598_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_18599_, _18598_, _18597_);
  and (_18600_, _18599_, _05352_);
  or (_18601_, _18600_, _18596_);
  or (_18602_, _18601_, _05373_);
  and (_18603_, _18602_, _05379_);
  and (_18604_, _18603_, _18592_);
  or (_18605_, _18604_, _18581_);
  and (_18606_, _18605_, _05361_);
  and (_18607_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_18608_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_18609_, _18608_, _18607_);
  and (_18610_, _18609_, _09527_);
  and (_18611_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_18612_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_18613_, _18612_, _18611_);
  and (_18614_, _18613_, _05352_);
  or (_18615_, _18614_, _18610_);
  or (_18616_, _18615_, _09540_);
  and (_18617_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_18618_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_18619_, _18618_, _18617_);
  and (_18620_, _18619_, _09527_);
  and (_18621_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_18622_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_18623_, _18622_, _18621_);
  and (_18624_, _18623_, _05352_);
  or (_18625_, _18624_, _18620_);
  or (_18626_, _18625_, _05373_);
  and (_18627_, _18626_, _09566_);
  and (_18628_, _18627_, _18616_);
  or (_18629_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_18630_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_18631_, _18630_, _05352_);
  and (_18632_, _18631_, _18629_);
  or (_18633_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_18634_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_18635_, _18634_, _09527_);
  and (_18636_, _18635_, _18633_);
  or (_18637_, _18636_, _18632_);
  or (_18638_, _18637_, _09540_);
  or (_18639_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_18640_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_18641_, _18640_, _05352_);
  and (_18642_, _18641_, _18639_);
  or (_18643_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_18644_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_18645_, _18644_, _09527_);
  and (_18646_, _18645_, _18643_);
  or (_18647_, _18646_, _18642_);
  or (_18648_, _18647_, _05373_);
  and (_18649_, _18648_, _05379_);
  and (_18650_, _18649_, _18638_);
  or (_18651_, _18650_, _18628_);
  and (_18652_, _18651_, _09581_);
  or (_18653_, _18652_, _18606_);
  and (_18654_, _18653_, _09682_);
  and (_18655_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and (_18656_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_18657_, _18656_, _18655_);
  and (_18658_, _18657_, _09527_);
  and (_18659_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and (_18660_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_18661_, _18660_, _18659_);
  and (_18662_, _18661_, _05352_);
  or (_18663_, _18662_, _18658_);
  and (_18664_, _18663_, _05373_);
  and (_18665_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and (_18666_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_18667_, _18666_, _18665_);
  and (_18668_, _18667_, _09527_);
  and (_18669_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and (_18670_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_18671_, _18670_, _18669_);
  and (_18672_, _18671_, _05352_);
  or (_18673_, _18672_, _18668_);
  and (_18674_, _18673_, _09540_);
  or (_18675_, _18674_, _18664_);
  and (_18676_, _18675_, _09566_);
  or (_18677_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_18679_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_18680_, _18679_, _05352_);
  and (_18681_, _18680_, _18677_);
  or (_18682_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_18683_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and (_18684_, _18683_, _09527_);
  and (_18685_, _18684_, _18682_);
  or (_18686_, _18685_, _18681_);
  and (_18687_, _18686_, _05373_);
  or (_18688_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_18689_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and (_18690_, _18689_, _05352_);
  and (_18691_, _18690_, _18688_);
  or (_18692_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_18693_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and (_18694_, _18693_, _09527_);
  and (_18695_, _18694_, _18692_);
  or (_18696_, _18695_, _18691_);
  and (_18697_, _18696_, _09540_);
  or (_18698_, _18697_, _18687_);
  and (_18699_, _18698_, _05379_);
  or (_18700_, _18699_, _18676_);
  and (_18701_, _18700_, _09581_);
  and (_18702_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_18703_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_18704_, _18703_, _18702_);
  and (_18705_, _18704_, _09527_);
  and (_18706_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_18707_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_18708_, _18707_, _18706_);
  and (_18709_, _18708_, _05352_);
  or (_18710_, _18709_, _18705_);
  and (_18711_, _18710_, _05373_);
  and (_18712_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_18713_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_18714_, _18713_, _18712_);
  and (_18715_, _18714_, _09527_);
  and (_18716_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_18717_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_18718_, _18717_, _18716_);
  and (_18719_, _18718_, _05352_);
  or (_18720_, _18719_, _18715_);
  and (_18721_, _18720_, _09540_);
  or (_18722_, _18721_, _18711_);
  and (_18723_, _18722_, _09566_);
  or (_18724_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_18725_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_18726_, _18725_, _18724_);
  and (_18727_, _18726_, _09527_);
  or (_18728_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_18729_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_18730_, _18729_, _18728_);
  and (_18731_, _18730_, _05352_);
  or (_18732_, _18731_, _18727_);
  and (_18733_, _18732_, _05373_);
  or (_18734_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_18735_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_18736_, _18735_, _18734_);
  and (_18737_, _18736_, _09527_);
  or (_18738_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_18739_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_18740_, _18739_, _18738_);
  and (_18741_, _18740_, _05352_);
  or (_18742_, _18741_, _18737_);
  and (_18743_, _18742_, _09540_);
  or (_18744_, _18743_, _18733_);
  and (_18745_, _18744_, _05379_);
  or (_18746_, _18745_, _18723_);
  and (_18747_, _18746_, _05361_);
  or (_18748_, _18747_, _18701_);
  and (_18749_, _18748_, _05363_);
  or (_18750_, _18749_, _18654_);
  or (_18751_, _18750_, _05357_);
  and (_18752_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_18753_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_18754_, _18753_, _18752_);
  and (_18755_, _18754_, _09527_);
  and (_18756_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_18757_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_18758_, _18757_, _18756_);
  and (_18759_, _18758_, _05352_);
  or (_18760_, _18759_, _18755_);
  or (_18761_, _18760_, _09540_);
  and (_18762_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_18763_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_18764_, _18763_, _18762_);
  and (_18765_, _18764_, _09527_);
  and (_18766_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_18767_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_18768_, _18767_, _18766_);
  and (_18769_, _18768_, _05352_);
  or (_18770_, _18769_, _18765_);
  or (_18771_, _18770_, _05373_);
  and (_18772_, _18771_, _09566_);
  and (_18773_, _18772_, _18761_);
  or (_18774_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_18775_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_18776_, _18775_, _05352_);
  and (_18777_, _18776_, _18774_);
  or (_18778_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_18779_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_18780_, _18779_, _09527_);
  and (_18781_, _18780_, _18778_);
  or (_18782_, _18781_, _18777_);
  or (_18783_, _18782_, _09540_);
  or (_18784_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_18785_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_18786_, _18785_, _05352_);
  and (_18787_, _18786_, _18784_);
  or (_18788_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_18790_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_18791_, _18790_, _09527_);
  and (_18792_, _18791_, _18788_);
  or (_18793_, _18792_, _18787_);
  or (_18794_, _18793_, _05373_);
  and (_18795_, _18794_, _05379_);
  and (_18796_, _18795_, _18783_);
  or (_18797_, _18796_, _18773_);
  and (_18798_, _18797_, _09581_);
  and (_18799_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_18800_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_18801_, _18800_, _18799_);
  and (_18802_, _18801_, _09527_);
  and (_18803_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_18804_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_18805_, _18804_, _18803_);
  and (_18806_, _18805_, _05352_);
  or (_18807_, _18806_, _18802_);
  or (_18808_, _18807_, _09540_);
  and (_18809_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_18810_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_18811_, _18810_, _18809_);
  and (_18812_, _18811_, _09527_);
  and (_18813_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_18814_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_18815_, _18814_, _18813_);
  and (_18816_, _18815_, _05352_);
  or (_18817_, _18816_, _18812_);
  or (_18818_, _18817_, _05373_);
  and (_18819_, _18818_, _09566_);
  and (_18820_, _18819_, _18808_);
  or (_18821_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_18822_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_18823_, _18822_, _18821_);
  and (_18824_, _18823_, _09527_);
  or (_18825_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_18826_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_18827_, _18826_, _18825_);
  and (_18828_, _18827_, _05352_);
  or (_18829_, _18828_, _18824_);
  or (_18830_, _18829_, _09540_);
  or (_18831_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_18832_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_18833_, _18832_, _18831_);
  and (_18834_, _18833_, _09527_);
  or (_18835_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_18836_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_18837_, _18836_, _18835_);
  and (_18838_, _18837_, _05352_);
  or (_18839_, _18838_, _18834_);
  or (_18840_, _18839_, _05373_);
  and (_18841_, _18840_, _05379_);
  and (_18842_, _18841_, _18830_);
  or (_18843_, _18842_, _18820_);
  and (_18844_, _18843_, _05361_);
  or (_18845_, _18844_, _18798_);
  and (_18846_, _18845_, _09682_);
  or (_18847_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_18848_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_18849_, _18848_, _18847_);
  and (_18850_, _18849_, _09527_);
  or (_18851_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_18852_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_18853_, _18852_, _18851_);
  and (_18854_, _18853_, _05352_);
  or (_18855_, _18854_, _18850_);
  and (_18856_, _18855_, _09540_);
  or (_18857_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_18858_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_18859_, _18858_, _18857_);
  and (_18860_, _18859_, _09527_);
  or (_18861_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_18862_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_18863_, _18862_, _18861_);
  and (_18864_, _18863_, _05352_);
  or (_18865_, _18864_, _18860_);
  and (_18866_, _18865_, _05373_);
  or (_18867_, _18866_, _18856_);
  and (_18868_, _18867_, _05379_);
  and (_18869_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_18870_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_18871_, _18870_, _18869_);
  and (_18872_, _18871_, _09527_);
  and (_18873_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_18874_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_18875_, _18874_, _18873_);
  and (_18876_, _18875_, _05352_);
  or (_18877_, _18876_, _18872_);
  and (_18878_, _18877_, _09540_);
  and (_18879_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_18880_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_18881_, _18880_, _18879_);
  and (_18882_, _18881_, _09527_);
  and (_18883_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_18884_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_18885_, _18884_, _18883_);
  and (_18886_, _18885_, _05352_);
  or (_18887_, _18886_, _18882_);
  and (_18888_, _18887_, _05373_);
  or (_18889_, _18888_, _18878_);
  and (_18890_, _18889_, _09566_);
  or (_18891_, _18890_, _18868_);
  and (_18892_, _18891_, _05361_);
  or (_18893_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_18894_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and (_18895_, _18894_, _05352_);
  and (_18896_, _18895_, _18893_);
  or (_18897_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_18898_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_18899_, _18898_, _09527_);
  and (_18900_, _18899_, _18897_);
  or (_18901_, _18900_, _18896_);
  and (_18902_, _18901_, _09540_);
  or (_18903_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_18904_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_18905_, _18904_, _05352_);
  and (_18906_, _18905_, _18903_);
  or (_18907_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_18908_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and (_18909_, _18908_, _09527_);
  and (_18910_, _18909_, _18907_);
  or (_18911_, _18910_, _18906_);
  and (_18912_, _18911_, _05373_);
  or (_18913_, _18912_, _18902_);
  and (_18914_, _18913_, _05379_);
  and (_18915_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_18916_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_18917_, _18916_, _18915_);
  and (_18918_, _18917_, _09527_);
  and (_18919_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_18920_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_18921_, _18920_, _18919_);
  and (_18922_, _18921_, _05352_);
  or (_18923_, _18922_, _18918_);
  and (_18924_, _18923_, _09540_);
  and (_18925_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_18926_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_18927_, _18926_, _18925_);
  and (_18928_, _18927_, _09527_);
  and (_18929_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_18930_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_18931_, _18930_, _18929_);
  and (_18932_, _18931_, _05352_);
  or (_18933_, _18932_, _18928_);
  and (_18934_, _18933_, _05373_);
  or (_18935_, _18934_, _18924_);
  and (_18936_, _18935_, _09566_);
  or (_18937_, _18936_, _18914_);
  and (_18938_, _18937_, _09581_);
  or (_18939_, _18938_, _18892_);
  and (_18940_, _18939_, _05363_);
  or (_18941_, _18940_, _18846_);
  or (_18942_, _18941_, _09739_);
  and (_18943_, _18942_, _18751_);
  or (_18944_, _18943_, _04360_);
  and (_18945_, _18944_, _18559_);
  or (_18946_, _18945_, _05401_);
  or (_18947_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_18948_, _18947_, _22761_);
  and (_10902_, _18948_, _18946_);
  and (_18949_, _15481_, _23676_);
  and (_18950_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_10905_, _18950_, _18949_);
  and (_18951_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_18952_, _09519_, _23718_);
  or (_27102_, _18952_, _18951_);
  and (_18953_, _24209_, _23676_);
  and (_18954_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_27281_, _18954_, _18953_);
  and (_18955_, _17312_, _23718_);
  and (_18956_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_26938_, _18956_, _18955_);
  and (_18957_, _17038_, _23589_);
  and (_18958_, _17040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or (_27309_, _18958_, _18957_);
  and (_18959_, _16443_, _23676_);
  and (_18960_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or (_26960_, _18960_, _18959_);
  and (_18961_, _15895_, _23635_);
  and (_18962_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_26981_, _18962_, _18961_);
  and (_18963_, _25118_, _24671_);
  nand (_18964_, _18963_, _23522_);
  or (_18965_, _18963_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_18966_, _18965_, _24629_);
  and (_18967_, _18966_, _18964_);
  nand (_18968_, _25124_, _23585_);
  or (_18969_, _25124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_18970_, _18969_, _23880_);
  and (_18971_, _18970_, _18968_);
  and (_18972_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_18973_, _18972_, rst);
  or (_18974_, _18973_, _18971_);
  or (_10929_, _18974_, _18967_);
  and (_18975_, _25400_, _23791_);
  and (_18976_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_27241_, _18976_, _18975_);
  and (_18977_, _16443_, _23791_);
  and (_18978_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or (_26961_, _18978_, _18977_);
  and (_18979_, _16443_, _23838_);
  and (_18980_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or (_26962_, _18980_, _18979_);
  and (_18981_, _25309_, _24671_);
  nand (_18982_, _18981_, _23522_);
  or (_18983_, _18981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_18984_, _18983_, _24629_);
  and (_18985_, _18984_, _18982_);
  nand (_18986_, _25317_, _23585_);
  or (_18987_, _25317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_18988_, _18987_, _23880_);
  and (_18989_, _18988_, _18986_);
  and (_18990_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_18991_, _18990_, rst);
  or (_18992_, _18991_, _18989_);
  or (_10945_, _18992_, _18985_);
  and (_18993_, _15895_, _23589_);
  and (_18994_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_26983_, _18994_, _18993_);
  and (_18995_, _16443_, _23635_);
  and (_18996_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or (_26963_, _18996_, _18995_);
  and (_18997_, _16443_, _23755_);
  and (_18998_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or (_26964_, _18998_, _18997_);
  nand (_18999_, _25615_, _24491_);
  or (_26871_[2], _18999_, _24531_);
  and (_19000_, _15895_, _23755_);
  and (_19001_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_26982_, _19001_, _19000_);
  and (_19002_, _24577_, _23791_);
  and (_19003_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or (_27230_, _19003_, _19002_);
  and (_19004_, _15995_, _23755_);
  and (_19005_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or (_26994_, _19005_, _19004_);
  and (_19006_, _25407_, _24671_);
  nand (_19007_, _19006_, _23522_);
  or (_19008_, _19006_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_19009_, _19008_, _24629_);
  and (_19010_, _19009_, _19007_);
  nand (_19011_, _25413_, _23585_);
  or (_19012_, _25413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_19013_, _19012_, _23880_);
  and (_19014_, _19013_, _19011_);
  and (_19015_, _25129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_19016_, _19015_, rst);
  or (_19017_, _19016_, _19014_);
  or (_10963_, _19017_, _19010_);
  and (_19018_, _16443_, _23589_);
  and (_19019_, _16445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or (_26965_, _19019_, _19018_);
  and (_19020_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and (_19021_, _13826_, _23635_);
  or (_27115_, _19021_, _19020_);
  nand (_19022_, _23927_, _23628_);
  and (_19023_, _24152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_19024_, _24165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_19025_, _24155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand (_19026_, _19025_, _24154_);
  nor (_19027_, _19026_, _24156_);
  nor (_19028_, _19027_, _19024_);
  nor (_19029_, _19028_, _23921_);
  or (_19030_, _19029_, _19023_);
  or (_19031_, _19030_, _23927_);
  and (_19032_, _19031_, _22761_);
  and (_10977_, _19032_, _19022_);
  and (_19033_, _13485_, _23676_);
  and (_19034_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_26967_, _19034_, _19033_);
  and (_19035_, _04532_, _23982_);
  and (_19036_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_27178_, _19036_, _19035_);
  and (_19037_, _13485_, _23718_);
  and (_19038_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_26968_, _19038_, _19037_);
  and (_19039_, _13485_, _23982_);
  and (_19040_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_26970_, _19040_, _19039_);
  and (_19041_, _13827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  and (_19042_, _13826_, _23755_);
  or (_27116_, _19042_, _19041_);
  and (_19043_, _04532_, _23838_);
  and (_19044_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_27177_, _19044_, _19043_);
  and (_19045_, _17990_, _23718_);
  and (_19046_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or (_27257_, _19046_, _19045_);
  and (_19047_, _25400_, _23676_);
  and (_19048_, _25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_27240_, _19048_, _19047_);
  and (_19049_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_19050_, _09519_, _23791_);
  or (_27101_, _19050_, _19049_);
  and (_19051_, _02785_, _23635_);
  and (_19052_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  or (_27185_, _19052_, _19051_);
  and (_19053_, _13485_, _23635_);
  and (_19054_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_26971_, _19054_, _19053_);
  and (_19055_, _17990_, _23791_);
  and (_19056_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or (_27256_, _19056_, _19055_);
  and (_19057_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_19058_, _17978_, _23589_);
  or (_27239_, _19058_, _19057_);
  and (_19059_, _17990_, _23676_);
  and (_19060_, _17992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or (_27255_, _19060_, _19059_);
  and (_19061_, _24567_, _23982_);
  and (_19062_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or (_27086_, _19062_, _19061_);
  not (_19063_, _24259_);
  nand (_19064_, _24307_, _19063_);
  nor (_19065_, _19064_, _24432_);
  and (_19066_, _22764_, _24270_);
  and (_19067_, _19066_, _25615_);
  and (_19068_, _19067_, _24359_);
  and (_19069_, _24381_, _24335_);
  and (_19070_, _19069_, _19068_);
  and (_19071_, _24405_, _24282_);
  and (_19072_, _19071_, _19070_);
  and (_26907_, _19072_, _19065_);
  and (_19073_, _17972_, _23635_);
  and (_19074_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_11035_, _19074_, _19073_);
  and (_19075_, _24577_, _23718_);
  and (_19076_, _24579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or (_27231_, _19076_, _19075_);
  and (_19077_, _13485_, _23755_);
  and (_19078_, _13487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_11041_, _19078_, _19077_);
  and (_19079_, _17972_, _23589_);
  and (_19080_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_11043_, _19080_, _19079_);
  and (_19081_, _23843_, _23718_);
  and (_19082_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or (_26942_, _19082_, _19081_);
  and (_19083_, _23838_, _23652_);
  and (_19084_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or (_11048_, _19084_, _19083_);
  and (_19085_, _15481_, _23755_);
  and (_19086_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or (_11051_, _19086_, _19085_);
  and (_19087_, _23982_, _23855_);
  and (_19088_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or (_11057_, _19088_, _19087_);
  and (_19089_, _23855_, _23718_);
  and (_19090_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or (_11061_, _19090_, _19089_);
  and (_19091_, _23850_, _23589_);
  and (_19092_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_11063_, _19092_, _19091_);
  and (_19093_, _15481_, _23589_);
  and (_19094_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or (_11065_, _19094_, _19093_);
  and (_19095_, _24547_, _23676_);
  and (_19096_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_11068_, _19096_, _19095_);
  and (_19097_, _24080_, _23791_);
  and (_19098_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_27295_, _19098_, _19097_);
  and (_19099_, _23855_, _23838_);
  and (_19100_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or (_26939_, _19100_, _19099_);
  and (_19101_, _23755_, _23652_);
  and (_19102_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or (_27294_, _19102_, _19101_);
  and (_19103_, _17972_, _23755_);
  and (_19104_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_27254_, _19104_, _19103_);
  and (_19105_, _17001_, _23635_);
  and (_19106_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_11079_, _19106_, _19105_);
  and (_19107_, _23807_, _23676_);
  and (_19108_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_11083_, _19108_, _19107_);
  and (_19109_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and (_19110_, _02858_, _23635_);
  or (_11085_, _19110_, _19109_);
  and (_19111_, _23811_, _23718_);
  and (_19112_, _23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or (_11090_, _19112_, _19111_);
  and (_19113_, _24547_, _23838_);
  and (_19114_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_11097_, _19114_, _19113_);
  and (_19115_, _04532_, _23635_);
  and (_19116_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_11100_, _19116_, _19115_);
  and (_19117_, _24547_, _23635_);
  and (_19118_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_11102_, _19118_, _19117_);
  and (_19119_, _23843_, _23676_);
  and (_19120_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or (_11104_, _19120_, _19119_);
  and (_19121_, _23855_, _23635_);
  and (_19122_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or (_26940_, _19122_, _19121_);
  and (_19123_, _24080_, _23982_);
  and (_19124_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_11108_, _19124_, _19123_);
  and (_19125_, _23855_, _23755_);
  and (_19126_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or (_26941_, _19126_, _19125_);
  and (_19127_, _16703_, _23755_);
  and (_19128_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or (_11112_, _19128_, _19127_);
  and (_19129_, _23963_, _23838_);
  and (_19130_, _23966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_11114_, _19130_, _19129_);
  and (_19131_, _24547_, _23718_);
  and (_19132_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_11116_, _19132_, _19131_);
  and (_19133_, _24547_, _23982_);
  and (_19134_, _24550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_11119_, _19134_, _19133_);
  and (_19135_, _23855_, _23589_);
  and (_19136_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or (_11123_, _19136_, _19135_);
  and (_19137_, _16703_, _23589_);
  and (_19138_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_11125_, _19138_, _19137_);
  and (_19139_, _03296_, _23676_);
  and (_19140_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_11129_, _19140_, _19139_);
  and (_19141_, _12516_, _23755_);
  and (_19142_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or (_11132_, _19142_, _19141_);
  and (_19143_, _23982_, _23807_);
  and (_19144_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_11137_, _19144_, _19143_);
  and (_19145_, _23807_, _23755_);
  and (_19146_, _23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_11139_, _19146_, _19145_);
  and (_19147_, _24123_, _23755_);
  and (_19148_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_11141_, _19148_, _19147_);
  and (_19149_, _23982_, _23029_);
  and (_19150_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_11144_, _19150_, _19149_);
  and (_19151_, _15895_, _23791_);
  and (_19152_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_11147_, _19152_, _19151_);
  and (_19153_, _23850_, _23718_);
  and (_19154_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or (_11149_, _19154_, _19153_);
  and (_19155_, _23982_, _23850_);
  and (_19156_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or (_11151_, _19156_, _19155_);
  and (_19157_, _17312_, _23589_);
  and (_19158_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_11154_, _19158_, _19157_);
  and (_19159_, _23855_, _23676_);
  and (_19160_, _23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or (_11159_, _19160_, _19159_);
  and (_19161_, _23850_, _23635_);
  and (_19162_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or (_11161_, _19162_, _19161_);
  and (_19163_, _12516_, _23838_);
  and (_19164_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or (_26974_, _19164_, _19163_);
  and (_19165_, _23791_, _23029_);
  and (_19166_, _23591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_11168_, _19166_, _19165_);
  and (_19167_, _17312_, _23635_);
  and (_19168_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_11170_, _19168_, _19167_);
  and (_19169_, _24209_, _23589_);
  and (_19170_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_27285_, _19170_, _19169_);
  and (_19171_, _23850_, _23791_);
  and (_19172_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or (_11180_, _19172_, _19171_);
  and (_19173_, _24209_, _23982_);
  and (_19174_, _24211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_11182_, _19174_, _19173_);
  and (_19175_, _23850_, _23838_);
  and (_19176_, _23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or (_11187_, _19176_, _19175_);
  and (_19177_, _17312_, _23755_);
  and (_19178_, _17314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_11192_, _19178_, _19177_);
  and (_19179_, _24123_, _23718_);
  and (_19180_, _24125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_11196_, _19180_, _19179_);
  and (_19181_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_19182_, _02858_, _23982_);
  or (_11201_, _19182_, _19181_);
  and (_19183_, _04532_, _23791_);
  and (_19184_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_11206_, _19184_, _19183_);
  and (_19185_, _23982_, _23652_);
  and (_19186_, _23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or (_11213_, _19186_, _19185_);
  and (_19187_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_19188_, _02858_, _23838_);
  or (_11217_, _19188_, _19187_);
  and (_19189_, _04532_, _23676_);
  and (_19190_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_27175_, _19190_, _19189_);
  and (_19191_, _15895_, _23838_);
  and (_19192_, _15897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_11222_, _19192_, _19191_);
  and (_19193_, _24567_, _23676_);
  and (_19194_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or (_11226_, _19194_, _19193_);
  and (_19195_, _15995_, _23791_);
  and (_19196_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or (_11235_, _19196_, _19195_);
  and (_19197_, _24119_, _23838_);
  and (_19198_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_11237_, _19198_, _19197_);
  and (_19199_, _24119_, _23791_);
  and (_19200_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_11240_, _19200_, _19199_);
  and (_19201_, _25088_, _23982_);
  and (_19202_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or (_11242_, _19202_, _19201_);
  and (_19203_, _25088_, _23718_);
  and (_19204_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or (_27224_, _19204_, _19203_);
  and (_19205_, _15481_, _23718_);
  and (_19206_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or (_11245_, _19206_, _19205_);
  and (_19207_, _25046_, _23755_);
  and (_19208_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or (_11247_, _19208_, _19207_);
  and (_19209_, _25046_, _23791_);
  and (_19210_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or (_27222_, _19210_, _19209_);
  and (_19211_, _24991_, _23589_);
  and (_19212_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_11255_, _19212_, _19211_);
  and (_19213_, _15481_, _23791_);
  and (_19214_, _15483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_11257_, _19214_, _19213_);
  and (_19215_, _24991_, _23718_);
  and (_19216_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_11263_, _19216_, _19215_);
  and (_19217_, _24925_, _23589_);
  and (_19218_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_11265_, _19218_, _19217_);
  and (_19219_, _24925_, _23718_);
  and (_19220_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_11280_, _19220_, _19219_);
  and (_19221_, _24909_, _23838_);
  and (_19222_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or (_11283_, _19222_, _19221_);
  and (_19223_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and (_19224_, _02840_, _23676_);
  or (_11285_, _19224_, _19223_);
  and (_19225_, _24909_, _23676_);
  and (_19226_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or (_11287_, _19226_, _19225_);
  and (_19227_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_19228_, _09519_, _23982_);
  or (_11289_, _19228_, _19227_);
  and (_19229_, _24833_, _23589_);
  and (_19230_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or (_11291_, _19230_, _19229_);
  and (_19231_, _24833_, _23635_);
  and (_19232_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or (_27217_, _19232_, _19231_);
  and (_19233_, _24833_, _23791_);
  and (_19234_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or (_11294_, _19234_, _19233_);
  and (_19235_, _24610_, _23755_);
  and (_19236_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_11297_, _19236_, _19235_);
  and (_19237_, _16850_, _23676_);
  and (_19238_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or (_11300_, _19238_, _19237_);
  and (_19239_, _16850_, _23718_);
  and (_19240_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or (_11305_, _19240_, _19239_);
  and (_19241_, _24605_, _23838_);
  and (_19242_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_11307_, _19242_, _19241_);
  and (_19243_, _24722_, _23755_);
  and (_19244_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or (_11310_, _19244_, _19243_);
  and (_19245_, _24722_, _23982_);
  and (_19246_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or (_11312_, _19246_, _19245_);
  and (_19247_, _24722_, _23676_);
  and (_19248_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or (_27208_, _19248_, _19247_);
  and (_19249_, _24680_, _23589_);
  and (_19250_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or (_11317_, _19250_, _19249_);
  and (_19251_, _24680_, _23982_);
  and (_19252_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or (_27205_, _19252_, _19251_);
  and (_19253_, _24680_, _23676_);
  and (_19254_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or (_11320_, _19254_, _19253_);
  and (_19255_, _24622_, _23635_);
  and (_19256_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_11325_, _19256_, _19255_);
  and (_19257_, _04532_, _23718_);
  and (_19258_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_27176_, _19258_, _19257_);
  and (_19259_, _24610_, _23718_);
  and (_19260_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_11329_, _19260_, _19259_);
  and (_19261_, _16703_, _23791_);
  and (_19262_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_11344_, _19262_, _19261_);
  and (_19263_, _25088_, _23755_);
  and (_19264_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or (_11346_, _19264_, _19263_);
  and (_19265_, _25046_, _23838_);
  and (_19266_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or (_11352_, _19266_, _19265_);
  and (_19267_, _16081_, _23635_);
  and (_19268_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or (_11356_, _19268_, _19267_);
  and (_19269_, _24991_, _23982_);
  and (_19270_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_11364_, _19270_, _19269_);
  and (_19271_, _24925_, _23982_);
  and (_19272_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_11366_, _19272_, _19271_);
  and (_19273_, _16081_, _23982_);
  and (_19274_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or (_26978_, _19274_, _19273_);
  and (_19275_, _24925_, _23676_);
  and (_19276_, _24927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_27220_, _19276_, _19275_);
  and (_19277_, _24909_, _23635_);
  and (_19278_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or (_11370_, _19278_, _19277_);
  and (_19279_, _16703_, _23676_);
  and (_19280_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or (_11372_, _19280_, _19279_);
  and (_19281_, _16850_, _23791_);
  and (_19282_, _16852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or (_11380_, _19282_, _19281_);
  and (_19283_, _24680_, _23718_);
  and (_19284_, _24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or (_11386_, _19284_, _19283_);
  and (_19285_, _24622_, _23589_);
  and (_19286_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_11388_, _19286_, _19285_);
  and (_19287_, _24119_, _23635_);
  and (_19288_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_11392_, _19288_, _19287_);
  and (_19289_, _25046_, _23589_);
  and (_19290_, _25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or (_11394_, _19290_, _19289_);
  and (_19291_, _24909_, _23791_);
  and (_19292_, _24911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or (_11397_, _19292_, _19291_);
  and (_19293_, _24833_, _23718_);
  and (_19294_, _24835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or (_27215_, _19294_, _19293_);
  and (_19295_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_19296_, _17978_, _23676_);
  or (_27237_, _19296_, _19295_);
  and (_19297_, _24605_, _23676_);
  and (_19298_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_27209_, _19298_, _19297_);
  and (_19299_, _24722_, _23791_);
  and (_19300_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or (_11403_, _19300_, _19299_);
  and (_19301_, _24610_, _23838_);
  and (_19302_, _24612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_11405_, _19302_, _19301_);
  and (_19303_, _24991_, _23676_);
  and (_19304_, _24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_11408_, _19304_, _19303_);
  and (_19305_, _16703_, _23982_);
  and (_19306_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_11410_, _19306_, _19305_);
  and (_19307_, _24605_, _23755_);
  and (_19308_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_11412_, _19308_, _19307_);
  and (_19309_, _24593_, _23755_);
  and (_19310_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or (_11422_, _19310_, _19309_);
  and (_19311_, _16703_, _23838_);
  and (_19312_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or (_11424_, _19312_, _19311_);
  and (_19313_, _16703_, _23718_);
  and (_19314_, _16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_11428_, _19314_, _19313_);
  and (_19315_, _01802_, _23791_);
  and (_19316_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_27037_, _19316_, _19315_);
  and (_19317_, _02200_, _23982_);
  and (_19318_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_11431_, _19318_, _19317_);
  and (_19319_, _02221_, _23755_);
  and (_19320_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_26992_, _19320_, _19319_);
  and (_19321_, _02221_, _23676_);
  and (_19322_, _02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_11435_, _19322_, _19321_);
  and (_19323_, _24934_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_19324_, _24850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_19325_, _24850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_19326_, _19325_, _19324_);
  nor (_19327_, _19326_, _24933_);
  or (_19328_, _19327_, _24847_);
  or (_19329_, _19328_, _19323_);
  or (_19330_, _19326_, _24938_);
  and (_19331_, _19330_, _22761_);
  and (_11447_, _19331_, _19329_);
  and (_19332_, _03189_, _23718_);
  and (_19333_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_11450_, _19333_, _19332_);
  or (_19334_, _25001_, _24945_);
  and (_19335_, _19334_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_19336_, _19335_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_19337_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_19338_, _24850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_19339_, _19338_, _19337_);
  or (_19340_, _19339_, _24849_);
  nor (_19341_, _02148_, _02117_);
  nor (_19342_, _19341_, _24849_);
  not (_19343_, _19342_);
  and (_19344_, _19343_, _19340_);
  nand (_19345_, _19344_, _19336_);
  nand (_19346_, _19345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_19347_, _19346_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_19348_, _23875_, _23887_);
  nor (_19349_, _24630_, _19348_);
  or (_19350_, _19349_, _19347_);
  nand (_19351_, _19349_, _23812_);
  and (_19352_, _19351_, _19350_);
  nand (_19353_, _19352_, _24802_);
  nand (_19354_, _24801_, _23784_);
  and (_19355_, _19354_, _22761_);
  and (_11460_, _19355_, _19353_);
  and (_11482_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _22761_);
  and (_19356_, _16081_, _23589_);
  and (_19357_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or (_11485_, _19357_, _19356_);
  and (_19358_, _03648_, _23635_);
  and (_19359_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_11490_, _19359_, _19358_);
  or (_19360_, _03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_11492_, _19360_, _03392_);
  and (_19361_, _16707_, _23982_);
  and (_19362_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_27279_, _19362_, _19361_);
  and (_19363_, _16081_, _23755_);
  and (_19364_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or (_26979_, _19364_, _19363_);
  and (_19365_, _05445_, _23635_);
  and (_19366_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or (_11501_, _19366_, _19365_);
  and (_19367_, _05445_, _23982_);
  and (_19368_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  or (_27173_, _19368_, _19367_);
  not (_19369_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_19370_, _19335_, _19369_);
  not (_19371_, _19341_);
  or (_19372_, _19371_, _19340_);
  or (_19373_, _19372_, _19370_);
  and (_19374_, _19373_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_19375_, _19374_, _04626_);
  and (_19376_, _24631_, _23875_);
  and (_19377_, _19376_, _24671_);
  or (_19378_, _19377_, _19375_);
  nand (_19379_, _19377_, _23522_);
  and (_19380_, _19379_, _19378_);
  or (_19381_, _19380_, _24801_);
  nand (_19382_, _24801_, _23585_);
  and (_19383_, _19382_, _22761_);
  and (_11510_, _19383_, _19381_);
  and (_11516_, _26272_, _22761_);
  and (_19384_, _24798_, _24688_);
  or (_19385_, _19384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_19386_, _19385_, _24802_);
  nand (_19387_, _19384_, _23522_);
  and (_19388_, _19387_, _19386_);
  nor (_19389_, _24802_, _23748_);
  or (_19390_, _19389_, _19388_);
  and (_11523_, _19390_, _22761_);
  and (_19391_, _24877_, _24865_);
  nand (_19392_, _24881_, _19391_);
  or (_19393_, _24892_, _24881_);
  and (_19394_, _19393_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_19395_, _19394_, _19392_);
  or (_19396_, _19395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nand (_19397_, _24902_, _24933_);
  or (_19398_, _24874_, _24855_);
  and (_19399_, _19398_, _19397_);
  or (_19400_, _19399_, _24921_);
  and (_19401_, _24921_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_19402_, _19401_, _24938_);
  and (_19403_, _19402_, _22761_);
  and (_19404_, _19403_, _19400_);
  and (_11529_, _19404_, _19396_);
  and (_11532_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _22761_);
  or (_19405_, _19393_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_19406_, _19405_, _19399_);
  or (_19407_, _19337_, _24847_);
  or (_19408_, _19407_, _19406_);
  and (_19409_, _19392_, _24848_);
  or (_19410_, _19409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_19411_, _19410_, _22761_);
  and (_11534_, _19411_, _19408_);
  and (_11536_, _00364_, _22761_);
  not (_19412_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_19413_, _19412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_19414_, _19342_, _19339_);
  not (_19415_, _19414_);
  or (_19416_, _19415_, _19370_);
  and (_19417_, _19416_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_19418_, _19417_, _19413_);
  and (_19419_, _19376_, _23919_);
  or (_19420_, _19419_, _19418_);
  nand (_19421_, _19419_, _23522_);
  and (_19422_, _19421_, _19420_);
  or (_19423_, _19422_, _24801_);
  nand (_19424_, _24801_, _23628_);
  and (_19425_, _19424_, _22761_);
  and (_11550_, _19425_, _19423_);
  and (_19426_, _16707_, _23838_);
  and (_19427_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_11554_, _19427_, _19426_);
  and (_19428_, _19376_, _23925_);
  and (_19429_, _19428_, _23812_);
  nand (_19430_, _25953_, _23888_);
  nand (_19431_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_19432_, _19414_, _19336_);
  or (_19433_, _19432_, _19431_);
  or (_19434_, _19433_, _19428_);
  nand (_19435_, _19434_, _19430_);
  or (_19436_, _19435_, _19429_);
  nand (_19437_, _24801_, _23832_);
  and (_19438_, _19437_, _22761_);
  and (_11558_, _19438_, _19436_);
  and (_19439_, _24671_, _24634_);
  nand (_19440_, _19439_, _23522_);
  or (_19441_, _19439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_19442_, _19441_, _24653_);
  and (_19443_, _19442_, _19440_);
  nor (_19444_, _24653_, _23585_);
  or (_19445_, _19444_, _19443_);
  and (_11561_, _19445_, _22761_);
  and (_19446_, _16081_, _23676_);
  and (_19447_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or (_11563_, _19447_, _19446_);
  and (_19448_, _25529_, _23982_);
  and (_19449_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_11567_, _19449_, _19448_);
  and (_19450_, _02092_, _23838_);
  and (_19451_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_11569_, _19451_, _19450_);
  and (_19452_, _16081_, _23791_);
  and (_19453_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or (_11574_, _19453_, _19452_);
  and (_19454_, _09520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and (_19455_, _09519_, _23635_);
  or (_11577_, _19455_, _19454_);
  nand (_19456_, _24934_, _24849_);
  nand (_19457_, _19324_, _24847_);
  and (_19458_, _19457_, _22761_);
  and (_11586_, _19458_, _19456_);
  and (_19459_, _02750_, _23838_);
  and (_19460_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_11588_, _19460_, _19459_);
  and (_19461_, _03010_, _23635_);
  and (_19462_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_11591_, _19462_, _19461_);
  and (_19463_, _16707_, _23718_);
  and (_19464_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_27278_, _19464_, _19463_);
  and (_19465_, _24708_, _24671_);
  or (_19466_, _19465_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_19467_, _19466_, _24716_);
  nand (_19468_, _19465_, _23522_);
  and (_19469_, _19468_, _19467_);
  nor (_19470_, _24716_, _23585_);
  or (_19471_, _19470_, _19469_);
  and (_11597_, _19471_, _22761_);
  not (_19472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_19473_, _23938_, _19472_);
  or (_19474_, _19473_, _02413_);
  and (_19475_, _19474_, _24147_);
  or (_19476_, _19473_, _02422_);
  and (_19477_, _19476_, _24191_);
  nand (_19478_, _23938_, _23946_);
  and (_19479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_19480_, _19479_, _19478_);
  or (_19481_, _19480_, _15456_);
  or (_19482_, _19481_, _19477_);
  or (_19483_, _19482_, _19475_);
  nor (_19484_, _23927_, rst);
  and (_19485_, _19484_, _23922_);
  and (_11603_, _19485_, _19483_);
  and (_19486_, _03273_, _23755_);
  and (_19487_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_11605_, _19487_, _19486_);
  and (_19488_, _03648_, _23676_);
  and (_19489_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_11610_, _19489_, _19488_);
  and (_19490_, _03189_, _23838_);
  and (_19491_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_11639_, _19491_, _19490_);
  and (_19492_, _03302_, _23676_);
  and (_19493_, _03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  or (_11642_, _19493_, _19492_);
  nor (_11644_, _00759_, rst);
  and (_11646_, _00366_, _22761_);
  and (_11650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _22761_);
  and (_19494_, _05445_, _23755_);
  and (_19495_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  or (_27174_, _19495_, _19494_);
  and (_19496_, _17001_, _23982_);
  and (_19497_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or (_11680_, _19497_, _19496_);
  and (_19498_, _02092_, _23982_);
  and (_19499_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_11685_, _19499_, _19498_);
  and (_19500_, _03010_, _23755_);
  and (_19501_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_11688_, _19501_, _19500_);
  and (_19502_, _06255_, _23676_);
  and (_19503_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or (_11691_, _19503_, _19502_);
  and (_19504_, _24573_, _23755_);
  and (_19505_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or (_11698_, _19505_, _19504_);
  and (_19506_, _16081_, _23718_);
  and (_19507_, _16083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or (_11701_, _19507_, _19506_);
  and (_19508_, _23982_, _23843_);
  and (_19509_, _23845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or (_11703_, _19509_, _19508_);
  and (_11721_, _00538_, _22761_);
  and (_11732_, _16332_, _24847_);
  and (_11734_, _00454_, _22761_);
  and (_19510_, _02069_, _23838_);
  and (_19511_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_27253_, _19511_, _19510_);
  or (_19512_, _02086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_19513_, _19512_, _22761_);
  nand (_19514_, _02086_, _23914_);
  and (_11753_, _19514_, _19513_);
  and (_11755_, _00675_, _22761_);
  and (_11757_, _26372_, _22761_);
  or (_19515_, _03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_11762_, _19515_, _03381_);
  and (_11764_, _00620_, _22761_);
  or (_19516_, _03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_11766_, _19516_, _03399_);
  and (_19517_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_19518_, _17978_, _23791_);
  or (_11774_, _19518_, _19517_);
  and (_19519_, _03340_, _23791_);
  and (_19520_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_11779_, _19520_, _19519_);
  and (_19521_, _03340_, _23635_);
  and (_19522_, _03343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_11784_, _19522_, _19521_);
  and (_19523_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_19524_, _17978_, _23838_);
  or (_27238_, _19524_, _19523_);
  and (_19525_, _03273_, _23635_);
  and (_19526_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_11796_, _19526_, _19525_);
  and (_19527_, _03273_, _23838_);
  and (_19528_, _03275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_11798_, _19528_, _19527_);
  and (_19529_, _02845_, _23676_);
  and (_19530_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_11803_, _19530_, _19529_);
  and (_19531_, _03214_, _23718_);
  and (_19532_, _03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_11808_, _19532_, _19531_);
  and (_19533_, _17979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_19534_, _17978_, _23718_);
  or (_11816_, _19534_, _19533_);
  and (_19535_, _03154_, _23676_);
  and (_19536_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_11837_, _19536_, _19535_);
  and (_19537_, _03189_, _23635_);
  and (_19538_, _03192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_11839_, _19538_, _19537_);
  and (_19539_, _03154_, _23982_);
  and (_19540_, _03156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_11841_, _19540_, _19539_);
  and (_19541_, _02436_, _23718_);
  and (_19542_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or (_27093_, _19542_, _19541_);
  and (_19543_, _03032_, _23755_);
  and (_19544_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_11847_, _19544_, _19543_);
  and (_19545_, _03032_, _23838_);
  and (_19546_, _03034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_27293_, _19546_, _19545_);
  and (_19547_, _05445_, _23676_);
  and (_19548_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  or (_11853_, _19548_, _19547_);
  and (_19549_, _03010_, _23982_);
  and (_19550_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_11856_, _19550_, _19549_);
  and (_19551_, _16707_, _23755_);
  and (_19552_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_11859_, _19552_, _19551_);
  and (_19553_, _02947_, _23718_);
  and (_19554_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_11864_, _19554_, _19553_);
  and (_19555_, _02947_, _23676_);
  and (_19556_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_11869_, _19556_, _19555_);
  and (_19557_, _02947_, _23589_);
  and (_19558_, _02950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_11877_, _19558_, _19557_);
  and (_19559_, _15899_, _23982_);
  and (_19560_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or (_11879_, _19560_, _19559_);
  and (_19561_, _03358_, _23589_);
  and (_19562_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or (_11882_, _19562_, _19561_);
  and (_19563_, _02768_, _23982_);
  and (_19564_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_26945_, _19564_, _19563_);
  and (_19565_, _02768_, _23718_);
  and (_19566_, _02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_11886_, _19566_, _19565_);
  and (_19567_, _02750_, _23718_);
  and (_19568_, _02752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_11888_, _19568_, _19567_);
  and (_19569_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  and (_19570_, _02840_, _23755_);
  or (_11891_, _19570_, _19569_);
  and (_19571_, _25517_, _23635_);
  and (_19572_, _25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_11898_, _19572_, _19571_);
  and (_19573_, _16707_, _23635_);
  and (_19574_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_11911_, _19574_, _19573_);
  and (_19575_, _24777_, _23718_);
  and (_19576_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or (_11913_, _19576_, _19575_);
  and (_19577_, _24777_, _23982_);
  and (_19578_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or (_11915_, _19578_, _19577_);
  and (_19579_, _02092_, _23718_);
  and (_19580_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_11917_, _19580_, _19579_);
  and (_19581_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  and (_19582_, _02840_, _23635_);
  or (_11919_, _19582_, _19581_);
  and (_19583_, _24777_, _23838_);
  and (_19584_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or (_11921_, _19584_, _19583_);
  and (_19585_, _05445_, _23718_);
  and (_19586_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or (_27172_, _19586_, _19585_);
  and (_19587_, _01802_, _23982_);
  and (_19588_, _01804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_27038_, _19588_, _19587_);
  and (_19589_, _15899_, _23755_);
  and (_19590_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or (_11941_, _19590_, _19589_);
  and (_19591_, _25611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or (_11943_, _19591_, _03529_);
  and (_19592_, _25529_, _23838_);
  and (_19593_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_11945_, _19593_, _19592_);
  and (_19594_, _25529_, _23676_);
  and (_19595_, _25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_11947_, _19595_, _19594_);
  and (_19596_, _25468_, _23718_);
  and (_19597_, _25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_11949_, _19597_, _19596_);
  and (_19598_, _02342_, _23791_);
  and (_19599_, _02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_11952_, _19599_, _19598_);
  and (_19600_, _24593_, _23838_);
  and (_19601_, _24595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or (_11955_, _19601_, _19600_);
  and (_19602_, _24584_, _23838_);
  and (_19603_, _24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or (_11957_, _19603_, _19602_);
  and (_19604_, _03296_, _23838_);
  and (_19605_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_11962_, _19605_, _19604_);
  nor (_19606_, _23531_, _26378_);
  and (_19607_, _23531_, _26378_);
  or (_19608_, _19607_, _19606_);
  and (_11972_, _19608_, _22761_);
  and (_19609_, _05445_, _23791_);
  and (_19610_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or (_11974_, _19610_, _19609_);
  and (_11977_, _01204_, _22761_);
  and (_11983_, _00939_, _22761_);
  and (_11985_, _00461_, _22761_);
  and (_11988_, _01057_, _22761_);
  and (_11990_, _01272_, _22761_);
  and (_11992_, _00378_, _22761_);
  and (_11996_, _01342_, _22761_);
  and (_11998_, _26546_, _22761_);
  and (_12000_, _01115_, _22761_);
  and (_12002_, _03846_, _22761_);
  and (_12005_, _00625_, _22761_);
  and (_12009_, _00553_, _22761_);
  and (_12028_, _00682_, _22761_);
  and (_19611_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_19612_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_19613_, _19612_, _19611_);
  and (_19614_, _19613_, _09527_);
  and (_19615_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_19616_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_19617_, _19616_, _19615_);
  and (_19618_, _19617_, _05352_);
  or (_19619_, _19618_, _19614_);
  or (_19620_, _19619_, _09540_);
  and (_19621_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_19622_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_19623_, _19622_, _19621_);
  and (_19624_, _19623_, _09527_);
  and (_19625_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and (_19626_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_19627_, _19626_, _19625_);
  and (_19628_, _19627_, _05352_);
  or (_19629_, _19628_, _19624_);
  or (_19630_, _19629_, _05373_);
  and (_19631_, _19630_, _09566_);
  and (_19632_, _19631_, _19620_);
  or (_19633_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_19634_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_19635_, _19634_, _19633_);
  and (_19636_, _19635_, _09527_);
  or (_19637_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_19638_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and (_19639_, _19638_, _19637_);
  and (_19640_, _19639_, _05352_);
  or (_19641_, _19640_, _19636_);
  or (_19642_, _19641_, _09540_);
  or (_19643_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_19644_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_19645_, _19644_, _19643_);
  and (_19646_, _19645_, _09527_);
  or (_19647_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_19648_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_19649_, _19648_, _19647_);
  and (_19650_, _19649_, _05352_);
  or (_19651_, _19650_, _19646_);
  or (_19652_, _19651_, _05373_);
  and (_19653_, _19652_, _05379_);
  and (_19654_, _19653_, _19642_);
  or (_19655_, _19654_, _19632_);
  and (_19656_, _19655_, _05361_);
  and (_19657_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_19658_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_19659_, _19658_, _19657_);
  and (_19660_, _19659_, _09527_);
  and (_19661_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and (_19662_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_19663_, _19662_, _19661_);
  and (_19664_, _19663_, _05352_);
  or (_19665_, _19664_, _19660_);
  or (_19666_, _19665_, _09540_);
  and (_19667_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_19668_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_19669_, _19668_, _19667_);
  and (_19670_, _19669_, _09527_);
  and (_19671_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_19672_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_19673_, _19672_, _19671_);
  and (_19674_, _19673_, _05352_);
  or (_19675_, _19674_, _19670_);
  or (_19676_, _19675_, _05373_);
  and (_19677_, _19676_, _09566_);
  and (_19678_, _19677_, _19666_);
  or (_19679_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_19680_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_19681_, _19680_, _05352_);
  and (_19682_, _19681_, _19679_);
  or (_19683_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_19684_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_19685_, _19684_, _09527_);
  and (_19686_, _19685_, _19683_);
  or (_19687_, _19686_, _19682_);
  or (_19688_, _19687_, _09540_);
  or (_19689_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_19690_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_19691_, _19690_, _05352_);
  and (_19692_, _19691_, _19689_);
  or (_19693_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_19694_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and (_19695_, _19694_, _09527_);
  and (_19696_, _19695_, _19693_);
  or (_19698_, _19696_, _19692_);
  or (_19699_, _19698_, _05373_);
  and (_19700_, _19699_, _05379_);
  and (_19701_, _19700_, _19688_);
  or (_19702_, _19701_, _19678_);
  and (_19703_, _19702_, _09581_);
  or (_19704_, _19703_, _19656_);
  and (_19705_, _19704_, _09682_);
  and (_19706_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_19707_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_19708_, _19707_, _19706_);
  and (_19709_, _19708_, _09527_);
  and (_19710_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_19711_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_19712_, _19711_, _19710_);
  and (_19713_, _19712_, _05352_);
  or (_19714_, _19713_, _19709_);
  and (_19715_, _19714_, _05373_);
  and (_19716_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_19717_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_19718_, _19717_, _19716_);
  and (_19719_, _19718_, _09527_);
  and (_19720_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_19721_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_19722_, _19721_, _19720_);
  and (_19723_, _19722_, _05352_);
  or (_19724_, _19723_, _19719_);
  and (_19725_, _19724_, _09540_);
  or (_19726_, _19725_, _19715_);
  and (_19727_, _19726_, _09566_);
  or (_19728_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_19729_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_19730_, _19729_, _05352_);
  and (_19731_, _19730_, _19728_);
  or (_19732_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_19733_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_19734_, _19733_, _09527_);
  and (_19735_, _19734_, _19732_);
  or (_19736_, _19735_, _19731_);
  and (_19737_, _19736_, _05373_);
  or (_19738_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_19739_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_19740_, _19739_, _05352_);
  and (_19741_, _19740_, _19738_);
  or (_19742_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_19743_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_19744_, _19743_, _09527_);
  and (_19745_, _19744_, _19742_);
  or (_19746_, _19745_, _19741_);
  and (_19747_, _19746_, _09540_);
  or (_19748_, _19747_, _19737_);
  and (_19749_, _19748_, _05379_);
  or (_19750_, _19749_, _19727_);
  and (_19751_, _19750_, _09581_);
  and (_19752_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_19753_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_19754_, _19753_, _19752_);
  and (_19755_, _19754_, _09527_);
  and (_19756_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_19757_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_19758_, _19757_, _19756_);
  and (_19759_, _19758_, _05352_);
  or (_19760_, _19759_, _19755_);
  and (_19761_, _19760_, _05373_);
  and (_19762_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_19763_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_19764_, _19763_, _19762_);
  and (_19765_, _19764_, _09527_);
  and (_19766_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_19767_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_19768_, _19767_, _19766_);
  and (_19769_, _19768_, _05352_);
  or (_19770_, _19769_, _19765_);
  and (_19771_, _19770_, _09540_);
  or (_19772_, _19771_, _19761_);
  and (_19773_, _19772_, _09566_);
  or (_19774_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_19775_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_19776_, _19775_, _19774_);
  and (_19777_, _19776_, _09527_);
  or (_19778_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_19779_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_19780_, _19779_, _19778_);
  and (_19781_, _19780_, _05352_);
  or (_19782_, _19781_, _19777_);
  and (_19783_, _19782_, _05373_);
  or (_19784_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_19785_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_19786_, _19785_, _19784_);
  and (_19787_, _19786_, _09527_);
  or (_19789_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_19790_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_19791_, _19790_, _19789_);
  and (_19792_, _19791_, _05352_);
  or (_19793_, _19792_, _19787_);
  and (_19794_, _19793_, _09540_);
  or (_19795_, _19794_, _19783_);
  and (_19796_, _19795_, _05379_);
  or (_19797_, _19796_, _19773_);
  and (_19798_, _19797_, _05361_);
  or (_19799_, _19798_, _19751_);
  and (_19800_, _19799_, _05363_);
  or (_19801_, _19800_, _19705_);
  or (_19802_, _19801_, _05357_);
  and (_19803_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and (_19804_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_19805_, _19804_, _19803_);
  and (_19806_, _19805_, _09527_);
  and (_19807_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_19808_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_19809_, _19808_, _19807_);
  and (_19810_, _19809_, _05352_);
  or (_19811_, _19810_, _19806_);
  or (_19812_, _19811_, _09540_);
  and (_19813_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_19814_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_19815_, _19814_, _19813_);
  and (_19816_, _19815_, _09527_);
  and (_19817_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_19818_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_19819_, _19818_, _19817_);
  and (_19820_, _19819_, _05352_);
  or (_19821_, _19820_, _19816_);
  or (_19822_, _19821_, _05373_);
  and (_19823_, _19822_, _09566_);
  and (_19824_, _19823_, _19812_);
  or (_19825_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_19826_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_19827_, _19826_, _05352_);
  and (_19828_, _19827_, _19825_);
  or (_19829_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_19830_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_19831_, _19830_, _09527_);
  and (_19832_, _19831_, _19829_);
  or (_19833_, _19832_, _19828_);
  or (_19834_, _19833_, _09540_);
  or (_19835_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_19836_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_19837_, _19836_, _05352_);
  and (_19838_, _19837_, _19835_);
  or (_19839_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_19840_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and (_19841_, _19840_, _09527_);
  and (_19842_, _19841_, _19839_);
  or (_19843_, _19842_, _19838_);
  or (_19844_, _19843_, _05373_);
  and (_19845_, _19844_, _05379_);
  and (_19846_, _19845_, _19834_);
  or (_19847_, _19846_, _19824_);
  and (_19848_, _19847_, _09581_);
  and (_19849_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_19850_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_19851_, _19850_, _19849_);
  and (_19852_, _19851_, _09527_);
  and (_19853_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_19854_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_19855_, _19854_, _19853_);
  and (_19856_, _19855_, _05352_);
  or (_19857_, _19856_, _19852_);
  or (_19858_, _19857_, _09540_);
  and (_19859_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_19860_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_19861_, _19860_, _19859_);
  and (_19862_, _19861_, _09527_);
  and (_19863_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_19864_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_19865_, _19864_, _19863_);
  and (_19866_, _19865_, _05352_);
  or (_19867_, _19866_, _19862_);
  or (_19868_, _19867_, _05373_);
  and (_19869_, _19868_, _09566_);
  and (_19870_, _19869_, _19858_);
  or (_19871_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_19872_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_19873_, _19872_, _19871_);
  and (_19874_, _19873_, _09527_);
  or (_19875_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_19876_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_19877_, _19876_, _19875_);
  and (_19878_, _19877_, _05352_);
  or (_19879_, _19878_, _19874_);
  or (_19880_, _19879_, _09540_);
  or (_19881_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_19882_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_19883_, _19882_, _19881_);
  and (_19884_, _19883_, _09527_);
  or (_19885_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_19886_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_19887_, _19886_, _19885_);
  and (_19888_, _19887_, _05352_);
  or (_19889_, _19888_, _19884_);
  or (_19890_, _19889_, _05373_);
  and (_19891_, _19890_, _05379_);
  and (_19892_, _19891_, _19880_);
  or (_19893_, _19892_, _19870_);
  and (_19894_, _19893_, _05361_);
  or (_19895_, _19894_, _19848_);
  and (_19896_, _19895_, _09682_);
  or (_19897_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_19898_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and (_19899_, _19898_, _19897_);
  and (_19900_, _19899_, _09527_);
  or (_19901_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_19902_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_19903_, _19902_, _19901_);
  and (_19904_, _19903_, _05352_);
  or (_19905_, _19904_, _19900_);
  and (_19906_, _19905_, _09540_);
  or (_19907_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_19908_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_19909_, _19908_, _19907_);
  and (_19910_, _19909_, _09527_);
  or (_19911_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_19912_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and (_19913_, _19912_, _19911_);
  and (_19914_, _19913_, _05352_);
  or (_19915_, _19914_, _19910_);
  and (_19916_, _19915_, _05373_);
  or (_19917_, _19916_, _19906_);
  and (_19918_, _19917_, _05379_);
  and (_19919_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_19920_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_19921_, _19920_, _19919_);
  and (_19922_, _19921_, _09527_);
  and (_19923_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_19924_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_19925_, _19924_, _19923_);
  and (_19926_, _19925_, _05352_);
  or (_19927_, _19926_, _19922_);
  and (_19928_, _19927_, _09540_);
  and (_19929_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_19930_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_19931_, _19930_, _19929_);
  and (_19932_, _19931_, _09527_);
  and (_19933_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_19934_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_19935_, _19934_, _19933_);
  and (_19936_, _19935_, _05352_);
  or (_19937_, _19936_, _19932_);
  and (_19938_, _19937_, _05373_);
  or (_19940_, _19938_, _19928_);
  and (_19941_, _19940_, _09566_);
  or (_19942_, _19941_, _19918_);
  and (_19943_, _19942_, _05361_);
  or (_19944_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_19945_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and (_19946_, _19945_, _05352_);
  and (_19947_, _19946_, _19944_);
  or (_19948_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_19949_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and (_19950_, _19949_, _09527_);
  and (_19951_, _19950_, _19948_);
  or (_19952_, _19951_, _19947_);
  and (_19953_, _19952_, _09540_);
  or (_19954_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_19955_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and (_19956_, _19955_, _05352_);
  and (_19957_, _19956_, _19954_);
  or (_19958_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_19959_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and (_19960_, _19959_, _09527_);
  and (_19961_, _19960_, _19958_);
  or (_19962_, _19961_, _19957_);
  and (_19963_, _19962_, _05373_);
  or (_19964_, _19963_, _19953_);
  and (_19965_, _19964_, _05379_);
  and (_19966_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and (_19967_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_19968_, _19967_, _19966_);
  and (_19969_, _19968_, _09527_);
  and (_19970_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and (_19971_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_19972_, _19971_, _19970_);
  and (_19973_, _19972_, _05352_);
  or (_19974_, _19973_, _19969_);
  and (_19975_, _19974_, _09540_);
  and (_19976_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and (_19977_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_19978_, _19977_, _19976_);
  and (_19979_, _19978_, _09527_);
  and (_19980_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and (_19981_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_19982_, _19981_, _19980_);
  and (_19983_, _19982_, _05352_);
  or (_19984_, _19983_, _19979_);
  and (_19985_, _19984_, _05373_);
  or (_19986_, _19985_, _19975_);
  and (_19987_, _19986_, _09566_);
  or (_19988_, _19987_, _19965_);
  and (_19989_, _19988_, _09581_);
  or (_19990_, _19989_, _19943_);
  and (_19991_, _19990_, _05363_);
  or (_19992_, _19991_, _19896_);
  or (_19993_, _19992_, _09739_);
  and (_19994_, _19993_, _19802_);
  or (_19995_, _19994_, _26838_);
  and (_19996_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_19997_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_19998_, _19997_, _19996_);
  and (_19999_, _19998_, _09527_);
  and (_20000_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_20001_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_20002_, _20001_, _20000_);
  and (_20003_, _20002_, _05352_);
  or (_20004_, _20003_, _19999_);
  or (_20005_, _20004_, _09540_);
  and (_20006_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_20007_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_20008_, _20007_, _20006_);
  and (_20009_, _20008_, _09527_);
  and (_20010_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_20011_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_20012_, _20011_, _20010_);
  and (_20013_, _20012_, _05352_);
  or (_20014_, _20013_, _20009_);
  or (_20015_, _20014_, _05373_);
  and (_20016_, _20015_, _09566_);
  and (_20017_, _20016_, _20005_);
  or (_20018_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_20019_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_20020_, _20019_, _20018_);
  and (_20021_, _20020_, _09527_);
  or (_20022_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_20023_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_20024_, _20023_, _20022_);
  and (_20025_, _20024_, _05352_);
  or (_20026_, _20025_, _20021_);
  or (_20027_, _20026_, _09540_);
  or (_20028_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_20029_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_20030_, _20029_, _20028_);
  and (_20031_, _20030_, _09527_);
  or (_20032_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_20033_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_20034_, _20033_, _20032_);
  and (_20035_, _20034_, _05352_);
  or (_20036_, _20035_, _20031_);
  or (_20037_, _20036_, _05373_);
  and (_20038_, _20037_, _05379_);
  and (_20039_, _20038_, _20027_);
  or (_20040_, _20039_, _20017_);
  and (_20041_, _20040_, _05361_);
  and (_20042_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_20043_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_20044_, _20043_, _20042_);
  and (_20045_, _20044_, _09527_);
  and (_20046_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_20047_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_20048_, _20047_, _20046_);
  and (_20049_, _20048_, _05352_);
  or (_20050_, _20049_, _20045_);
  or (_20051_, _20050_, _09540_);
  and (_20052_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_20053_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_20054_, _20053_, _20052_);
  and (_20055_, _20054_, _09527_);
  and (_20056_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_20057_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_20058_, _20057_, _20056_);
  and (_20059_, _20058_, _05352_);
  or (_20060_, _20059_, _20055_);
  or (_20061_, _20060_, _05373_);
  and (_20062_, _20061_, _09566_);
  and (_20063_, _20062_, _20051_);
  or (_20064_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_20065_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_20066_, _20065_, _05352_);
  and (_20067_, _20066_, _20064_);
  or (_20068_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_20069_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_20070_, _20069_, _09527_);
  and (_20071_, _20070_, _20068_);
  or (_20072_, _20071_, _20067_);
  or (_20073_, _20072_, _09540_);
  or (_20074_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_20075_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_20076_, _20075_, _05352_);
  and (_20077_, _20076_, _20074_);
  or (_20078_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_20079_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_20080_, _20079_, _09527_);
  and (_20081_, _20080_, _20078_);
  or (_20082_, _20081_, _20077_);
  or (_20083_, _20082_, _05373_);
  and (_20084_, _20083_, _05379_);
  and (_20085_, _20084_, _20073_);
  or (_20086_, _20085_, _20063_);
  and (_20087_, _20086_, _09581_);
  or (_20088_, _20087_, _20041_);
  and (_20089_, _20088_, _09682_);
  and (_20090_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_20091_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_20092_, _20091_, _20090_);
  and (_20093_, _20092_, _09527_);
  and (_20094_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_20095_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_20096_, _20095_, _20094_);
  and (_20097_, _20096_, _05352_);
  or (_20098_, _20097_, _20093_);
  and (_20099_, _20098_, _05373_);
  and (_20100_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_20101_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_20102_, _20101_, _20100_);
  and (_20103_, _20102_, _09527_);
  and (_20104_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_20105_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_20106_, _20105_, _20104_);
  and (_20107_, _20106_, _05352_);
  or (_20108_, _20107_, _20103_);
  and (_20109_, _20108_, _09540_);
  or (_20110_, _20109_, _20099_);
  and (_20111_, _20110_, _09566_);
  or (_20112_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_20113_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_20114_, _20113_, _05352_);
  and (_20115_, _20114_, _20112_);
  or (_20116_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_20117_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_20118_, _20117_, _09527_);
  and (_20119_, _20118_, _20116_);
  or (_20120_, _20119_, _20115_);
  and (_20121_, _20120_, _05373_);
  or (_20122_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_20123_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_20124_, _20123_, _05352_);
  and (_20125_, _20124_, _20122_);
  or (_20126_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_20127_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_20128_, _20127_, _09527_);
  and (_20129_, _20128_, _20126_);
  or (_20130_, _20129_, _20125_);
  and (_20131_, _20130_, _09540_);
  or (_20132_, _20131_, _20121_);
  and (_20133_, _20132_, _05379_);
  or (_20134_, _20133_, _20111_);
  and (_20135_, _20134_, _09581_);
  and (_20136_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_20137_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_20138_, _20137_, _20136_);
  and (_20139_, _20138_, _09527_);
  and (_20140_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_20141_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_20142_, _20141_, _20140_);
  and (_20143_, _20142_, _05352_);
  or (_20144_, _20143_, _20139_);
  and (_20145_, _20144_, _05373_);
  and (_20146_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_20147_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_20148_, _20147_, _20146_);
  and (_20149_, _20148_, _09527_);
  and (_20150_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_20151_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_20152_, _20151_, _20150_);
  and (_20153_, _20152_, _05352_);
  or (_20154_, _20153_, _20149_);
  and (_20155_, _20154_, _09540_);
  or (_20156_, _20155_, _20145_);
  and (_20157_, _20156_, _09566_);
  or (_20158_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_20159_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_20160_, _20159_, _20158_);
  and (_20161_, _20160_, _09527_);
  or (_20162_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_20163_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_20164_, _20163_, _20162_);
  and (_20165_, _20164_, _05352_);
  or (_20166_, _20165_, _20161_);
  and (_20167_, _20166_, _05373_);
  or (_20168_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_20169_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_20170_, _20169_, _20168_);
  and (_20171_, _20170_, _09527_);
  or (_20172_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_20173_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_20174_, _20173_, _20172_);
  and (_20175_, _20174_, _05352_);
  or (_20176_, _20175_, _20171_);
  and (_20177_, _20176_, _09540_);
  or (_20178_, _20177_, _20167_);
  and (_20179_, _20178_, _05379_);
  or (_20180_, _20179_, _20157_);
  and (_20181_, _20180_, _05361_);
  or (_20182_, _20181_, _20135_);
  and (_20183_, _20182_, _05363_);
  or (_20184_, _20183_, _20089_);
  or (_20185_, _20184_, _05357_);
  and (_20186_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_20187_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_20188_, _20187_, _20186_);
  and (_20189_, _20188_, _09527_);
  and (_20190_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_20191_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_20192_, _20191_, _20190_);
  and (_20193_, _20192_, _05352_);
  or (_20194_, _20193_, _20189_);
  or (_20195_, _20194_, _09540_);
  and (_20196_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_20197_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_20198_, _20197_, _20196_);
  and (_20199_, _20198_, _09527_);
  and (_20200_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_20201_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_20202_, _20201_, _20200_);
  and (_20203_, _20202_, _05352_);
  or (_20204_, _20203_, _20199_);
  or (_20205_, _20204_, _05373_);
  and (_20206_, _20205_, _09566_);
  and (_20207_, _20206_, _20195_);
  or (_20208_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_20209_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_20211_, _20209_, _05352_);
  and (_20212_, _20211_, _20208_);
  or (_20213_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_20214_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_20215_, _20214_, _09527_);
  and (_20216_, _20215_, _20213_);
  or (_20217_, _20216_, _20212_);
  or (_20218_, _20217_, _09540_);
  or (_20219_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_20220_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_20221_, _20220_, _05352_);
  and (_20222_, _20221_, _20219_);
  or (_20223_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_20224_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_20225_, _20224_, _09527_);
  and (_20226_, _20225_, _20223_);
  or (_20227_, _20226_, _20222_);
  or (_20228_, _20227_, _05373_);
  and (_20229_, _20228_, _05379_);
  and (_20230_, _20229_, _20218_);
  or (_20231_, _20230_, _20207_);
  and (_20232_, _20231_, _09581_);
  and (_20233_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_20234_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_20235_, _20234_, _20233_);
  and (_20236_, _20235_, _09527_);
  and (_20237_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_20238_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_20239_, _20238_, _20237_);
  and (_20240_, _20239_, _05352_);
  or (_20241_, _20240_, _20236_);
  or (_20242_, _20241_, _09540_);
  and (_20243_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_20244_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_20245_, _20244_, _20243_);
  and (_20246_, _20245_, _09527_);
  and (_20247_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_20248_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_20249_, _20248_, _20247_);
  and (_20250_, _20249_, _05352_);
  or (_20251_, _20250_, _20246_);
  or (_20252_, _20251_, _05373_);
  and (_20253_, _20252_, _09566_);
  and (_20254_, _20253_, _20242_);
  or (_20255_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_20256_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_20257_, _20256_, _20255_);
  and (_20258_, _20257_, _09527_);
  or (_20259_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_20260_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_20261_, _20260_, _20259_);
  and (_20262_, _20261_, _05352_);
  or (_20263_, _20262_, _20258_);
  or (_20264_, _20263_, _09540_);
  or (_20265_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_20266_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_20267_, _20266_, _20265_);
  and (_20268_, _20267_, _09527_);
  or (_20269_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_20270_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_20271_, _20270_, _20269_);
  and (_20272_, _20271_, _05352_);
  or (_20273_, _20272_, _20268_);
  or (_20274_, _20273_, _05373_);
  and (_20275_, _20274_, _05379_);
  and (_20276_, _20275_, _20264_);
  or (_20277_, _20276_, _20254_);
  and (_20278_, _20277_, _05361_);
  or (_20279_, _20278_, _20232_);
  and (_20280_, _20279_, _09682_);
  or (_20281_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_20282_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_20283_, _20282_, _20281_);
  and (_20284_, _20283_, _09527_);
  or (_20285_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_20286_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_20287_, _20286_, _20285_);
  and (_20288_, _20287_, _05352_);
  or (_20289_, _20288_, _20284_);
  and (_20290_, _20289_, _09540_);
  or (_20291_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_20292_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_20293_, _20292_, _20291_);
  and (_20294_, _20293_, _09527_);
  or (_20295_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_20296_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_20297_, _20296_, _20295_);
  and (_20298_, _20297_, _05352_);
  or (_20299_, _20298_, _20294_);
  and (_20300_, _20299_, _05373_);
  or (_20301_, _20300_, _20290_);
  and (_20302_, _20301_, _05379_);
  and (_20303_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_20304_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_20305_, _20304_, _20303_);
  and (_20306_, _20305_, _09527_);
  and (_20307_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_20308_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_20309_, _20308_, _20307_);
  and (_20310_, _20309_, _05352_);
  or (_20311_, _20310_, _20306_);
  and (_20312_, _20311_, _09540_);
  and (_20313_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_20314_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_20315_, _20314_, _20313_);
  and (_20316_, _20315_, _09527_);
  and (_20317_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_20318_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_20319_, _20318_, _20317_);
  and (_20320_, _20319_, _05352_);
  or (_20321_, _20320_, _20316_);
  and (_20322_, _20321_, _05373_);
  or (_20323_, _20322_, _20312_);
  and (_20324_, _20323_, _09566_);
  or (_20325_, _20324_, _20302_);
  and (_20326_, _20325_, _05361_);
  or (_20327_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_20328_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_20329_, _20328_, _05352_);
  and (_20330_, _20329_, _20327_);
  or (_20331_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_20332_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_20333_, _20332_, _09527_);
  and (_20334_, _20333_, _20331_);
  or (_20335_, _20334_, _20330_);
  and (_20336_, _20335_, _09540_);
  or (_20337_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_20338_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_20339_, _20338_, _05352_);
  and (_20340_, _20339_, _20337_);
  or (_20341_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_20342_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_20343_, _20342_, _09527_);
  and (_20344_, _20343_, _20341_);
  or (_20345_, _20344_, _20340_);
  and (_20346_, _20345_, _05373_);
  or (_20347_, _20346_, _20336_);
  and (_20348_, _20347_, _05379_);
  and (_20349_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_20350_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_20351_, _20350_, _20349_);
  and (_20352_, _20351_, _09527_);
  and (_20353_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_20354_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_20355_, _20354_, _20353_);
  and (_20356_, _20355_, _05352_);
  or (_20357_, _20356_, _20352_);
  and (_20358_, _20357_, _09540_);
  and (_20359_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_20360_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_20361_, _20360_, _20359_);
  and (_20362_, _20361_, _09527_);
  and (_20363_, _09530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_20364_, _05388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_20365_, _20364_, _20363_);
  and (_20366_, _20365_, _05352_);
  or (_20367_, _20366_, _20362_);
  and (_20368_, _20367_, _05373_);
  or (_20369_, _20368_, _20358_);
  and (_20370_, _20369_, _09566_);
  or (_20371_, _20370_, _20348_);
  and (_20372_, _20371_, _09581_);
  or (_20373_, _20372_, _20326_);
  and (_20374_, _20373_, _05363_);
  or (_20375_, _20374_, _20280_);
  or (_20376_, _20375_, _09739_);
  and (_20377_, _20376_, _20185_);
  or (_20378_, _20377_, _04360_);
  and (_20379_, _20378_, _19995_);
  or (_20380_, _20379_, _05401_);
  or (_20381_, _10445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_20382_, _20381_, _22761_);
  and (_12045_, _20382_, _20380_);
  and (_20383_, _17001_, _23755_);
  and (_20384_, _17003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or (_12096_, _20384_, _20383_);
  and (_20385_, _24119_, _23589_);
  and (_20386_, _24121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_12109_, _20386_, _20385_);
  nor (_26896_[4], _00136_, rst);
  nor (_26896_[5], _00021_, rst);
  and (_20387_, _15899_, _23791_);
  and (_20388_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or (_12153_, _20388_, _20387_);
  and (_20389_, _02845_, _23755_);
  and (_20390_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_27277_, _20390_, _20389_);
  and (_20391_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and (_20392_, _02858_, _23589_);
  or (_12158_, _20392_, _20391_);
  and (_20393_, _12516_, _23635_);
  and (_20394_, _12519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or (_12160_, _20394_, _20393_);
  and (_20395_, _02069_, _23755_);
  and (_20396_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_12162_, _20396_, _20395_);
  and (_20397_, _17972_, _23676_);
  and (_20398_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_12164_, _20398_, _20397_);
  and (_20399_, _02785_, _23589_);
  and (_20401_, _02787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or (_12167_, _20401_, _20399_);
  and (_20402_, _15899_, _23676_);
  and (_20403_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or (_12169_, _20403_, _20402_);
  and (_20404_, _02069_, _23589_);
  and (_20405_, _02071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_12172_, _20405_, _20404_);
  and (_20406_, _15995_, _23718_);
  and (_20407_, _15997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or (_26993_, _20407_, _20406_);
  and (_20408_, _02859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_20409_, _02858_, _23755_);
  or (_12175_, _20409_, _20408_);
  and (_20410_, _03358_, _23718_);
  and (_20411_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or (_27168_, _20411_, _20410_);
  and (_20412_, _02436_, _23982_);
  and (_20413_, _02438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or (_12186_, _20413_, _20412_);
  and (_20414_, _02845_, _23635_);
  and (_20415_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_27276_, _20415_, _20414_);
  and (_20416_, _15899_, _23718_);
  and (_20417_, _15901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or (_12191_, _20417_, _20416_);
  and (_20418_, _03358_, _23982_);
  and (_20419_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or (_12198_, _20419_, _20418_);
  and (_20420_, _06255_, _23718_);
  and (_20421_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or (_12211_, _20421_, _20420_);
  and (_12219_, _01001_, _22761_);
  and (_20422_, _15909_, _23635_);
  and (_20423_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_12371_, _20423_, _20422_);
  and (_20424_, _13736_, _23718_);
  and (_20425_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_12404_, _20425_, _20424_);
  and (_20426_, _15909_, _23982_);
  and (_20427_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_12423_, _20427_, _20426_);
  and (_20428_, _13696_, _23755_);
  and (_20429_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or (_27171_, _20429_, _20428_);
  and (_20430_, _17972_, _23838_);
  and (_20431_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_12434_, _20431_, _20430_);
  and (_20432_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20433_, _20432_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20434_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_20435_, _20434_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_20436_, _20435_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_20437_, _20436_, _20433_);
  and (_20438_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_20439_, _20438_, _20437_);
  and (_20440_, _20439_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_20441_, _20440_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_20442_, _20441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_20443_, _20442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_20444_, _20443_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20445_, _20443_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20446_, _20445_, _20444_);
  nor (_20447_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20448_, _20447_);
  nor (_20449_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20450_, _22798_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20451_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _22794_);
  nor (_20452_, _20451_, _20450_);
  and (_20453_, _20452_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20454_, _20453_, _20449_);
  not (_20455_, _20454_);
  and (_20456_, _20432_, _22802_);
  nor (_20457_, _20432_, _22802_);
  nor (_20458_, _20457_, _20456_);
  nor (_20459_, _20458_, _22789_);
  and (_20460_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _22789_);
  nor (_20461_, _20460_, _20459_);
  nor (_20462_, _20461_, _05456_);
  and (_20463_, _20461_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_20464_, _20463_, _20462_);
  nor (_20465_, _20464_, _20455_);
  and (_20466_, _20461_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_20467_, _20461_, _05493_);
  nor (_20468_, _20467_, _20466_);
  nor (_20469_, _20468_, _20454_);
  nor (_20470_, _20469_, _20465_);
  nor (_20471_, _20470_, _20448_);
  and (_20472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _22789_);
  not (_20473_, _20472_);
  not (_20474_, _20461_);
  nor (_20475_, _20454_, _05479_);
  and (_20476_, _20454_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_20477_, _20476_, _20475_);
  nor (_20478_, _20477_, _20474_);
  nor (_20479_, _20454_, _06111_);
  and (_20480_, _20454_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_20481_, _20480_, _20479_);
  nor (_20482_, _20481_, _20461_);
  nor (_20483_, _20482_, _20478_);
  nor (_20484_, _20483_, _20473_);
  nor (_20485_, _20484_, _20471_);
  and (_20486_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20487_, _20486_);
  not (_20488_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_20489_, _20454_, _20488_);
  and (_20490_, _20454_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_20491_, _20490_, _20489_);
  nor (_20492_, _20491_, _20474_);
  nor (_20493_, _20454_, _05526_);
  and (_20494_, _20454_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_20495_, _20494_, _20493_);
  nor (_20496_, _20495_, _20461_);
  nor (_20497_, _20496_, _20492_);
  nor (_20498_, _20497_, _20487_);
  and (_20499_, _22794_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20500_, _20499_);
  nor (_20501_, _20461_, _05504_);
  and (_20502_, _20461_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_20503_, _20502_, _20501_);
  nor (_20504_, _20503_, _20455_);
  nor (_20505_, _20461_, _06073_);
  and (_20506_, _20461_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_20507_, _20506_, _20505_);
  nor (_20508_, _20507_, _20454_);
  nor (_20509_, _20508_, _20504_);
  nor (_20510_, _20509_, _20500_);
  nor (_20511_, _20510_, _20498_);
  and (_20512_, _20511_, _20485_);
  and (_20513_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_20514_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_20515_, _20514_, _20513_);
  and (_20516_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_20517_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_20518_, _20517_, _20516_);
  and (_20519_, _20518_, _20515_);
  and (_20520_, _20519_, _20455_);
  and (_20521_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_20522_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_20523_, _20522_, _20521_);
  and (_20524_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_20525_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_20526_, _20525_, _20524_);
  and (_20527_, _20526_, _20523_);
  and (_20528_, _20527_, _20454_);
  or (_20529_, _20528_, _20474_);
  nor (_20530_, _20529_, _20520_);
  and (_20531_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_20532_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_20533_, _20532_, _20531_);
  and (_20534_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_20535_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_20536_, _20535_, _20534_);
  and (_20537_, _20536_, _20533_);
  nor (_20538_, _20537_, _20454_);
  and (_20539_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_20540_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_20541_, _20540_, _20539_);
  and (_20542_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_20543_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_20544_, _20543_, _20542_);
  and (_20545_, _20544_, _20541_);
  nor (_20546_, _20545_, _20455_);
  or (_20547_, _20546_, _20538_);
  and (_20548_, _20547_, _20474_);
  nor (_20549_, _20548_, _20530_);
  nor (_20550_, _20549_, _20512_);
  and (_20551_, _20550_, _20446_);
  nor (_20552_, _20550_, _20446_);
  nor (_20553_, _20552_, _20551_);
  and (_20554_, _20442_, _22844_);
  nor (_20555_, _20442_, _22844_);
  nor (_20556_, _20555_, _20554_);
  not (_20557_, _20556_);
  and (_20558_, _20557_, _20550_);
  nor (_20559_, _20557_, _20550_);
  nor (_20560_, _20441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20561_, _20560_, _20442_);
  and (_20562_, _20561_, _20550_);
  nor (_20563_, _20440_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_20564_, _20563_, _20441_);
  and (_20565_, _20564_, _20550_);
  nor (_20566_, _20564_, _20550_);
  nor (_20567_, _20439_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_20568_, _20567_, _20440_);
  and (_20569_, _20568_, _20550_);
  nor (_20570_, _20568_, _20550_);
  nor (_20571_, _20570_, _20569_);
  not (_20572_, _20571_);
  and (_20573_, _20437_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20574_, _20573_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_20575_, _20574_, _20439_);
  and (_20576_, _20575_, _20550_);
  nor (_20577_, _20437_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20578_, _20577_, _20573_);
  and (_20579_, _20578_, _20550_);
  nor (_20580_, _20575_, _20550_);
  nor (_20581_, _20580_, _20576_);
  and (_20582_, _20435_, _20433_);
  nor (_20583_, _20582_, _22820_);
  and (_20584_, _20582_, _22820_);
  nor (_20585_, _20584_, _20583_);
  not (_20586_, _20585_);
  and (_20587_, _20586_, _20550_);
  nor (_20588_, _20586_, _20550_);
  and (_20589_, _20434_, _20433_);
  nor (_20590_, _20589_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_20591_, _20590_, _20582_);
  and (_20592_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_20593_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_20594_, _20593_, _20592_);
  and (_20595_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_20596_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_20597_, _20596_, _20595_);
  and (_20598_, _20597_, _20594_);
  and (_20599_, _20598_, _20455_);
  and (_20600_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_20601_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_20602_, _20601_, _20600_);
  and (_20603_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_20604_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_20605_, _20604_, _20603_);
  and (_20606_, _20605_, _20602_);
  and (_20607_, _20606_, _20454_);
  or (_20608_, _20607_, _20474_);
  nor (_20609_, _20608_, _20599_);
  and (_20610_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_20611_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_20612_, _20611_, _20610_);
  and (_20613_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_20614_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_20615_, _20614_, _20613_);
  and (_20616_, _20615_, _20612_);
  nor (_20617_, _20616_, _20454_);
  and (_20618_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_20619_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_20620_, _20619_, _20618_);
  and (_20621_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_20622_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_20623_, _20622_, _20621_);
  and (_20624_, _20623_, _20620_);
  nor (_20625_, _20624_, _20455_);
  or (_20626_, _20625_, _20617_);
  and (_20627_, _20626_, _20474_);
  nor (_20628_, _20627_, _20609_);
  nor (_20629_, _20628_, _20512_);
  and (_20630_, _20629_, _20591_);
  nor (_20631_, _20629_, _20591_);
  nor (_20632_, _20631_, _20630_);
  not (_20633_, _20632_);
  and (_20634_, _20433_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20635_, _20634_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_20636_, _20635_, _20589_);
  and (_20637_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_20638_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_20639_, _20638_, _20637_);
  and (_20640_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_20641_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_20642_, _20641_, _20640_);
  and (_20643_, _20642_, _20639_);
  and (_20644_, _20643_, _20455_);
  and (_20645_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_20646_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_20647_, _20646_, _20645_);
  and (_20648_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_20649_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_20650_, _20649_, _20648_);
  and (_20651_, _20650_, _20647_);
  and (_20652_, _20651_, _20454_);
  or (_20653_, _20652_, _20474_);
  nor (_20654_, _20653_, _20644_);
  and (_20655_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_20656_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_20657_, _20656_, _20655_);
  and (_20658_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_20659_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_20660_, _20659_, _20658_);
  and (_20661_, _20660_, _20657_);
  nor (_20662_, _20661_, _20454_);
  and (_20663_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_20664_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_20665_, _20664_, _20663_);
  and (_20666_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_20667_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_20668_, _20667_, _20666_);
  and (_20669_, _20668_, _20665_);
  nor (_20670_, _20669_, _20455_);
  or (_20671_, _20670_, _20662_);
  and (_20672_, _20671_, _20474_);
  nor (_20673_, _20672_, _20654_);
  nor (_20674_, _20673_, _20512_);
  and (_20675_, _20674_, _20636_);
  nor (_20676_, _20674_, _20636_);
  nor (_20677_, _20676_, _20675_);
  not (_20678_, _20677_);
  and (_20679_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_20680_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_20681_, _20680_, _20679_);
  and (_20682_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_20683_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_20684_, _20683_, _20682_);
  and (_20685_, _20684_, _20681_);
  and (_20686_, _20685_, _20455_);
  and (_20687_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_20688_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_20689_, _20688_, _20687_);
  and (_20690_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_20691_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_20692_, _20691_, _20690_);
  and (_20693_, _20692_, _20689_);
  and (_20694_, _20693_, _20454_);
  or (_20695_, _20694_, _20474_);
  nor (_20696_, _20695_, _20686_);
  and (_20697_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_20698_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_20699_, _20698_, _20697_);
  and (_20700_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_20701_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_20702_, _20701_, _20700_);
  and (_20703_, _20702_, _20699_);
  and (_20704_, _20703_, _20455_);
  and (_20705_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_20706_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_20707_, _20706_, _20705_);
  and (_20708_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_20709_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_20710_, _20709_, _20708_);
  and (_20711_, _20710_, _20707_);
  and (_20712_, _20711_, _20454_);
  or (_20713_, _20712_, _20461_);
  nor (_20714_, _20713_, _20704_);
  nor (_20715_, _20714_, _20696_);
  nor (_20716_, _20715_, _20512_);
  nor (_20717_, _20433_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20718_, _20717_, _20634_);
  and (_20719_, _20718_, _20716_);
  not (_20720_, _20458_);
  and (_20721_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_20722_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_20723_, _20722_, _20721_);
  and (_20724_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_20725_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_20726_, _20725_, _20724_);
  and (_20727_, _20726_, _20723_);
  and (_20728_, _20727_, _20455_);
  and (_20729_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_20730_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_20731_, _20730_, _20729_);
  and (_20732_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_20733_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_20734_, _20733_, _20732_);
  and (_20735_, _20734_, _20731_);
  and (_20736_, _20735_, _20454_);
  or (_20737_, _20736_, _20461_);
  nor (_20738_, _20737_, _20728_);
  and (_20739_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_20740_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_20741_, _20740_, _20739_);
  and (_20742_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_20743_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_20744_, _20743_, _20742_);
  and (_20745_, _20744_, _20741_);
  and (_20746_, _20745_, _20455_);
  and (_20747_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_20748_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_20749_, _20748_, _20747_);
  and (_20750_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_20751_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_20752_, _20751_, _20750_);
  and (_20753_, _20752_, _20749_);
  and (_20754_, _20753_, _20454_);
  or (_20755_, _20754_, _20474_);
  nor (_20756_, _20755_, _20746_);
  nor (_20757_, _20756_, _20738_);
  nor (_20758_, _20757_, _20512_);
  and (_20759_, _20758_, _20720_);
  nor (_20760_, _20758_, _20720_);
  nor (_20761_, _20760_, _20759_);
  not (_20762_, _20761_);
  not (_20763_, _20452_);
  and (_20764_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_20765_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_20766_, _20765_, _20764_);
  and (_20767_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_20768_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_20769_, _20768_, _20767_);
  and (_20770_, _20769_, _20766_);
  and (_20771_, _20770_, _20455_);
  and (_20772_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_20773_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_20774_, _20773_, _20772_);
  and (_20775_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_20776_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_20777_, _20776_, _20775_);
  and (_20778_, _20777_, _20774_);
  and (_20779_, _20778_, _20454_);
  or (_20780_, _20779_, _20461_);
  nor (_20781_, _20780_, _20771_);
  and (_20782_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_20783_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_20784_, _20783_, _20782_);
  and (_20785_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_20786_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_20787_, _20786_, _20785_);
  and (_20788_, _20787_, _20784_);
  nor (_20789_, _20788_, _20454_);
  and (_20790_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_20791_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_20792_, _20791_, _20790_);
  and (_20793_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_20794_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_20795_, _20794_, _20793_);
  and (_20796_, _20795_, _20792_);
  nor (_20797_, _20796_, _20455_);
  or (_20798_, _20797_, _20789_);
  and (_20799_, _20798_, _20461_);
  nor (_20800_, _20799_, _20781_);
  nor (_20801_, _20800_, _20512_);
  and (_20802_, _20801_, _20763_);
  and (_20803_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_20804_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_20805_, _20804_, _20803_);
  and (_20806_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_20807_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_20808_, _20807_, _20806_);
  and (_20809_, _20808_, _20805_);
  and (_20810_, _20809_, _20455_);
  and (_20811_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_20812_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_20813_, _20812_, _20811_);
  and (_20814_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_20815_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_20816_, _20815_, _20814_);
  and (_20817_, _20816_, _20813_);
  and (_20818_, _20817_, _20454_);
  or (_20819_, _20818_, _20474_);
  nor (_20820_, _20819_, _20810_);
  and (_20821_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_20822_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_20823_, _20822_, _20821_);
  and (_20824_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_20825_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_20826_, _20825_, _20824_);
  and (_20827_, _20826_, _20823_);
  nor (_20828_, _20827_, _20454_);
  and (_20829_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_20830_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_20831_, _20830_, _20829_);
  and (_20832_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_20833_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_20834_, _20833_, _20832_);
  and (_20835_, _20834_, _20831_);
  nor (_20836_, _20835_, _20455_);
  or (_20837_, _20836_, _20828_);
  and (_20838_, _20837_, _20474_);
  nor (_20839_, _20838_, _20820_);
  nor (_20840_, _20839_, _20512_);
  and (_20841_, _20840_, _22794_);
  and (_20842_, _20472_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_20843_, _20447_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_20844_, _20843_, _20842_);
  and (_20845_, _20499_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_20846_, _20486_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_20847_, _20846_, _20845_);
  and (_20848_, _20847_, _20844_);
  and (_20849_, _20848_, _20455_);
  and (_20850_, _20472_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_20851_, _20486_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_20852_, _20851_, _20850_);
  and (_20853_, _20499_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_20854_, _20447_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_20855_, _20854_, _20853_);
  and (_20856_, _20855_, _20852_);
  and (_20857_, _20856_, _20454_);
  or (_20858_, _20857_, _20474_);
  nor (_20859_, _20858_, _20849_);
  and (_20860_, _20472_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_20861_, _20486_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_20862_, _20861_, _20860_);
  and (_20863_, _20499_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_20864_, _20447_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_20865_, _20864_, _20863_);
  and (_20866_, _20865_, _20862_);
  nor (_20867_, _20866_, _20454_);
  and (_20868_, _20499_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_20869_, _20486_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_20870_, _20869_, _20868_);
  and (_20871_, _20472_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_20872_, _20447_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_20873_, _20872_, _20871_);
  and (_20874_, _20873_, _20870_);
  nor (_20875_, _20874_, _20455_);
  or (_20876_, _20875_, _20867_);
  and (_20877_, _20876_, _20474_);
  nor (_20878_, _20877_, _20859_);
  nor (_20879_, _20878_, _20512_);
  and (_20880_, _20879_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20881_, _20840_, _22794_);
  nor (_20882_, _20881_, _20841_);
  and (_20883_, _20882_, _20880_);
  nor (_20884_, _20883_, _20841_);
  nor (_20885_, _20801_, _20763_);
  nor (_20886_, _20885_, _20802_);
  not (_20887_, _20886_);
  nor (_20888_, _20887_, _20884_);
  nor (_20889_, _20888_, _20802_);
  nor (_20890_, _20889_, _20762_);
  nor (_20891_, _20890_, _20759_);
  nor (_20892_, _20718_, _20716_);
  nor (_20893_, _20892_, _20719_);
  not (_20894_, _20893_);
  nor (_20895_, _20894_, _20891_);
  nor (_20896_, _20895_, _20719_);
  nor (_20897_, _20896_, _20678_);
  nor (_20898_, _20897_, _20675_);
  nor (_20899_, _20898_, _20633_);
  nor (_20900_, _20899_, _20630_);
  nor (_20901_, _20900_, _20588_);
  or (_20902_, _20901_, _20587_);
  nor (_20903_, _20578_, _20550_);
  nor (_20904_, _20903_, _20579_);
  and (_20905_, _20904_, _20902_);
  and (_20906_, _20905_, _20581_);
  or (_20907_, _20906_, _20579_);
  nor (_20908_, _20907_, _20576_);
  nor (_20909_, _20908_, _20572_);
  nor (_20910_, _20909_, _20569_);
  nor (_20911_, _20910_, _20566_);
  or (_20912_, _20911_, _20565_);
  nor (_20913_, _20561_, _20550_);
  nor (_20914_, _20913_, _20562_);
  and (_20915_, _20914_, _20912_);
  nor (_20916_, _20915_, _20562_);
  nor (_20917_, _20916_, _20559_);
  or (_20918_, _20917_, _20558_);
  and (_20919_, _20918_, _20553_);
  nor (_20920_, _20918_, _20553_);
  nor (_20921_, _20920_, _20919_);
  nand (_20922_, _20921_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_20923_, _20921_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_20924_, _20923_, _20922_);
  nor (_20925_, _20919_, _20551_);
  not (_20926_, _20925_);
  nor (_20927_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_20928_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_20929_, _20928_, _20927_);
  not (_20930_, _20929_);
  and (_20931_, _20930_, _20444_);
  nor (_20932_, _20930_, _20444_);
  nor (_20933_, _20932_, _20931_);
  nor (_20934_, _20933_, _20550_);
  and (_20935_, _20933_, _20550_);
  nor (_20936_, _20935_, _20934_);
  nor (_20937_, _20936_, _20926_);
  and (_20938_, _20936_, _20926_);
  nor (_20939_, _20556_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_20940_, _20556_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_20941_, _20940_, _20939_);
  not (_20942_, _20941_);
  and (_20943_, _20942_, _20550_);
  nor (_20944_, _20942_, _20550_);
  nor (_20945_, _20944_, _20943_);
  nor (_20946_, _20945_, _20916_);
  or (_20947_, _20564_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_20948_, _20564_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_20949_, _20948_, _20947_);
  or (_20950_, _20949_, _20550_);
  nand (_20951_, _20949_, _20550_);
  and (_20952_, _20951_, _20950_);
  not (_20953_, _20952_);
  nand (_20954_, _20953_, _20910_);
  or (_20955_, _20953_, _20910_);
  and (_20956_, _20955_, _20954_);
  and (_20957_, _20908_, _20572_);
  nor (_20958_, _20957_, _20909_);
  nor (_20959_, _20958_, _22853_);
  and (_20960_, _20958_, _22853_);
  nor (_20961_, _20904_, _20902_);
  nor (_20962_, _20961_, _20905_);
  nor (_20963_, _20962_, _22824_);
  nor (_20964_, _20587_, _20588_);
  nor (_20965_, _20964_, _20900_);
  and (_20966_, _20964_, _20900_);
  or (_20967_, _20966_, _20965_);
  and (_20968_, _20967_, _23972_);
  nor (_20969_, _20967_, _23972_);
  and (_20970_, _20898_, _20633_);
  nor (_20971_, _20970_, _20899_);
  nor (_20972_, _20971_, _26118_);
  and (_20973_, _20971_, _26118_);
  and (_20974_, _20896_, _20678_);
  nor (_20975_, _20974_, _20897_);
  and (_20976_, _20975_, _26122_);
  nor (_20977_, _20975_, _26122_);
  and (_20978_, _20894_, _20891_);
  nor (_20979_, _20978_, _20895_);
  and (_20980_, _20979_, _22807_);
  nor (_20981_, _20979_, _22807_);
  and (_20982_, _20889_, _20762_);
  nor (_20983_, _20982_, _20890_);
  nor (_20984_, _20983_, _26129_);
  and (_20985_, _20983_, _26129_);
  and (_20986_, _20887_, _20884_);
  nor (_20987_, _20986_, _20888_);
  nor (_20988_, _20987_, _26133_);
  nor (_20989_, _20882_, _20880_);
  nor (_20990_, _20989_, _20883_);
  and (_20991_, _20990_, _26137_);
  and (_20992_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20993_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_20994_, _20993_, _20992_);
  and (_20995_, _20994_, _20879_);
  nor (_20996_, _20994_, _20879_);
  or (_20997_, _20996_, _20995_);
  nor (_20998_, _20990_, _26137_);
  or (_20999_, _20998_, _20997_);
  or (_21000_, _20999_, _20991_);
  and (_21001_, _20987_, _26133_);
  or (_21002_, _21001_, _21000_);
  or (_21003_, _21002_, _20988_);
  or (_21004_, _21003_, _20985_);
  or (_21005_, _21004_, _20984_);
  or (_21006_, _21005_, _20981_);
  or (_21007_, _21006_, _20980_);
  or (_21008_, _21007_, _20977_);
  or (_21009_, _21008_, _20976_);
  or (_21010_, _21009_, _20973_);
  or (_21011_, _21010_, _20972_);
  or (_21012_, _21011_, _20969_);
  or (_21013_, _21012_, _20968_);
  or (_21014_, _21013_, _20963_);
  nor (_21015_, _20905_, _20579_);
  and (_21016_, _20581_, _24590_);
  nor (_21017_, _20581_, _24590_);
  nor (_21018_, _21017_, _21016_);
  not (_21019_, _21018_);
  nor (_21020_, _21019_, _21015_);
  and (_21021_, _20962_, _22824_);
  and (_21022_, _21019_, _21015_);
  or (_21023_, _21022_, _21021_);
  or (_21024_, _21023_, _21020_);
  or (_21025_, _21024_, _21014_);
  or (_21026_, _21025_, _20960_);
  or (_21027_, _21026_, _20959_);
  or (_21028_, _21027_, _20956_);
  or (_21029_, _21028_, _20946_);
  nor (_21030_, _20914_, _20912_);
  nor (_21031_, _21030_, _20915_);
  nor (_21032_, _21031_, _22776_);
  and (_21033_, _20945_, _20916_);
  and (_21034_, _21031_, _22776_);
  or (_21035_, _21034_, _21033_);
  or (_21036_, _21035_, _21032_);
  or (_21037_, _21036_, _21029_);
  or (_21038_, _21037_, _20938_);
  or (_21039_, _21038_, _20937_);
  or (_21040_, _21039_, _20924_);
  or (_21041_, \oc8051_symbolic_cxrom1.regvalid [13], _26129_);
  or (_21042_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21043_, _21042_, _21041_);
  and (_21044_, _26133_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21045_, _21044_, _21043_);
  or (_21046_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21047_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_21048_, \oc8051_symbolic_cxrom1.regvalid [1], _26129_);
  and (_21049_, _21048_, _21047_);
  and (_21050_, _21049_, _21046_);
  or (_21051_, _21050_, _21045_);
  nor (_21052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21053_, _21052_, _26133_);
  nor (_21054_, _21053_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21055_, _21053_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21056_, _21055_, _21054_);
  and (_21057_, _21056_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_21058_, _21052_, _26133_);
  nor (_21059_, _21058_, _21053_);
  nand (_21060_, \oc8051_symbolic_cxrom1.regvalid [7], _26129_);
  nand (_21061_, _21060_, _21059_);
  or (_21062_, _21061_, _21057_);
  and (_21063_, _21062_, _26137_);
  nand (_21064_, _21056_, _06111_);
  or (_21065_, _21056_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_21066_, _21065_, _21064_);
  or (_21067_, _21059_, _21066_);
  and (_21068_, _21067_, _21063_);
  or (_21069_, _21068_, _21051_);
  and (_21070_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21071_, \oc8051_symbolic_cxrom1.regvalid [0], _26129_);
  or (_21072_, _21071_, _21070_);
  and (_21073_, _21072_, _26133_);
  and (_21074_, \oc8051_symbolic_cxrom1.regvalid [4], _26129_);
  and (_21075_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21076_, _21075_, _21074_);
  and (_21077_, _21076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21078_, _21077_, _21073_);
  and (_21079_, _21078_, _26137_);
  and (_21080_, _21047_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21081_, _21080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21082_, _21080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21083_, _21082_, _21081_);
  or (_21084_, _21083_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_21085_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21086_, _21085_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_21087_, _21086_, _21080_);
  and (_21088_, _21087_, _21041_);
  and (_21089_, _21088_, _21084_);
  or (_21090_, _21083_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_21091_, _21087_);
  nand (_21092_, _21083_, _05493_);
  and (_21093_, _21092_, _21091_);
  and (_21094_, _21093_, _21090_);
  or (_21095_, _21094_, _21089_);
  and (_21096_, _21095_, _21079_);
  or (_21097_, _21083_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_21098_, \oc8051_symbolic_cxrom1.regvalid [15], _26129_);
  and (_21099_, _21098_, _21087_);
  and (_21100_, _21099_, _21097_);
  or (_21101_, _21083_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_21102_, _21083_, _06111_);
  and (_21103_, _21102_, _21091_);
  and (_21104_, _21103_, _21101_);
  or (_21105_, _21104_, _21100_);
  and (_21106_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21107_, \oc8051_symbolic_cxrom1.regvalid [6], _26129_);
  or (_21108_, _21107_, _26133_);
  or (_21109_, _21108_, _21106_);
  or (_21110_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21111_, \oc8051_symbolic_cxrom1.regvalid [10], _26129_);
  and (_21112_, _21111_, _21110_);
  or (_21113_, _21112_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21114_, _21113_, _21109_);
  and (_21115_, _21114_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21116_, _21076_, _21044_);
  or (_21117_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21118_, \oc8051_symbolic_cxrom1.regvalid [0], _26129_);
  and (_21119_, _21118_, _21047_);
  and (_21120_, _21119_, _21117_);
  or (_21121_, _21120_, _21116_);
  and (_21122_, _21121_, _21115_);
  and (_21123_, _21122_, _21105_);
  or (_21124_, _21123_, _21096_);
  or (_21125_, _21121_, _21114_);
  and (_21126_, _21125_, _26141_);
  and (_21127_, _21126_, _21124_);
  and (_21128_, _21127_, _21069_);
  or (_21129_, \oc8051_symbolic_cxrom1.regvalid [2], _26137_);
  or (_21130_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21131_, _21130_, _21129_);
  or (_21132_, _21131_, _21056_);
  or (_21133_, \oc8051_symbolic_cxrom1.regvalid [10], _26137_);
  or (_21134_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_21135_, _21134_, _21133_);
  and (_21136_, _21135_, _21056_);
  nor (_21137_, _21136_, _21059_);
  and (_21138_, _21137_, _21132_);
  and (_21139_, _21056_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_21140_, _21074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_21141_, _21140_, _21139_);
  and (_21142_, _21056_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_21143_, _21107_, _26137_);
  or (_21144_, _21143_, _21142_);
  and (_21145_, _21144_, _21059_);
  and (_21146_, _21145_, _21141_);
  or (_21147_, _21146_, _21138_);
  or (_21148_, _21083_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_21149_, \oc8051_symbolic_cxrom1.regvalid [14], _26129_);
  and (_21150_, _21149_, _21148_);
  or (_21151_, _21150_, _21091_);
  nand (_21152_, _21083_, _06073_);
  or (_21153_, _21083_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_21154_, _21153_, _21152_);
  or (_21155_, _21154_, _21087_);
  and (_21156_, _21155_, _21151_);
  or (_21157_, _21156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_21158_, _21083_, _20488_);
  and (_21159_, _21083_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_21160_, _21159_, _21158_);
  and (_21161_, _21160_, _21091_);
  or (_21162_, _21083_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_21163_, \oc8051_symbolic_cxrom1.regvalid [12], _26129_);
  and (_21164_, _21163_, _21087_);
  and (_21165_, _21164_, _21162_);
  or (_21166_, _21165_, _26137_);
  or (_21167_, _21166_, _21161_);
  or (_21168_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21169_, _21168_, _21098_);
  or (_21170_, _21169_, _26133_);
  or (_21171_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21172_, \oc8051_symbolic_cxrom1.regvalid [11], _26129_);
  and (_21173_, _21172_, _21171_);
  or (_21174_, _21173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21175_, _21174_, _21170_);
  and (_21176_, _21175_, _21085_);
  and (_21177_, _26137_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_21178_, _21043_, _26133_);
  or (_21179_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21180_, \oc8051_symbolic_cxrom1.regvalid [9], _26129_);
  and (_21181_, _21180_, _21179_);
  or (_21182_, _21181_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21183_, _21182_, _21178_);
  and (_21184_, _21183_, _21177_);
  or (_21185_, _21184_, _21176_);
  and (_21186_, _21175_, _26137_);
  or (_21187_, _21186_, _21051_);
  and (_21188_, _21187_, _21185_);
  and (_21189_, _21188_, _21167_);
  and (_21190_, _21189_, _21157_);
  and (_21191_, _21190_, _21147_);
  or (_21192_, _21191_, _21128_);
  nor (_21193_, _20447_, _22798_);
  and (_21194_, _20449_, _22794_);
  nor (_21195_, _21194_, _21193_);
  not (_21196_, _21195_);
  and (_21197_, _21193_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21198_, _21193_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21199_, _21198_, _21197_);
  and (_21200_, _21199_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_21201_, _21199_, _05479_);
  or (_21202_, _21201_, _21200_);
  and (_21203_, _21202_, _21196_);
  nand (_21204_, _21199_, _05487_);
  nor (_21205_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21206_, _21205_, _21196_);
  and (_21207_, _21206_, _21204_);
  or (_21208_, _21207_, _21203_);
  and (_21209_, _21208_, _20447_);
  and (_21210_, _21199_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_21211_, _21199_, _20488_);
  or (_21212_, _21211_, _21210_);
  and (_21213_, _21212_, _21196_);
  or (_21214_, _21199_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_21215_, \oc8051_symbolic_cxrom1.regvalid [12], _22802_);
  nor (_21216_, _21215_, _21196_);
  and (_21217_, _21216_, _21214_);
  or (_21218_, _21217_, _21213_);
  and (_21219_, _21218_, _20499_);
  or (_21220_, _21219_, _21209_);
  and (_21221_, _21199_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_21222_, _21199_, _05519_);
  or (_21223_, _21222_, _21221_);
  and (_21224_, _21223_, _21196_);
  nand (_21225_, _21199_, _05504_);
  nor (_21226_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21227_, _21226_, _21196_);
  and (_21228_, _21227_, _21225_);
  or (_21229_, _21228_, _21224_);
  and (_21230_, _21229_, _20486_);
  and (_21231_, _21199_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_21232_, _21199_, _05885_);
  or (_21233_, _21232_, _21231_);
  and (_21234_, _21233_, _21196_);
  nand (_21235_, _21199_, _05456_);
  nor (_21236_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21237_, _21236_, _21196_);
  and (_21238_, _21237_, _21235_);
  or (_21239_, _21238_, _21234_);
  and (_21240_, _21239_, _20472_);
  or (_21241_, _21240_, _21230_);
  or (_21242_, _21241_, _21220_);
  and (_21243_, _05487_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21244_, _21243_);
  nor (_21245_, _21205_, _22798_);
  and (_21246_, _21245_, _21244_);
  and (_21247_, _06111_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21248_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21249_, _21248_, _21247_);
  and (_21250_, _21249_, _22798_);
  nor (_21251_, _21250_, _21246_);
  nor (_21252_, _21251_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21253_, _05456_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21254_, _21253_, _21236_);
  and (_21255_, _21254_, _20450_);
  or (_21256_, _21255_, _21252_);
  and (_21257_, _21256_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21258_, _05504_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21259_, _21258_);
  nor (_21260_, _21226_, _22798_);
  and (_21261_, _21260_, _21259_);
  and (_21262_, _06073_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21263_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21264_, _21263_, _21262_);
  and (_21265_, _21264_, _22798_);
  nor (_21266_, _21265_, _21261_);
  nor (_21267_, _21266_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21268_, _20488_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21269_, _21268_);
  not (_21270_, _20432_);
  nor (_21271_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21272_, _21271_, _21270_);
  and (_21273_, _21272_, _21269_);
  nor (_21274_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21275_, _21274_, _21215_);
  and (_21276_, _21275_, _20450_);
  or (_21277_, _21276_, _21273_);
  or (_21278_, _21277_, _21267_);
  and (_21279_, _21278_, _22789_);
  and (_21280_, _05885_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21281_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21282_, _21281_, _22798_);
  nor (_21283_, _21282_, _21280_);
  and (_21284_, _21283_, _20486_);
  or (_21285_, _21284_, _21279_);
  or (_21286_, _21285_, _21257_);
  nor (_21287_, _21266_, _22794_);
  nor (_21288_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21289_, _05526_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21290_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21291_, _21290_, _21289_);
  and (_21292_, _21291_, _21288_);
  and (_21293_, _21275_, _20451_);
  or (_21294_, _21293_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_21295_, _21294_, _21292_);
  nor (_21296_, _21295_, _21287_);
  nor (_21297_, _21251_, _22794_);
  nor (_21298_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_21299_, _05493_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21300_, _21299_, _21298_);
  and (_21301_, _21300_, _21288_);
  and (_21302_, _21254_, _20451_);
  or (_21303_, _21302_, _22789_);
  or (_21304_, _21303_, _21301_);
  nor (_21305_, _21304_, _21297_);
  nor (_21306_, _21305_, _21296_);
  not (_21307_, _22770_);
  nor (_21308_, _21307_, first_instr);
  and (_21309_, _21308_, _21306_);
  and (_21310_, _21309_, _21286_);
  nand (_21311_, _21310_, _21242_);
  nor (_21312_, _21311_, _20512_);
  and (_21313_, _21312_, _21192_);
  nor (_21314_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21315_, _07000_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21316_, _21315_, _21314_);
  and (_21317_, _21316_, _20451_);
  nor (_21318_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21319_, _06502_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21320_, _21319_, _21318_);
  and (_21321_, _21320_, _21288_);
  nor (_21322_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21323_, _07267_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21324_, _21323_, _21322_);
  and (_21325_, _21324_, _20432_);
  or (_21326_, _21325_, _21321_);
  nor (_21327_, _21326_, _21317_);
  nor (_21328_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21329_, _06751_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21330_, _21329_, _21328_);
  and (_21331_, _21330_, _20450_);
  nor (_21332_, _21331_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_21333_, _21332_, _21327_);
  nor (_21334_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21335_, _08334_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21336_, _21335_, _21334_);
  and (_21337_, _21336_, _20432_);
  nor (_21338_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21339_, _08053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21340_, _21339_, _21338_);
  and (_21341_, _21340_, _20451_);
  nor (_21342_, _21341_, _21337_);
  nor (_21343_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21344_, _07761_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21345_, _21344_, _21343_);
  and (_21346_, _21345_, _20450_);
  nor (_21347_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21348_, _07551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21349_, _21348_, _21347_);
  and (_21350_, _21349_, _21288_);
  nor (_21351_, _21350_, _21346_);
  and (_21352_, _21351_, _21342_);
  and (_21353_, _21352_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21354_, _21353_, _21333_);
  and (_21355_, _21354_, _21306_);
  nor (_21356_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21357_, _06731_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21358_, _21357_, _21356_);
  and (_21359_, _21358_, _20450_);
  nor (_21360_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21361_, _06979_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21362_, _21361_, _21360_);
  and (_21363_, _21362_, _20451_);
  nor (_21364_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21365_, _06478_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21366_, _21365_, _21364_);
  and (_21367_, _21366_, _21288_);
  nor (_21368_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21369_, _07248_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21370_, _21369_, _21368_);
  and (_21371_, _21370_, _20432_);
  or (_21372_, _21371_, _21367_);
  or (_21373_, _21372_, _21363_);
  or (_21374_, _21373_, _21359_);
  and (_21375_, _21374_, _22802_);
  nor (_21376_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21377_, _07743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21378_, _21377_, _21376_);
  and (_21379_, _21378_, _20450_);
  nor (_21380_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21381_, _08043_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21382_, _21381_, _21380_);
  and (_21383_, _21382_, _20451_);
  nor (_21384_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21385_, _07532_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21386_, _21385_, _21384_);
  and (_21387_, _21386_, _21288_);
  nor (_21388_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21389_, _08320_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21390_, _21389_, _21388_);
  and (_21391_, _21390_, _20432_);
  or (_21392_, _21391_, _21387_);
  or (_21393_, _21392_, _21383_);
  or (_21394_, _21393_, _21379_);
  and (_21395_, _21394_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21396_, _21395_, _21375_);
  and (_21397_, _21396_, _21306_);
  nor (_21398_, _21397_, _21355_);
  nor (_21399_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21400_, _07061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21401_, _21400_, _21399_);
  and (_21402_, _21401_, _20451_);
  nor (_21403_, _21402_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21404_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21405_, _06804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21406_, _21405_, _21404_);
  and (_21407_, _21406_, _20450_);
  nor (_21408_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21409_, _06568_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21410_, _21409_, _21408_);
  and (_21411_, _21410_, _21288_);
  nor (_21412_, _21411_, _21407_);
  nor (_21413_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21414_, _07341_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21415_, _21414_, _21413_);
  and (_21416_, _21415_, _20432_);
  not (_21417_, _21416_);
  and (_21418_, _21417_, _21412_);
  and (_21419_, _21418_, _21403_);
  nor (_21420_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21421_, _08110_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21422_, _21421_, _21420_);
  and (_21423_, _21422_, _20451_);
  nor (_21424_, _21423_, _22802_);
  nor (_21425_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21426_, _07601_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21427_, _21426_, _21425_);
  and (_21428_, _21427_, _21288_);
  not (_21429_, _21428_);
  nor (_21430_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21431_, _07814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21432_, _21431_, _21430_);
  and (_21433_, _21432_, _20450_);
  nor (_21434_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21435_, _08391_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21436_, _21435_, _21434_);
  and (_21437_, _21436_, _20432_);
  nor (_21438_, _21437_, _21433_);
  and (_21439_, _21438_, _21429_);
  and (_21440_, _21439_, _21424_);
  nor (_21441_, _21440_, _21419_);
  and (_21442_, _21441_, _21306_);
  nor (_21443_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21444_, _06792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21445_, _21444_, _21443_);
  and (_21446_, _21445_, _20450_);
  nor (_21447_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21448_, _07047_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21449_, _21448_, _21447_);
  and (_21450_, _21449_, _20451_);
  nor (_21451_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21452_, _06551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21453_, _21452_, _21451_);
  and (_21454_, _21453_, _21288_);
  nor (_21455_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21456_, _07321_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21457_, _21456_, _21455_);
  and (_21458_, _21457_, _20432_);
  or (_21459_, _21458_, _21454_);
  or (_21460_, _21459_, _21450_);
  or (_21461_, _21460_, _21446_);
  and (_21462_, _21461_, _22802_);
  nor (_21463_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21464_, _07800_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21465_, _21464_, _21463_);
  and (_21466_, _21465_, _20450_);
  nor (_21467_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21468_, _08098_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21469_, _21468_, _21467_);
  and (_21470_, _21469_, _20451_);
  nor (_21471_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21472_, _07589_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21473_, _21472_, _21471_);
  and (_21474_, _21473_, _21288_);
  nor (_21475_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21476_, _08379_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21477_, _21476_, _21475_);
  and (_21478_, _21477_, _20432_);
  or (_21479_, _21478_, _21474_);
  or (_21480_, _21479_, _21470_);
  or (_21481_, _21480_, _21466_);
  and (_21482_, _21481_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21483_, _21482_, _21462_);
  and (_21484_, _21483_, _21306_);
  nor (_21485_, _21484_, _21442_);
  and (_21486_, _21485_, _21398_);
  nor (_21487_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21488_, _06766_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21489_, _21488_, _21487_);
  and (_21490_, _21489_, _20450_);
  nor (_21491_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21492_, _07016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21493_, _21492_, _21491_);
  and (_21494_, _21493_, _20451_);
  nor (_21495_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21496_, _06516_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21497_, _21496_, _21495_);
  and (_21498_, _21497_, _21288_);
  nor (_21499_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21500_, _07287_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21501_, _21500_, _21499_);
  and (_21502_, _21501_, _20432_);
  or (_21503_, _21502_, _21498_);
  or (_21504_, _21503_, _21494_);
  or (_21505_, _21504_, _21490_);
  and (_21506_, _21505_, _22802_);
  nor (_21507_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21508_, _07772_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21509_, _21508_, _21507_);
  and (_21510_, _21509_, _20450_);
  nor (_21511_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21512_, _08072_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21513_, _21512_, _21511_);
  and (_21514_, _21513_, _20451_);
  nor (_21515_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21516_, _07564_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21517_, _21516_, _21515_);
  and (_21518_, _21517_, _21288_);
  nor (_21519_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21520_, _08349_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21521_, _21520_, _21519_);
  and (_21522_, _21521_, _20432_);
  or (_21523_, _21522_, _21518_);
  or (_21524_, _21523_, _21514_);
  or (_21525_, _21524_, _21510_);
  and (_21526_, _21525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21527_, _21526_, _21506_);
  and (_21528_, _21527_, _21306_);
  nor (_21529_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21530_, _06779_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21531_, _21530_, _21529_);
  and (_21532_, _21531_, _20450_);
  nor (_21533_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21534_, _07033_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21535_, _21534_, _21533_);
  and (_21536_, _21535_, _20451_);
  nor (_21537_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21538_, _07303_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21539_, _21538_, _21537_);
  and (_21540_, _21539_, _20432_);
  nor (_21541_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21542_, _06536_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21543_, _21542_, _21541_);
  and (_21544_, _21543_, _21288_);
  or (_21545_, _21544_, _21540_);
  or (_21546_, _21545_, _21536_);
  or (_21547_, _21546_, _21532_);
  and (_21548_, _21547_, _22802_);
  nor (_21549_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21550_, _07786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21551_, _21550_, _21549_);
  and (_21552_, _21551_, _20450_);
  nor (_21553_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21554_, _08085_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21555_, _21554_, _21553_);
  and (_21556_, _21555_, _20451_);
  nor (_21557_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21558_, _08363_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21559_, _21558_, _21557_);
  and (_21560_, _21559_, _20432_);
  nor (_21561_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21562_, _07576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21563_, _21562_, _21561_);
  and (_21564_, _21563_, _21288_);
  or (_21565_, _21564_, _21560_);
  or (_21566_, _21565_, _21556_);
  or (_21567_, _21566_, _21552_);
  and (_21568_, _21567_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21569_, _21568_, _21548_);
  and (_21570_, _21569_, _21306_);
  nor (_21571_, _21570_, _21528_);
  nor (_21572_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21573_, _05539_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21574_, _21573_, _21572_);
  and (_21575_, _21574_, _21288_);
  nor (_21576_, _21575_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21577_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21578_, _05551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21579_, _21578_, _21577_);
  and (_21580_, _21579_, _20451_);
  not (_21581_, _21580_);
  nor (_21582_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21583_, _05556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21585_, _21583_, _21582_);
  and (_21586_, _21585_, _20450_);
  nor (_21587_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21588_, _05546_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21589_, _21588_, _21587_);
  and (_21590_, _21589_, _20432_);
  nor (_21591_, _21590_, _21586_);
  and (_21592_, _21591_, _21581_);
  and (_21593_, _21592_, _21576_);
  nor (_21594_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21595_, _05564_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21596_, _21595_, _21594_);
  and (_21597_, _21596_, _21288_);
  nor (_21598_, _21597_, _22802_);
  nor (_21599_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21600_, _05570_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21601_, _21600_, _21599_);
  and (_21602_, _21601_, _20451_);
  not (_21603_, _21602_);
  nor (_21604_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21605_, _05584_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21606_, _21605_, _21604_);
  and (_21607_, _21606_, _20450_);
  nor (_21608_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21609_, _05576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21610_, _21609_, _21608_);
  and (_21611_, _21610_, _20432_);
  nor (_21612_, _21611_, _21607_);
  and (_21613_, _21612_, _21603_);
  and (_21614_, _21613_, _21598_);
  nor (_21615_, _21614_, _21593_);
  and (_21616_, _21615_, _21306_);
  not (_21617_, _21616_);
  nor (_21618_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21619_, _06817_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21620_, _21619_, _21618_);
  and (_21621_, _21620_, _20450_);
  nor (_21622_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21623_, _07074_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21624_, _21623_, _21622_);
  and (_21625_, _21624_, _20451_);
  nor (_21626_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21627_, _06582_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21628_, _21627_, _21626_);
  and (_21629_, _21628_, _21288_);
  nor (_21630_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21631_, _07361_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21632_, _21631_, _21630_);
  and (_21633_, _21632_, _20432_);
  or (_21634_, _21633_, _21629_);
  or (_21635_, _21634_, _21625_);
  or (_21636_, _21635_, _21621_);
  and (_21637_, _21636_, _22802_);
  nor (_21638_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21639_, _07829_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21640_, _21639_, _21638_);
  and (_21641_, _21640_, _20450_);
  nor (_21642_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21643_, _08121_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21644_, _21643_, _21642_);
  and (_21645_, _21644_, _20451_);
  nor (_21646_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21647_, _07614_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21648_, _21647_, _21646_);
  and (_21649_, _21648_, _21288_);
  nor (_21650_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21651_, _08406_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21652_, _21651_, _21650_);
  and (_21653_, _21652_, _20432_);
  or (_21654_, _21653_, _21649_);
  or (_21655_, _21654_, _21645_);
  or (_21656_, _21655_, _21641_);
  and (_21657_, _21656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21658_, _21657_, _21637_);
  nor (_21659_, _21658_, _21617_);
  and (_21660_, _21659_, _21571_);
  and (_21661_, _21660_, _21486_);
  and (_21662_, _21661_, _21313_);
  and (_21663_, _21662_, _21040_);
  and (_21664_, _21658_, _21306_);
  not (_21665_, _21397_);
  not (_21666_, _21570_);
  not (_21667_, _21355_);
  and (_21668_, _21528_, _21667_);
  and (_21669_, _21668_, _21666_);
  and (_21670_, _21669_, _21665_);
  and (_21671_, _21527_, _21355_);
  and (_21672_, _21483_, _21442_);
  and (_21673_, _21672_, _21671_);
  and (_21674_, _21571_, _21665_);
  and (_21675_, _21674_, _21355_);
  and (_21676_, _21569_, _21442_);
  and (_21677_, _21676_, _21483_);
  or (_21678_, _21677_, _21675_);
  or (_21679_, _21678_, _21673_);
  or (_21680_, _21679_, _21670_);
  and (_21681_, _21680_, _21664_);
  not (_21682_, _21442_);
  nor (_21683_, _21658_, _21682_);
  and (_21684_, _21683_, _21669_);
  and (_21685_, _21669_, _21397_);
  and (_21686_, _21685_, _21682_);
  or (_21687_, _21686_, _21684_);
  or (_21688_, _21687_, _21681_);
  and (_21689_, _21688_, _21617_);
  not (_21690_, _21484_);
  and (_21691_, _21685_, _21690_);
  not (_21692_, _21441_);
  and (_21693_, _21616_, _21692_);
  and (_21694_, _21693_, _21674_);
  or (_21695_, _21694_, _21691_);
  and (_21696_, _21695_, _21664_);
  and (_21697_, _21675_, _21682_);
  and (_21698_, _21664_, _21441_);
  and (_21699_, _21698_, _21685_);
  or (_21700_, _21699_, _21697_);
  and (_21701_, _21700_, _21616_);
  and (_21702_, _21659_, _21692_);
  and (_21703_, _21702_, _21484_);
  and (_21704_, _21703_, _21669_);
  nor (_21705_, _21682_, _21396_);
  and (_21706_, _21705_, _21571_);
  and (_21707_, _21671_, _21690_);
  and (_21708_, _21570_, _21690_);
  or (_21709_, _21708_, _21707_);
  or (_21710_, _21709_, _21706_);
  and (_21711_, _21710_, _21659_);
  or (_21712_, _21711_, _21704_);
  or (_21713_, _21712_, _21701_);
  or (_21714_, _21713_, _21696_);
  or (_21715_, _21714_, _21689_);
  nor (_21716_, _20561_, _22776_);
  and (_21717_, _20561_, _22776_);
  or (_21718_, _21717_, _21716_);
  nor (_21719_, _20446_, _22784_);
  or (_21720_, _21719_, _21718_);
  nand (_21721_, _20446_, _22784_);
  nand (_21722_, _21721_, _20933_);
  or (_21723_, _21722_, _20942_);
  or (_21724_, _21723_, _21720_);
  nor (_21725_, _20591_, _26118_);
  nor (_21726_, _20452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21727_, _20452_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21728_, _21727_, _21726_);
  nor (_21729_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_21730_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_21731_, _21730_, _21729_);
  not (_21732_, _21731_);
  and (_21733_, _21732_, _20433_);
  or (_21734_, _21733_, _21728_);
  and (_21735_, _20458_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21736_, _20458_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21737_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21738_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21739_, _21738_, _21737_);
  nand (_21740_, _21739_, _20994_);
  nor (_21741_, _21732_, _20433_);
  or (_21742_, _21741_, _21740_);
  or (_21743_, _21742_, _21736_);
  or (_21744_, _21743_, _21735_);
  or (_21745_, _21744_, _21734_);
  and (_21746_, _20591_, _26118_);
  or (_21747_, _21746_, _21745_);
  or (_21748_, _21747_, _21725_);
  or (_21749_, _20578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_21750_, _20578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_21751_, _21750_, _21749_);
  nor (_21752_, _20636_, _26122_);
  and (_21753_, _20636_, _26122_);
  or (_21754_, _21753_, _21752_);
  nor (_21755_, _20585_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_21756_, _20585_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_21757_, _21756_, _21755_);
  or (_21758_, _21757_, _21754_);
  or (_21759_, _21758_, _21751_);
  or (_21760_, _21759_, _21748_);
  nor (_21761_, _20568_, _22853_);
  and (_21762_, _20568_, _22853_);
  or (_21763_, _21762_, _21761_);
  nor (_21764_, _20575_, _24590_);
  and (_21765_, _20575_, _24590_);
  or (_21766_, _21765_, _21764_);
  or (_21767_, _21766_, _20949_);
  or (_21768_, _21767_, _21763_);
  or (_21769_, _21768_, _21760_);
  or (_21770_, _21769_, _21724_);
  and (_21771_, _21770_, _21715_);
  and (_21772_, _21684_, _21690_);
  and (_21773_, _21528_, _21665_);
  and (_21774_, _21773_, _21666_);
  or (_21775_, _21705_, _21676_);
  or (_21776_, _21775_, _21774_);
  and (_21777_, _21776_, _21664_);
  or (_21778_, _21777_, _21772_);
  and (_21779_, _21778_, _21616_);
  not (_21780_, _21664_);
  and (_21781_, _21396_, _21355_);
  and (_21782_, _21781_, _21571_);
  and (_21783_, _21670_, _21485_);
  or (_21784_, _21783_, _21782_);
  and (_21785_, _21784_, _21780_);
  nor (_21786_, _21617_, _21569_);
  and (_21787_, _21786_, _21781_);
  or (_21788_, _21787_, _21707_);
  and (_21789_, _21788_, _21664_);
  and (_21790_, _21780_, _21570_);
  not (_21791_, _21615_);
  and (_21792_, _21484_, _21692_);
  or (_21793_, _21792_, _21791_);
  and (_21794_, _21793_, _21790_);
  nor (_21795_, _21615_, _21441_);
  and (_21796_, _21795_, _21570_);
  and (_21797_, _21708_, _21664_);
  or (_21798_, _21797_, _21796_);
  or (_21799_, _21798_, _21794_);
  or (_21800_, _21799_, _21789_);
  nor (_21801_, _21664_, _21616_);
  and (_21802_, _21773_, _21682_);
  or (_21803_, _21802_, _21486_);
  and (_21804_, _21803_, _21801_);
  and (_21805_, _21792_, _21666_);
  or (_21806_, _21805_, _21801_);
  and (_21807_, _21806_, _21671_);
  or (_21808_, _21807_, _21804_);
  or (_21809_, _21808_, _21800_);
  or (_21810_, _21809_, _21785_);
  or (_21811_, _21810_, _21779_);
  and (_21812_, _20444_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21813_, _20443_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21814_, _21813_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21815_, _21814_, _21812_);
  and (_21816_, _21815_, _22784_);
  nor (_21817_, _21815_, _22784_);
  or (_21818_, _21817_, _21816_);
  and (_21819_, _20441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21820_, _21819_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_21821_, _21820_, _22844_);
  and (_21822_, _21820_, _22844_);
  nor (_21823_, _21822_, _21821_);
  and (_21824_, _21823_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_21825_, _21823_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_21826_, _21825_, _21824_);
  or (_21827_, _21826_, _21818_);
  and (_21828_, _20433_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21829_, _21828_, _20436_);
  and (_21830_, _21829_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_21831_, _21830_, _22828_);
  nor (_21832_, _21830_, _22828_);
  nor (_21833_, _21832_, _21831_);
  and (_21834_, _21833_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_21835_, _20564_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_21836_, _22837_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21837_, _21836_, _21835_);
  and (_21838_, _21837_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_21839_, _21812_, _20930_);
  or (_21840_, _21839_, _21838_);
  or (_21841_, _21840_, _21834_);
  nor (_21842_, _21833_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_21843_, _20582_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21844_, _21843_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_21845_, _21844_, _21829_);
  nor (_21846_, _21845_, _23972_);
  and (_21847_, _21845_, _23972_);
  or (_21848_, _21739_, _22789_);
  nand (_21849_, _21739_, _22789_);
  and (_21850_, _21849_, _21848_);
  nor (_21851_, _21828_, _21732_);
  and (_21852_, _21828_, _21732_);
  or (_21853_, _21852_, _20994_);
  nor (_21854_, _21853_, _21851_);
  nand (_21855_, _21854_, _21850_);
  or (_21856_, _21855_, _21847_);
  or (_21857_, _21856_, _21846_);
  nor (_21858_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_21859_, _21858_, _21843_);
  nor (_21860_, _21859_, _20590_);
  nor (_21861_, _21860_, _26118_);
  and (_21862_, _20461_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21863_, _20461_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21864_, _21863_, _21862_);
  nor (_21865_, _20454_, _26133_);
  and (_21866_, _20454_, _26133_);
  or (_21867_, _21866_, _21865_);
  or (_21868_, _21867_, _21864_);
  or (_21869_, _21868_, _21861_);
  or (_21870_, _21869_, _21857_);
  or (_21871_, _22811_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_21872_, _20636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21873_, _21872_, _21871_);
  and (_21874_, _21873_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_21875_, _21873_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_21876_, _21875_, _21874_);
  or (_21877_, _21876_, _21870_);
  or (_21878_, _21877_, _21842_);
  nor (_21879_, _21837_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_21880_, _21812_, _20930_);
  or (_21881_, _21880_, _21879_);
  or (_21882_, _21881_, _21878_);
  nor (_21883_, _21819_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_21884_, _21883_, _21820_);
  nand (_21885_, _21884_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_21886_, _21884_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_21887_, _21886_, _21885_);
  and (_21888_, _21829_, _20438_);
  and (_21889_, _21888_, _22833_);
  nor (_21890_, _21888_, _22833_);
  or (_21891_, _21890_, _21889_);
  and (_21892_, _21891_, _22853_);
  nor (_21893_, _21891_, _22853_);
  nor (_21894_, _21829_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_21896_, _21894_, _21830_);
  nor (_21897_, _21896_, _22824_);
  and (_21898_, _21896_, _22824_);
  or (_21899_, _21898_, _21897_);
  and (_21900_, _21860_, _26118_);
  or (_21901_, _21900_, _21899_);
  or (_21902_, _21901_, _21893_);
  or (_21903_, _21902_, _21892_);
  or (_21904_, _21903_, _21887_);
  or (_21905_, _21904_, _21882_);
  or (_21906_, _21905_, _21841_);
  or (_21907_, _21906_, _21827_);
  and (_21908_, _21907_, _21811_);
  and (_21909_, _21702_, _21691_);
  and (_21910_, _21571_, _21398_);
  and (_21911_, _21910_, _21703_);
  or (_21912_, _21911_, _21909_);
  and (_21913_, _21699_, _21484_);
  nor (_21914_, _21672_, _21780_);
  and (_21915_, _21914_, _21782_);
  or (_21916_, _21915_, _21913_);
  and (_21917_, _21916_, _21617_);
  or (_21918_, _21917_, _21912_);
  and (_21919_, _21197_, _20436_);
  and (_21920_, _21919_, _20438_);
  and (_21921_, _21920_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_21922_, _21921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_21923_, _21922_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_21924_, _21923_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_21925_, _21923_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_21927_, _21925_, _21924_);
  nor (_21928_, _21927_, _22780_);
  and (_21929_, _21924_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21930_, _21929_, _20930_);
  and (_21931_, _21929_, _20930_);
  or (_21932_, _21931_, _21930_);
  or (_21933_, _21932_, _21928_);
  nor (_21934_, _21924_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21935_, _21934_, _21929_);
  nor (_21936_, _21935_, _22784_);
  and (_21937_, _21935_, _22784_);
  or (_21938_, _21937_, _21936_);
  nor (_21939_, _21922_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_21940_, _21939_, _21923_);
  and (_21941_, _21940_, _22776_);
  nor (_21942_, _21940_, _22776_);
  and (_21943_, _21919_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_21944_, _21919_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_21945_, _21944_, _21943_);
  nor (_21946_, _21945_, _22824_);
  and (_21948_, _21945_, _22824_);
  or (_21949_, _21948_, _21946_);
  and (_21950_, _21197_, _20434_);
  and (_21951_, _21197_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_21952_, _21951_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_21953_, _21952_, _21950_);
  and (_21954_, _21953_, _26122_);
  nor (_21955_, _21953_, _26122_);
  or (_21956_, _21955_, _21954_);
  or (_21957_, _21956_, _21949_);
  and (_21958_, _21197_, _20435_);
  nor (_21959_, _21950_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_21960_, _21959_, _21958_);
  and (_21961_, _21960_, _26118_);
  or (_21962_, _21731_, _21197_);
  nand (_21963_, _21731_, _21197_);
  and (_21964_, _21963_, _21962_);
  or (_21965_, _21850_, _20994_);
  or (_21966_, _21965_, _21964_);
  nor (_21967_, _21195_, _26133_);
  and (_21969_, _21195_, _26133_);
  or (_21970_, _21969_, _21967_);
  and (_21971_, _21199_, _26129_);
  nor (_21972_, _21199_, _26129_);
  or (_21973_, _21972_, _21971_);
  or (_21974_, _21973_, _21970_);
  or (_21975_, _21974_, _21966_);
  or (_21976_, _21975_, _21961_);
  or (_21977_, _21976_, _21957_);
  nor (_21978_, _21920_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_21979_, _21978_, _21921_);
  nor (_21980_, _21979_, _22853_);
  and (_21981_, _21979_, _22853_);
  or (_21982_, _21981_, _21980_);
  or (_21983_, _21982_, _21977_);
  or (_21984_, _21983_, _21942_);
  or (_21985_, _21984_, _21941_);
  and (_21986_, _21927_, _22780_);
  nor (_21987_, _21921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_21988_, _21987_, _21922_);
  nor (_21989_, _21988_, _22772_);
  nor (_21990_, _21943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_21991_, _21990_, _21920_);
  and (_21992_, _21991_, _24590_);
  nor (_21993_, _21960_, _26118_);
  nor (_21994_, _21991_, _24590_);
  or (_21995_, _21994_, _21993_);
  or (_21996_, _21995_, _21992_);
  or (_21997_, _21996_, _21989_);
  and (_21998_, _21988_, _22772_);
  nor (_21999_, _21958_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22000_, _21999_, _21919_);
  and (_22001_, _22000_, _23972_);
  nor (_22002_, _22000_, _23972_);
  or (_22003_, _22002_, _22001_);
  or (_22004_, _22003_, _21998_);
  or (_22005_, _22004_, _21997_);
  or (_22006_, _22005_, _21986_);
  or (_22007_, _22006_, _21985_);
  or (_22008_, _22007_, _21938_);
  or (_22009_, _22008_, _21933_);
  and (_22010_, _22009_, _21918_);
  or (_22011_, _22010_, _21908_);
  or (_22012_, _22011_, _21771_);
  and (_22013_, _22012_, _21313_);
  nor (_22014_, _21442_, _22824_);
  and (_22015_, _21442_, _22824_);
  or (_22016_, _22015_, _22014_);
  nor (_22017_, _21664_, _24590_);
  and (_22018_, _21664_, _24590_);
  or (_22019_, _22018_, _22017_);
  or (_22020_, _22019_, _22016_);
  and (_22021_, _21616_, _22853_);
  nor (_22022_, _21616_, _22853_);
  or (_22023_, _22022_, _22021_);
  or (_22024_, _22023_, _20949_);
  or (_22025_, _22024_, _22020_);
  or (_22026_, _22025_, _21724_);
  or (_22027_, _20840_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_22028_, _20840_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22029_, _22028_, _22027_);
  nor (_22030_, _20879_, _26141_);
  and (_22031_, _20879_, _26141_);
  or (_22032_, _22031_, _22030_);
  or (_22033_, _22032_, _22029_);
  or (_22034_, _20758_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_22035_, _20758_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22036_, _22035_, _22034_);
  nor (_22037_, _20801_, _26133_);
  and (_22038_, _20801_, _26133_);
  or (_22039_, _22038_, _22037_);
  or (_22040_, _22039_, _22036_);
  or (_22041_, _22040_, _22033_);
  or (_22042_, _20674_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_22043_, _20674_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_22044_, _22043_, _22042_);
  nor (_22045_, _20716_, _22807_);
  and (_22046_, _20716_, _22807_);
  or (_22047_, _22046_, _22045_);
  or (_22048_, _22047_, _22044_);
  nor (_22049_, _20550_, _23972_);
  and (_22050_, _20550_, _23972_);
  or (_22051_, _22050_, _22049_);
  nor (_22052_, _20629_, _26118_);
  and (_22053_, _20629_, _26118_);
  or (_22054_, _22053_, _22052_);
  or (_22055_, _22054_, _22051_);
  or (_22056_, _22055_, _22048_);
  or (_22057_, _22056_, _22041_);
  or (_22058_, _22057_, _22026_);
  and (_22059_, _21397_, _21667_);
  and (_22060_, _22059_, _21571_);
  and (_22061_, _22060_, _21313_);
  and (_22062_, _22061_, _22058_);
  and (_22063_, _21539_, _20451_);
  and (_22064_, _21543_, _20432_);
  and (_22065_, _21535_, _20450_);
  or (_22066_, _22065_, _22064_);
  or (_22067_, _22066_, _22063_);
  and (_22068_, _21531_, _21288_);
  or (_22069_, _22068_, _20720_);
  or (_22070_, _22069_, _22067_);
  and (_22071_, _21555_, _20450_);
  or (_22072_, _22071_, _20458_);
  and (_22073_, _21563_, _20432_);
  and (_22074_, _21551_, _21288_);
  and (_22075_, _21559_, _20451_);
  or (_22076_, _22075_, _22074_);
  or (_22077_, _22076_, _22073_);
  or (_22078_, _22077_, _22072_);
  and (_22079_, _22078_, _22070_);
  and (_22080_, _22079_, _21286_);
  nand (_22081_, _22080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22082_, _22080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22083_, _22082_, _22081_);
  and (_22084_, _21521_, _20451_);
  and (_22085_, _21513_, _20450_);
  nor (_22086_, _22085_, _22084_);
  and (_22087_, _21509_, _21288_);
  and (_22088_, _21517_, _20432_);
  nor (_22089_, _22088_, _22087_);
  and (_22090_, _22089_, _22086_);
  nor (_22091_, _22090_, _20458_);
  and (_22092_, _21501_, _20451_);
  and (_22093_, _21493_, _20450_);
  nor (_22094_, _22093_, _22092_);
  and (_22095_, _21489_, _21288_);
  and (_22096_, _21497_, _20432_);
  nor (_22097_, _22096_, _22095_);
  and (_22098_, _22097_, _22094_);
  nor (_22099_, _22098_, _20720_);
  nor (_22100_, _22099_, _22091_);
  not (_22101_, _22100_);
  and (_22102_, _22101_, _21286_);
  and (_22103_, _22102_, _26133_);
  nor (_22104_, _22102_, _26133_);
  or (_22105_, _22104_, _22103_);
  or (_22106_, _22105_, _22083_);
  and (_22107_, _21370_, _20451_);
  or (_22108_, _22107_, _20720_);
  and (_22109_, _21366_, _20432_);
  and (_22110_, _21358_, _21288_);
  and (_22111_, _21362_, _20450_);
  or (_22112_, _22111_, _22110_);
  or (_22113_, _22112_, _22109_);
  or (_22114_, _22113_, _22108_);
  and (_22115_, _21382_, _20450_);
  and (_22116_, _21390_, _20451_);
  and (_22117_, _21386_, _20432_);
  or (_22118_, _22117_, _22116_);
  or (_22119_, _22118_, _22115_);
  and (_22120_, _21378_, _21288_);
  or (_22121_, _22120_, _20458_);
  or (_22122_, _22121_, _22119_);
  and (_22123_, _22122_, _22114_);
  and (_22124_, _22123_, _21286_);
  or (_22125_, _22124_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_22126_, _22124_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_22127_, _22126_, _22125_);
  and (_22128_, _21316_, _20450_);
  or (_22129_, _22128_, _20720_);
  and (_22130_, _21320_, _20432_);
  and (_22131_, _21330_, _21288_);
  or (_22132_, _22131_, _22130_);
  and (_22133_, _21324_, _20451_);
  or (_22134_, _22133_, _22132_);
  or (_22135_, _22134_, _22129_);
  and (_22136_, _21340_, _20450_);
  and (_22137_, _21336_, _20451_);
  and (_22138_, _21349_, _20432_);
  or (_22139_, _22138_, _22137_);
  or (_22140_, _22139_, _22136_);
  and (_22141_, _21345_, _21288_);
  or (_22142_, _22141_, _20458_);
  or (_22143_, _22142_, _22140_);
  and (_22144_, _22143_, _22135_);
  and (_22145_, _22144_, _21286_);
  nor (_22146_, _22145_, _26137_);
  and (_22147_, _22145_, _26137_);
  or (_22148_, _22147_, _22146_);
  or (_22149_, _22148_, _22127_);
  or (_22150_, _22149_, _22106_);
  and (_22151_, _21401_, _20450_);
  or (_22152_, _22151_, _20720_);
  and (_22153_, _21410_, _20432_);
  and (_22154_, _21406_, _21288_);
  or (_22155_, _22154_, _22153_);
  and (_22156_, _21415_, _20451_);
  or (_22157_, _22156_, _22155_);
  or (_22158_, _22157_, _22152_);
  and (_22159_, _21422_, _20450_);
  or (_22160_, _22159_, _20458_);
  and (_22161_, _21427_, _20432_);
  and (_22162_, _21432_, _21288_);
  and (_22163_, _21436_, _20451_);
  or (_22164_, _22163_, _22162_);
  or (_22165_, _22164_, _22161_);
  or (_22166_, _22165_, _22160_);
  and (_22167_, _22166_, _22158_);
  and (_22168_, _22167_, _21286_);
  nor (_22169_, _22168_, _26122_);
  and (_22170_, _22168_, _26122_);
  or (_22171_, _22170_, _22169_);
  and (_22172_, _21465_, _21288_);
  and (_22173_, _21477_, _20451_);
  and (_22174_, _21473_, _20432_);
  and (_22175_, _21469_, _20450_);
  or (_22176_, _22175_, _22174_);
  or (_22177_, _22176_, _22173_);
  or (_22178_, _22177_, _22172_);
  and (_22179_, _22178_, _20720_);
  and (_22180_, _21445_, _21288_);
  and (_22181_, _21457_, _20451_);
  and (_22182_, _21453_, _20432_);
  and (_22183_, _21449_, _20450_);
  or (_22184_, _22183_, _22182_);
  or (_22185_, _22184_, _22181_);
  or (_22186_, _22185_, _22180_);
  and (_22187_, _22186_, _20458_);
  or (_22188_, _22187_, _22179_);
  and (_22189_, _22188_, _21286_);
  and (_22190_, _22189_, _22807_);
  nor (_22191_, _22189_, _22807_);
  or (_22192_, _22191_, _22190_);
  or (_22193_, _22192_, _22171_);
  and (_22194_, _21585_, _21288_);
  and (_22195_, _21574_, _20432_);
  nor (_22196_, _22195_, _22194_);
  and (_22197_, _21589_, _20451_);
  and (_22198_, _21579_, _20450_);
  nor (_22199_, _22198_, _22197_);
  and (_22200_, _22199_, _22196_);
  and (_22201_, _22200_, _20458_);
  and (_22202_, _21610_, _20451_);
  and (_22203_, _21601_, _20450_);
  nor (_22204_, _22203_, _22202_);
  and (_22205_, _21596_, _20432_);
  and (_22206_, _21606_, _21288_);
  nor (_22207_, _22206_, _22205_);
  and (_22208_, _22207_, _22204_);
  and (_22209_, _22208_, _20720_);
  nor (_22210_, _22209_, _22201_);
  and (_22211_, _22210_, _21286_);
  nand (_22212_, _22211_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_22213_, _22211_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_22214_, _22213_, _22212_);
  and (_22215_, _21640_, _21288_);
  and (_22216_, _21652_, _20451_);
  and (_22217_, _21648_, _20432_);
  and (_22218_, _21644_, _20450_);
  or (_22219_, _22218_, _22217_);
  or (_22220_, _22219_, _22216_);
  or (_22221_, _22220_, _22215_);
  and (_22222_, _22221_, _20720_);
  and (_22223_, _21620_, _21288_);
  and (_22224_, _21632_, _20451_);
  and (_22225_, _21628_, _20432_);
  and (_22226_, _21624_, _20450_);
  or (_22227_, _22226_, _22225_);
  or (_22228_, _22227_, _22224_);
  or (_22229_, _22228_, _22223_);
  and (_22230_, _22229_, _20458_);
  or (_22231_, _22230_, _22222_);
  and (_22232_, _22231_, _21286_);
  nand (_22233_, _22232_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_22234_, _22232_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_22235_, _22234_, _22233_);
  or (_22236_, _22235_, _22214_);
  or (_22237_, _22236_, _22193_);
  or (_22238_, _22237_, _22150_);
  or (_22239_, _20840_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_22240_, _20840_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_22241_, _22240_, _22239_);
  and (_22242_, _20879_, _22824_);
  nor (_22243_, _20879_, _22824_);
  or (_22244_, _22243_, _22242_);
  or (_22245_, _22244_, _22241_);
  or (_22246_, _20758_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_22247_, _20758_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_22248_, _22247_, _22246_);
  nor (_22249_, _20801_, _22853_);
  and (_22250_, _20801_, _22853_);
  or (_22251_, _22250_, _22249_);
  or (_22252_, _22251_, _22248_);
  or (_22253_, _22252_, _22245_);
  or (_22254_, _20674_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_22255_, _20674_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22256_, _22255_, _22254_);
  and (_22257_, _20716_, _22776_);
  nor (_22258_, _20716_, _22776_);
  or (_22259_, _22258_, _22257_);
  or (_22260_, _22259_, _22256_);
  and (_22261_, _20550_, _04718_);
  nor (_22262_, _20550_, _04718_);
  or (_22263_, _22262_, _22261_);
  and (_22264_, _20629_, _22784_);
  nor (_22265_, _20629_, _22784_);
  or (_22266_, _22265_, _22264_);
  or (_22267_, _22266_, _22263_);
  or (_22268_, _22267_, _22260_);
  or (_22269_, _22268_, _22253_);
  or (_22270_, _22269_, _22238_);
  and (_22271_, _21801_, _21697_);
  and (_22272_, _22271_, _21313_);
  and (_22273_, _22272_, _22270_);
  or (_22274_, _22273_, _22062_);
  or (_22275_, _22274_, _22013_);
  or (property_invalid, _22275_, _21663_);
  and (_22276_, _13696_, _23718_);
  and (_22277_, _13698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or (_12449_, _22277_, _22276_);
  and (_22278_, _13690_, _23982_);
  and (_22279_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_27190_, _22279_, _22278_);
  and (_22280_, _02845_, _23982_);
  and (_22281_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_12454_, _22281_, _22280_);
  and (_22282_, _17972_, _23718_);
  and (_22283_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_12457_, _22283_, _22282_);
  and (_22284_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  and (_22285_, _02450_, _23635_);
  or (_12458_, _22285_, _22284_);
  and (_22286_, _05287_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_22287_, _24479_, _24486_);
  or (_22288_, _17153_, _22287_);
  or (_22289_, _22288_, _17164_);
  or (_22290_, _22289_, _24501_);
  or (_22291_, _26600_, _05307_);
  or (_22292_, _26711_, _26703_);
  and (_22293_, _24453_, _24486_);
  or (_22294_, _17172_, _22293_);
  or (_22295_, _22294_, _22292_);
  or (_22296_, _22295_, _22291_);
  and (_22297_, _24486_, _24391_);
  not (_22298_, _26707_);
  or (_22299_, _22298_, _26685_);
  or (_22300_, _22299_, _22297_);
  or (_22301_, _22300_, _17185_);
  or (_22302_, _22301_, _22296_);
  or (_22303_, _22302_, _22290_);
  and (_22304_, _22303_, _25615_);
  or (_26876_[0], _22304_, _22286_);
  and (_22305_, _21307_, first_instr);
  or (_00000_, _22305_, rst);
  and (_22306_, _13736_, _23635_);
  and (_22307_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_12464_, _22307_, _22306_);
  and (_22308_, _03296_, _23755_);
  and (_22309_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_27167_, _22309_, _22308_);
  and (_22310_, _17972_, _23791_);
  and (_22311_, _17974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_12480_, _22311_, _22310_);
  and (_22312_, _13846_, _23755_);
  and (_22313_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or (_27198_, _22313_, _22312_);
  and (_22314_, _06255_, _23982_);
  and (_22315_, _06257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or (_12483_, _22315_, _22314_);
  and (_22316_, _24777_, _23635_);
  and (_22317_, _24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_12495_, _22317_, _22316_);
  and (_22318_, _02845_, _23838_);
  and (_22319_, _02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_12497_, _22319_, _22318_);
  and (_22320_, _15909_, _23755_);
  and (_22321_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_12504_, _22321_, _22320_);
  and (_22322_, _15485_, _23589_);
  and (_22323_, _15487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or (_12506_, _22323_, _22322_);
  and (_22324_, _13846_, _23718_);
  and (_22325_, _13848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or (_12518_, _22325_, _22324_);
  and (_22326_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  and (_22327_, _02450_, _23982_);
  or (_12523_, _22327_, _22326_);
  and (_22328_, _06264_, _23589_);
  and (_22329_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_12532_, _22329_, _22328_);
  or (_22330_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_22331_, _22330_, _22761_);
  nand (_22332_, _23889_, _23784_);
  and (_12541_, _22332_, _22331_);
  nand (_22333_, _23884_, _23669_);
  or (_22334_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_22335_, _22334_, _22761_);
  and (_12546_, _22335_, _22333_);
  and (_22336_, _02322_, _23676_);
  and (_22337_, _02324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_12555_, _22337_, _22336_);
  or (_22338_, _17236_, _17232_);
  and (_22339_, _22338_, _22768_);
  and (_22340_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_22341_, _22340_, _17251_);
  or (_22342_, _22341_, _22339_);
  and (_26877_[0], _22342_, _22761_);
  and (_22343_, _06264_, _23755_);
  and (_22344_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_12559_, _22344_, _22343_);
  and (_22345_, _24622_, _23718_);
  and (_22346_, _24624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_27200_, _22346_, _22345_);
  and (_22347_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_22348_, _22347_, _17250_);
  and (_22349_, _22348_, _22761_);
  and (_22350_, _26716_, _24445_);
  or (_22351_, _22350_, _26664_);
  or (_22352_, _22351_, _17133_);
  or (_22353_, _22352_, _17239_);
  and (_22354_, _22353_, _25615_);
  or (_26877_[1], _22354_, _22349_);
  and (_22355_, _02451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  and (_22356_, _02450_, _23838_);
  or (_12563_, _22356_, _22355_);
  and (_22357_, _03358_, _23676_);
  and (_22358_, _03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or (_12564_, _22358_, _22357_);
  nand (_22359_, _23988_, _23784_);
  not (_22360_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_22361_, _24017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_22362_, _22361_, _24032_);
  and (_22363_, _22362_, _23996_);
  nor (_22364_, _22363_, _22360_);
  and (_22365_, _22363_, _22360_);
  or (_22366_, _22365_, _22364_);
  and (_22367_, _22366_, _23999_);
  and (_22368_, _24039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_22369_, _22368_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_22370_, _13639_);
  and (_22371_, _22370_, _24038_);
  and (_22372_, _22371_, _22369_);
  and (_22373_, _24050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_22374_, _22373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_22375_, _13634_, _24053_);
  and (_22376_, _22375_, _22374_);
  or (_22377_, _22376_, _22372_);
  or (_22378_, _22377_, _22367_);
  or (_22379_, _22378_, _23988_);
  and (_22380_, _22379_, _23995_);
  and (_22381_, _22380_, _22359_);
  and (_22382_, _23994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_22383_, _22382_, _22381_);
  and (_12568_, _22383_, _22761_);
  or (_22384_, _24034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_22385_, _22384_, _23999_);
  nor (_22386_, _22385_, _22363_);
  or (_22387_, _24039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_22388_, _22387_, _24038_);
  nor (_22389_, _22388_, _22368_);
  or (_22390_, _24023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_22391_, _22373_, _24054_);
  and (_22392_, _22391_, _22390_);
  or (_22393_, _22392_, _22389_);
  or (_22394_, _22393_, _22386_);
  or (_22395_, _22394_, _23988_);
  nand (_22396_, _23988_, _23669_);
  and (_22397_, _22396_, _22395_);
  or (_22398_, _22397_, _23994_);
  or (_22399_, _23995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_22400_, _22399_, _22761_);
  and (_12570_, _22400_, _22398_);
  and (_22401_, _13864_, _23635_);
  and (_22402_, _13866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_12575_, _22402_, _22401_);
  and (_22403_, _26728_, _25924_);
  or (_22404_, _26572_, _24472_);
  or (_22405_, _22404_, _22403_);
  and (_22406_, _02005_, _24489_);
  or (_22407_, _02260_, _22293_);
  or (_22408_, _22407_, _22406_);
  or (_22409_, _22408_, _22405_);
  or (_22410_, _17240_, _24488_);
  or (_22411_, _22410_, _24536_);
  or (_22412_, _22411_, _17133_);
  or (_22413_, _22412_, _22409_);
  or (_22414_, _24513_, _24420_);
  or (_22415_, _22414_, _24463_);
  or (_22416_, _22415_, _26653_);
  or (_22417_, _22416_, _02265_);
  or (_22418_, _22417_, _22413_);
  or (_22419_, _02006_, _24519_);
  or (_22420_, _02024_, _26821_);
  or (_22421_, _22420_, _22419_);
  and (_22422_, _02038_, _25924_);
  or (_22423_, _22422_, _24507_);
  or (_22424_, _17237_, _26819_);
  or (_22425_, _22424_, _02242_);
  or (_22426_, _22425_, _22423_);
  or (_22427_, _22426_, _22421_);
  or (_22428_, _22427_, _22418_);
  and (_22429_, _22428_, _22768_);
  and (_22430_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_22431_, _26824_, _24538_);
  or (_22432_, _22431_, _22430_);
  or (_22433_, _22432_, _22429_);
  and (_26878_[0], _22433_, _22761_);
  and (_22434_, _15537_, _23676_);
  and (_22435_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_12578_, _22435_, _22434_);
  and (_22436_, _15909_, _23718_);
  and (_22437_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_26976_, _22437_, _22436_);
  nand (_22438_, _23988_, _23748_);
  and (_22439_, _13606_, _24004_);
  or (_22440_, _22439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_22441_, _13606_, _24005_);
  and (_22442_, _22441_, _23998_);
  and (_22443_, _22442_, _22440_);
  and (_22444_, _24050_, _24004_);
  or (_22445_, _22444_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_22446_, _24051_, _24054_);
  and (_22447_, _22446_, _22445_);
  and (_22448_, _24039_, _24004_);
  and (_22449_, _22448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_22450_, _22449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_22451_, _22449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_22452_, _22451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_22453_, _22452_, _22450_);
  or (_22454_, _22453_, _22447_);
  or (_22455_, _22454_, _22443_);
  or (_22456_, _22455_, _23988_);
  and (_22457_, _22456_, _23995_);
  and (_22458_, _22457_, _22438_);
  and (_22459_, _23994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_22460_, _22459_, _22458_);
  and (_12591_, _22460_, _22761_);
  nand (_22461_, _23988_, _23628_);
  and (_22462_, _24039_, _24003_);
  or (_22463_, _22462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_22464_, _22448_);
  and (_22465_, _22464_, _24038_);
  and (_22466_, _22465_, _22463_);
  not (_22467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_22468_, _24034_, _24003_);
  nor (_22469_, _22468_, _22467_);
  and (_22470_, _22468_, _22467_);
  or (_22471_, _22470_, _22469_);
  and (_22472_, _22471_, _23999_);
  and (_22473_, _13636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_22474_, _22473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_22475_, _22474_, _22467_);
  nor (_22476_, _22444_, _24054_);
  and (_22477_, _22476_, _22475_);
  or (_22478_, _22477_, _22472_);
  or (_22479_, _22478_, _22466_);
  or (_22480_, _22479_, _23988_);
  and (_22481_, _22480_, _23995_);
  and (_22482_, _22481_, _22461_);
  and (_22483_, _23994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_22484_, _22483_, _22482_);
  and (_12594_, _22484_, _22761_);
  nand (_22485_, _23988_, _23914_);
  or (_22486_, _22473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_22487_, _22474_, _24053_);
  and (_22488_, _22487_, _22486_);
  and (_22489_, _24034_, _24002_);
  or (_22490_, _22489_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_22491_, _22490_, _23999_);
  nor (_22492_, _22491_, _22468_);
  and (_22493_, _24039_, _24002_);
  or (_22494_, _22493_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_22495_, _22462_);
  and (_22496_, _22495_, _24038_);
  and (_22497_, _22496_, _22494_);
  or (_22498_, _22497_, _22492_);
  or (_22499_, _22498_, _22488_);
  or (_22500_, _22499_, _23988_);
  and (_22501_, _22500_, _23995_);
  and (_22502_, _22501_, _22485_);
  and (_22503_, _23994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_22504_, _22503_, _22502_);
  and (_12596_, _22504_, _22761_);
  nand (_22505_, _23988_, _23832_);
  and (_22506_, _13629_, _23996_);
  or (_22507_, _22506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_22508_, _22506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_22509_, _22508_, _23999_);
  and (_22510_, _22509_, _22507_);
  and (_22511_, _24039_, _24001_);
  or (_22512_, _22511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_22513_, _22493_);
  and (_22514_, _22513_, _24038_);
  and (_22515_, _22514_, _22512_);
  or (_22516_, _13636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_22517_, _22473_, _24054_);
  and (_22518_, _22517_, _22516_);
  or (_22519_, _22518_, _22515_);
  or (_22520_, _22519_, _22510_);
  or (_22521_, _22520_, _23988_);
  and (_22522_, _22521_, _23995_);
  and (_22523_, _22522_, _22505_);
  and (_22524_, _23994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_22525_, _22524_, _22523_);
  and (_12598_, _22525_, _22761_);
  and (_22526_, _15537_, _23589_);
  and (_22527_, _15539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_12602_, _22527_, _22526_);
  and (_22528_, _15909_, _23791_);
  and (_22529_, _15911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_12604_, _22529_, _22528_);
  and (_22530_, _03296_, _23718_);
  and (_22531_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_12607_, _22531_, _22530_);
  or (_22532_, _23995_, _23709_);
  nor (_22533_, _24047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_22534_, _22533_, _24048_);
  and (_22535_, _13607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_22536_, _22535_, _22534_);
  nor (_22537_, _22536_, _23988_);
  and (_22538_, _23988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_22539_, _22538_, _22537_);
  or (_22540_, _22539_, _23994_);
  and (_22541_, _22540_, _22761_);
  and (_12614_, _22541_, _22532_);
  nor (_22542_, _24046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_22543_, _22542_, _24047_);
  and (_22544_, _13607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_22545_, _22544_, _22543_);
  nor (_22546_, _22545_, _23988_);
  and (_22547_, _23988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_22548_, _22547_, _22546_);
  and (_22549_, _22548_, _23995_);
  nor (_22550_, _23995_, _23784_);
  or (_22551_, _22550_, _22549_);
  and (_12616_, _22551_, _22761_);
  nor (_22552_, _24017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_22553_, _22552_, _24046_);
  and (_22554_, _22362_, _23997_);
  nor (_22555_, _22554_, _22553_);
  nor (_22556_, _22555_, _23988_);
  and (_22557_, _23988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_22558_, _22557_, _22556_);
  and (_22559_, _22558_, _23995_);
  and (_22560_, _23994_, _24763_);
  or (_22561_, _22560_, _22559_);
  and (_12623_, _22561_, _22761_);
  and (_22562_, _13736_, _23676_);
  and (_22563_, _13738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_27199_, _22563_, _22562_);
  and (_22564_, _16707_, _23676_);
  and (_22565_, _16709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_12626_, _22565_, _22564_);
  and (_22566_, _24491_, _24458_);
  nor (_22567_, _22566_, _24497_);
  nand (_22568_, _22567_, _26662_);
  or (_22569_, _17223_, _26735_);
  or (_22570_, _22569_, _22568_);
  not (_22571_, _26706_);
  or (_22572_, _22571_, _26683_);
  or (_22573_, _26728_, _24472_);
  or (_22574_, _22573_, _22572_);
  or (_22575_, _22574_, _22423_);
  or (_22576_, _22575_, _22570_);
  and (_22577_, _22424_, _24346_);
  or (_22578_, _22577_, _22416_);
  or (_22579_, _22578_, _22576_);
  or (_22580_, _22579_, _22421_);
  and (_22581_, _22580_, _22768_);
  and (_22582_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_22583_, _22582_, _22431_);
  or (_22584_, _22583_, _22581_);
  and (_26878_[1], _22584_, _22761_);
  and (_22585_, _13690_, _23755_);
  and (_22586_, _13692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_12631_, _22586_, _22585_);
  nand (_22587_, _23994_, _23914_);
  nand (_22588_, _13607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_22589_, _13602_);
  or (_22590_, _22589_, _24050_);
  and (_22591_, _22590_, _22588_);
  nor (_22592_, _22591_, _23988_);
  nand (_22593_, _13625_, _24050_);
  and (_22594_, _22593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_22595_, _22594_, _22592_);
  or (_22596_, _22595_, _23994_);
  and (_22597_, _22596_, _22761_);
  and (_12633_, _22597_, _22587_);
  and (_22598_, _24054_, _24050_);
  nand (_22599_, _22598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_22600_, _22599_, _23988_);
  and (_22601_, _22600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_22602_, _13607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_22603_, _22599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_22604_, _22603_, _22602_);
  nor (_22605_, _22604_, _23988_);
  or (_22606_, _22605_, _22601_);
  and (_22607_, _22606_, _23995_);
  nor (_22608_, _23995_, _23748_);
  or (_22609_, _22608_, _22607_);
  and (_12643_, _22609_, _22761_);
  and (_22610_, _06264_, _23718_);
  and (_22611_, _06267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_12645_, _22611_, _22610_);
  and (_22612_, _22600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand (_22613_, _13607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_22614_, _22599_, _22598_);
  and (_22615_, _22614_, _22613_);
  nor (_22616_, _22615_, _23988_);
  or (_22617_, _22616_, _22612_);
  and (_22618_, _22617_, _23995_);
  nor (_22619_, _23995_, _23628_);
  or (_22620_, _22619_, _22618_);
  and (_12647_, _22620_, _22761_);
  and (_22621_, _05323_, _23755_);
  and (_22622_, _05325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or (_12649_, _22622_, _22621_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _26852_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _26852_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _26852_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _26852_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _26852_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _26852_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _26852_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _26852_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _26868_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _26851_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _26851_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _26851_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _26851_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _26851_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _26851_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _26851_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _26851_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _26851_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _26851_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _26851_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _26851_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _26851_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _26851_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _26851_[15]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _26859_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _26859_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _26859_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _26859_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _26859_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _26859_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _26859_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _26859_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _26860_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _26860_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _26860_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _26860_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _26860_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _26860_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _26860_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _26860_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _26861_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _26861_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _26861_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _26861_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _26861_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _26861_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _26861_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _26861_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _26862_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _26862_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _26862_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _26862_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _26862_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _26862_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _26862_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _26862_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _26863_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _26863_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _26863_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _26863_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _26863_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _26863_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _26863_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _26863_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _26864_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _26864_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _26864_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _26864_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _26864_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _26864_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _26864_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _26864_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _26865_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _26865_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _26865_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _26865_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _26865_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _26865_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _26865_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _26865_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _26866_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _26866_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _26866_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _26866_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _26866_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _26866_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _26866_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _26866_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _26867_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _26867_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _26867_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _26867_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _26867_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _26867_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _26867_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _26867_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _26853_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _26853_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _26853_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _26853_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _26853_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _26853_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _26853_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _26853_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _26854_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _26854_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _26854_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _26854_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _26854_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _26854_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _26854_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _26854_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _26855_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _26855_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _26855_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _26855_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _26855_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _26855_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _26855_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _26855_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _26856_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _26856_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _26856_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _26856_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _26856_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _26856_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _26856_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _26856_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _26857_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _26857_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _26857_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _26857_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _26857_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _26857_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _26857_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _26857_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _26858_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _26858_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _26858_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _26858_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _26858_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _26858_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _26858_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _26858_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _11536_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _11516_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _09091_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _11482_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _11532_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _09097_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _09101_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _09083_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _11757_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11646_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _11734_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11721_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _11764_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _11755_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _11644_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _09094_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11972_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22694_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11983_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _12219_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11988_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _12000_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11977_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11990_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11996_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _12002_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11998_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11992_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11985_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _12009_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _12005_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _12028_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _26869_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _26869_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _26869_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _26869_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _26869_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _26869_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _26869_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _26869_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _26896_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _26896_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _26896_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _26896_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _26896_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _26896_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _26896_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _26896_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _26906_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _26906_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _26906_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _26906_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _26906_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _26906_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _26906_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _26906_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _26876_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _26876_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _26877_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _26877_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _26877_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _26878_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _26878_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _26878_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _26879_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _26879_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _26880_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _26880_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _26880_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _26880_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _26881_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _26881_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _26882_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _26870_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _26870_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _26870_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _26871_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _26871_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _26871_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _26872_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _26872_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _26873_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _26873_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _26873_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _26873_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _26873_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _26873_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _26873_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _26873_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _26874_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _26875_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _26875_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _26921_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _26883_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _26883_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _26883_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _26883_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _26883_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _26883_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _26883_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _26883_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _26884_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _26884_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _26884_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _26884_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _26884_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _26884_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _26884_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _26884_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _26885_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _26885_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _26885_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _26885_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _26885_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _26885_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _26885_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _26885_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _26886_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _26886_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _26886_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _26886_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _26886_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _26886_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _26886_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _26886_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _26887_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _26887_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _26887_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _26887_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _26887_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _26887_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _26887_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _26887_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _26888_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _26888_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _26888_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _26888_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _26888_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _26888_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _26888_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _26888_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _26889_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _26889_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _26889_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _26889_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _26889_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _26889_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _26889_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _26889_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _26890_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _26890_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _26890_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _26890_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _26890_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _26890_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _26890_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _26890_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _26894_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _26894_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _26894_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _26894_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _26894_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _26891_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _26891_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _26891_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _26891_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _26891_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _26891_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _26891_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _26891_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _26891_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _26891_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _26891_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _26891_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _26891_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _26891_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _26891_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _26891_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _26892_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26892_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26892_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _26892_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _26892_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _26892_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _26892_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _26892_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _26892_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _26892_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _26892_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26892_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _26892_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _26892_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _26892_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _26892_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _26912_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _26912_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _26912_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _26912_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _26912_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _26912_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _26912_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _26912_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _26912_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _26912_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _26912_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _26912_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _26912_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _26912_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _26912_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _26912_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _26912_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _26912_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _26912_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _26912_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _26912_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _26912_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _26912_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _26912_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _26912_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _26912_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _26912_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _26912_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _26912_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _26912_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _26912_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _26912_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _26893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _26895_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _26895_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _26895_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _26895_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _26895_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _26895_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _26895_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _26895_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _26897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _26898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _26899_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _26899_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _26899_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _26899_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _26899_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _26899_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _26899_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _26899_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _26899_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _26899_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _26899_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _26899_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _26899_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _26899_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _26899_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _26899_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _26900_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _26900_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _26900_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _26900_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _26900_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _26900_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _26900_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _26900_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _26900_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _26900_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _26900_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _26900_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _26900_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _26900_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _26900_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _26900_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _26901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _26903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _26902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _26904_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _26904_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _26904_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _26904_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _26904_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _26904_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _26904_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _26904_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _26905_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26905_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _26905_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _26907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _26908_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _26908_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _26908_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _26908_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _26908_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _26908_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _26908_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _26908_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _26909_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _26910_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _26911_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _26911_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _26911_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _26911_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _26913_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _26913_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _26913_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _26913_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _26913_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _26913_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _26913_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _26913_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _26913_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _26913_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _26913_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _26913_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _26913_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _26913_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _26913_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _26913_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _26913_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _26913_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _26913_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _26913_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _26913_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _26913_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _26913_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _26913_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _26913_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _26913_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _26913_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _26913_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _26913_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _26913_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _26913_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _26913_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _26914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _26915_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _26916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _26917_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _26917_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _26917_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _26917_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _26918_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _26919_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26920_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26920_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26920_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26920_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26920_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26920_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26920_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _26920_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _26922_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _26922_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _26922_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _22666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _22690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _22688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _22686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _11431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _22658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _22657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _22655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _11435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _26989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _26990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _26991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _22701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _22700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _26992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _22663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _22806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _26966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _11888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _11588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _22740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _22739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _22738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _22743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _22907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _22888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _11886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _23079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _26945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _26946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _22746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _22745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _22661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _27024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _11917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _11569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _11685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _22643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _27025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _22645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _11869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _23357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _11864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _23204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _23186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _23173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _23250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _11877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _04225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _27187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _27188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _27189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _27190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _04298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _12631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _04821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _04389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _04399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _12449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _04462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _04485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _27170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _27171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _04236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _27150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _05098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _05094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _27151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _05150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _12575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _27152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _05192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _27236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _10127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _11913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _11921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _11915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _12495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _25747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _10160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _10120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _01039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _02258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _27234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _27235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _07420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _03957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _10138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _10089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _07547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _04607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _10105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _05285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _07423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _27233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _23036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _07864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _27230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _27231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _27232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _10070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _07082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _07023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _09283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _07783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _08627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _10038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _10030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _11680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _11079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _12096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _10046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _27229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _09997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _26525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _10866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _08507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _08510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _10025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _08464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _12555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _10523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _07434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _08301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _23686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _06378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _07432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _22680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _08529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _09922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _27227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _09963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _27228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _07437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _01568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _03339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _09607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _11240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _09750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _11237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _09775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _11392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _01076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _12109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _27223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _09325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _27224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _27225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _11242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _09452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _11346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _09490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _08972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _27222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _08996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _11352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _09029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _09049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _11247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _11394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _08956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _09130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _10073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _08954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _10080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _27314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _08951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _10110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _27312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _09983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _08965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _27313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _10019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _08961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _10034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _08959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _11068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _27311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _11116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _11097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _11119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _11102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _09925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _08968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _08593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _11180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _11149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _11187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _11151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _11161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _27310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _11063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _10843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _10869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _07882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _27308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _10876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _10890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _10897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _27309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _07892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _10807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _07890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _10811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _08607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _10828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _07887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _10832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _27307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _07902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _10716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _07899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _10721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _08701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _10756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _07896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _10628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _07909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _27306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _07907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _10653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _08705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _08790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _10679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _11803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _27275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _10845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _12497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _12454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _27276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _27277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _09235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _10504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _27304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _07916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _10561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _07914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _10576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _27305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _10609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _09056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _10895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _26938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _08800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _09115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _11170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _11192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _11154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _08815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _10830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _26936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _10840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _10861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _08806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _10880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _26937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _10727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _09062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _10737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _26933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _10792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _26934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _26935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _09118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _26930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _10669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _08844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _26931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _10676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _08842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _26932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _10713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _07202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _05713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _26949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _07098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _05702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _07106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _26950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _06128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _08718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _07141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _08761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _09053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _26948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _09140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _07017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _09148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _07169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _07463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _07499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _07067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _07221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _07789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _07923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _07046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _06321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _27193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _24205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _06048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _06034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _06032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _06135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _06134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _06394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _06559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _06520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _24230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _25057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _06180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _06221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _06182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _27191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _27192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _06643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _01731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _06713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _06689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _01718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _06461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _06986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _01690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _07089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _01684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _06808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _06785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _01711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _06888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _11642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _26007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _24345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _05587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _26031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _26009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _24543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _25232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _25112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _25957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _27186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _25944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _22669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _00741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _00515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _25962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _09823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _10782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _25939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _24548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _25973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _24512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _02551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _02464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _07300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _07294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _01659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _27184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _25225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _27185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _22750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _12167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _07404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _07445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _07489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _07454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _24284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _07189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _07175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _01677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _24293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _07552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _07544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _01633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _27183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _07805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _24287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _07395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _09071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _08985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _27182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _08177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _08163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _08160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _08730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _08726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _09152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _09788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _09988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _01523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _08821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _08819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _08812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _27181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _08574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _27274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _10838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _26763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _26738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _07298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _09565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _09529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _27179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _27180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _10849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _24312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _10141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _01520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _10233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _01518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _27175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _11206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _27176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _27177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _27178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _11100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _00414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _25229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _11853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _11974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _27172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _00167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _27173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _11501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _27174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _00243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _12564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _00079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _27168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _00154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _12198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _27169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _24530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _11882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _11129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _24339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _12607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _11962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _00051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _24532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _27167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _00142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _02584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _23331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _23516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _02406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _27165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _27166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _10418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _00049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _27162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _27163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _10254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _05731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _02417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _27164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _11698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _23157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _11691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _02435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _12211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _02433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _12483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _02597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _27160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _27161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _25831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _11952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _02448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _27159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _02445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _06650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _02600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _22687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _22671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _27156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _02455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _22668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _27157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _06925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _02605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _27158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _07809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _25757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _27273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _26573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _22793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _23085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _23094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _07304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _27155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _22678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _22676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _02470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _22675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _02467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _22674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _02612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _02620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _22685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _02489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _22684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _02617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _22683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _22679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _02476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _19788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _07318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _22670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _22672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _22673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _27268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _27269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _01998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _07311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _27271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _22705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _22710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _22681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _27272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _22682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _10818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _02657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _27153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _22706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _02507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _22703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _27154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _22698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _22696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _27149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _02577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _08878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _02569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _08295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _02661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _00266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _26793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _22749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _02511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _22748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _02627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _27148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _04891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _02574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _09392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _27266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _01283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _01221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _10724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _07495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _23559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _24315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _23600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _00823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _00898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _00854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _10745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _27267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _11898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _10780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _13746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _09439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _07335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _27261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _27262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _04770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _04762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _04755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _05136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _05003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _10673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _27263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _03488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _03422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _27264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _04611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _10688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _11610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _25347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _25326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _27112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _25396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _11490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _25007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _25096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _07342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _09781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _09706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _09668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _10442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _10639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _08175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _06744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _26923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _11762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _26924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _25514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _11492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _25439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _11766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _25475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _24333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _24326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _11808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _24177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _24175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _24167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _24163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _24212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _24355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _24370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _27226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _11798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _24442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _11796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _11605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _24298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _27207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _11779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _24504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _24498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _24477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _11784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _24535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _24551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _27292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _23764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _23761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _27293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _23860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _23856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _11847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _23421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _11837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _23912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _23965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _23960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _11841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _27270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _24014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _24008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _24208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _24202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _11450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _11639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _24079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _11839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _24143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _24114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _23396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _23689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _23679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _23450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _11856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _11591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _11688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _23294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _02529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _27147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _02523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _23097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _02631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _23026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _02515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _22961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _26669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _02637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _26613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _26527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _02534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _27145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _25737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _27146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _02555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _26734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _02653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _26704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _26684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _02541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _27144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _26678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _05086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _24444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _05089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _05310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _24467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _27143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _05174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _24462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _05114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _05107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _05118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _24437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _27142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _24151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _04999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _24157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _04620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _03366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _27140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _05277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _05224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _27141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _05015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _05033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _04523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _04536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _03371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _04553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _03575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _04567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _04586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _04605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _04420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _04441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _27138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _27139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _03387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _04478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _03578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _04498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _04333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _03585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _04346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _04377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _03581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _04392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _04412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _03398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _04249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _04283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _03428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _03676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _04292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _04307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _03419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _04322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _27136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _04201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _03458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _27137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _03598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _04221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _04244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _03444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _27134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _27135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _04113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _03468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _04125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _04144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _03465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _04164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _03751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _27132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _03559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _03768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _03820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _27133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _03835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _03551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _04032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _27130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _04041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _04050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _27131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _04102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _03481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _03748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _03962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _03520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _27128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _03693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _27129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _03999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _03500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _04021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _03542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _03870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _03642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _03904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _03913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _03926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _03523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _27127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _24609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _24589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _24553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _25300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _25293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _25287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _05121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _24434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _05112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _25318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _25350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _25330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _05116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _25393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _25421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _25404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _27124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _24082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _24076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _24188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _24185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _24173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _05041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _25460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _27123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _25854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _24249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _24290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _05024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _24320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _24342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _24323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _25490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _25527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _25524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _25511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _05275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _25719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _25714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _05231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _04616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _27121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _25545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _05243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _25623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _25567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _27122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _25500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _04610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _01310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _01242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _27120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _10616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _09583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _24781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _00808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _27118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _02136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _04600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _03209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _03164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _04594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _27119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _01095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _09632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _09616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _02844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _04680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _04618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _04503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _04862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _27117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _04540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _10569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _10607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _04531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _08609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _07862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _05337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _05279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _04495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _10758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _10754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _27113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _27114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _27115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _27116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _10368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _22786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _04482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _03182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _11217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _11201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _11085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _12175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _12158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _23053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _22742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _27110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _12563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _12523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _12458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _04492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _22708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _04445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _01382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _01364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _04438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _03186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _27109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _01092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _04475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _01431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _01423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _04431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _03689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _03661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _03026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _27108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _25065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _02949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _27107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _05139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _04417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _06923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _06762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _04404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _03194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _09271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _27104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _04373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _27105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _08682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _27106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _08941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _08937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _09362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _09329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _10528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _27103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _09701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _02955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _09198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _09194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _04328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _27101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _27102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _10787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _11289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _11577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _02959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _09421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _11285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _04311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _22760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _27099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _27100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _11919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _11891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _04331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _03289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _00913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _02270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _02219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _04301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _04082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _04900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _27098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _27097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _06556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _06741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _06698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _04288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _09406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _08884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _04281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _08570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _02995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _27093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _22704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _12186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _27094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _07526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _23144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _22707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _22935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _26586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _02997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _08849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _27092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _08543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _08552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _23675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _10287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _04213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _03224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _08517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _27091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _08500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _04233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _04732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _04716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _04209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _22845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _04198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _09562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _27090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _04218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _07791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _25851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _09018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _04192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _07159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _23539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _04189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _10536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _10223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _07925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _10226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _27303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _10332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _07920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _10391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _10453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _09811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _09835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _09894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _08184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _09912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _08733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _27302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _10209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _08717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _10168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _27301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _09752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _08201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _09767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _09725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _08203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _10066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _10092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _08721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _27299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _27300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _07936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _10136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _07934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _09978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _09995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _27297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _08167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _10036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _08161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _27298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _08723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _25732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _25648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _11090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _23727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _09920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _09959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _08172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _09969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _00329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _00278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _00107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _11114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _27296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _25114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _25022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _25817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _25726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _27295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _22642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _00743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _11108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _26162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _26374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _26223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _11638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _20210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _14343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _11048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _11213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _25427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _27294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _04354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _27288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _11168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _27289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _27290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _11144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _27291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _01856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _24563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _27286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _01170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _11196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _01878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _01818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _01582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _11141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _27287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _27281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _07471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _07874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _27282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _11182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _27283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _27284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _27285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _10905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _11257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _11245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _07283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _04729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _04721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _11051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _11065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _11372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _11344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _11428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _11424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _11410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _27280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _11112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _11125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _12626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _07291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _27278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _11554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _27279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _11911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _11859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _10878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _08021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _04943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _08411_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _03842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _09838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _27242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _09897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _07442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _11408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _27221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _11263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _08658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _11364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _08780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _08852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _11255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _07452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _09233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _22665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _09729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _14495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _09150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _07868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _09821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _27220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _08374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _11280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _08392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _11366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _08475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _08595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _11265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _27240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _27241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _11935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _09754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _21947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _09746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _11111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _11495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _11287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _11397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _08181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _11283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _08224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _11370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _27218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _27219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _27237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _11774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _11816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _27238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _10729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _10611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _10567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _27239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _07877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _11294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _27215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _27216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _07976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _27217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _08063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _11291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _27212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _27213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _11329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _11405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _07709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _27214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _11297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _07831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _27209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _27210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _07484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _11307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _07516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _07690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _11412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _27211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _27208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _11403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _06935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _07105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _11312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _07183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _11310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _07210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _11320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _27203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _11386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _27204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _27205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _27206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _06852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _11317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _04577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _04590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _27200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _04574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _27201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _11325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _27202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _11388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _27199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _04317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _12404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _04324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _04550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _12464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _04555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _04546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _04647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _27197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _12518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _04694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _04691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _04669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _27198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _04543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _04748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _04745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _04725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _04723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _04788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _04784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _04782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _12506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _20400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _19939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _21968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _21895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _21584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _11943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _18030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _17708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _12578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _04885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _04877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _04872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _04941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _04934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _04927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _12602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _09798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _09847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _08976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _09889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _08973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _09900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _09112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _09142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _22644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _03933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _03258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _21926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _27065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _03959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _27066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _27067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _27068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _27069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _27070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _13781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _14645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _17209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _03970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _11687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _27040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _25931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _05581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _27041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _25947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _05579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _05748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _25919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _06145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _26997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _09947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _10008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _26998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _26999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _05915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _09069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _08989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _27000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _09159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _09155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _06291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _08777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _08772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _06297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _08696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _07414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _06173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _06087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _02461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _26995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _26996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _02648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _06199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _26972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _26649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _06206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _26973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _06072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _12649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _07416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _10162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _10172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _10193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _08927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _09731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _27315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _27316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _09051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _01367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _01354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _10718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _27265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _02641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _10710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _01070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _01116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _27255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _27256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _27257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _27258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _10592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _27259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _10630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _27260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _11300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _11380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _11305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _07355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _07816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _10815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _10872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _10835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _22729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _01215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _22695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _22652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _19697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _18556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _14741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _07364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _12164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _12480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _12457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _12434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _10554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _11035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _27254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _11043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _27251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _22632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _27252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _27253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _07080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _07362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _12162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _12172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _04117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _04791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _04137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _06722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _06592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _10268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _02085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _02068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _01407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _23957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _27249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _10490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _24878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _27250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _25062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _07367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _10348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _03022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _03649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _10328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _25698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _00164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _25912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _10437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _09205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _09202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _10213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _09281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _09251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _07401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _08888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _08787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _09109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _09106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _10219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _27245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _27246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _27247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _08741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _27248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _27125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _10167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _27126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _11957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _04997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _04991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _05053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _05036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _10469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _10354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _10331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _11955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _11143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _11031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _11422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _27111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _11947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _18475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _18678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _11945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _11567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _14596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _14374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _13902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _17026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _16909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _11949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _12030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _11746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _12299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _27095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _27096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _22653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _27037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _22624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _22623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _27038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _22628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _22627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _22626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _22697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _27088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _27089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _22664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _09027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _22689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _03786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _03856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _22709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _25768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _25535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _09719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _05716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _04120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _18789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _27084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _11226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _27085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _08939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _22625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _27086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _03011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _27087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _04176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _23201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _27083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _03146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _23048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _03851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _03845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _03268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _24231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _26425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _00681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _00592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _00511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _04099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _03230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _27080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _23905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _27082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _03807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _23400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _03771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _23272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _23343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _23336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _03818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _03739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _03765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _23708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _03153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _23970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _27081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _24066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _24060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _04053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _01193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _01413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _04090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _27078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _02051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _04084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _27079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _04047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _27072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _27073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _03045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _27074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _27075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _27076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _27077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _07957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _07729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _04038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _08829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _09285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _04029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _03240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _27071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _22659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _22654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _22656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _22662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _22660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _27064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _22631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _22630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _04008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _12238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _03995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _03252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _10243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _04024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _10904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _03049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _25480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _27060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _22882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _27061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _03129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _27062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _22755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _03873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _27063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _22699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _22741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _22737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _03906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _22667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _22693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _22692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _05366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _05711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _03036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _27058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _27059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _03060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _03071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _05340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _02965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _27055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _27056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _02999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _27057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _05383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _03020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _05370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _05422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _02907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _27052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _27053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _05406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _02946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _27054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _02952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _05467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _01566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _27043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _27044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _05722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _27045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _27046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _27047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _27048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _27049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _05432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _27050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _27051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _05429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _02846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _05629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _05491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _00162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _05652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _00460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _01494_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _05476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _01500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _05472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _05527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _05742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _26012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _27035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _27036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _26043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _05520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _26808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _00134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _05506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _00139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _05658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _27042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _00157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _05494_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _05729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _27039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _05516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _00071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _05664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _00077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _00085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _05512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _05737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _25969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _05540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _05745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _25982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _25992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _05535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _25998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _05531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _06914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _06892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _27033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _06890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _25951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _25954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _05572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _27034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _03243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _06498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _25894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _25884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _03131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _03123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _03108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _27032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _03333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _27030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _03401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _03377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _05818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _03200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _03172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _27031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _01758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _24455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _05841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _27194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _05844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _01779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _27195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _27196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _05828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _03502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _03484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _03590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _27029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _03561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _03347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _03342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _03948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _03936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _05830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _03640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _03673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _03668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _03762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _03741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _04275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _27027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _04396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _04380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _06463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _04063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _04058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _04185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _04173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _04127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _06468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _06024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _03813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _27028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _06473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _04490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _04471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _04548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _27026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _04581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _05837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _06096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _04286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _06028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _04697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _04685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _04666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _04738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _04768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _27023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _06453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _05071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _27020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _04806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _27021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _04809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _27022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _04914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _04903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _05672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _05667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _06400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _05734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _05725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _27016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _27017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _05132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _06405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _27018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _05209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _27019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _06102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _04986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _04982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _05075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _27014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _05859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _05812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _27015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _06392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _05880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _06389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _06039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _06068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _06153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _06141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _05863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _06105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _05995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _05992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _05949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _27013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _06232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _06226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _06372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _06266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _06295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _06272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _05868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _05883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _06109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _06523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _06518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _27010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _27011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _27012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _06584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _05878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _06374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _06365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _06354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _06440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _06447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _06442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _05873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _06830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _06825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _27006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _06657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _27007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _27008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _27009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _06700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _06975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _06966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _27005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _06750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _06771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _06756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _06349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _06819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _07042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _07027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _07114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _07100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _27004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _06904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _06897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _06988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _07514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _05902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _07350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _07345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _07330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _06333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _07418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _27003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _07187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _07178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _07148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _07252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _07247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _07232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _05897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _07020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _07787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _06319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _07823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _07819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _06314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _07460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _07451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _06324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _08923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _05910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _08170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _27001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _08196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _08189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _27002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _06050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _06160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _11235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _26993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _06163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _06091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _06170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _26994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _06167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _10175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _06287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _26987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _10231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _05927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _06119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _26988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _01618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _06263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _26984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _26985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _10507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _06278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _26986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _10813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _10150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _11563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _11574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _11701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _06252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _26978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _11356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _26979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _11485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _06122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _11147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _26980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _11222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _05937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _26981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _26982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _26983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _12169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _12153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _12191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _05969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _11879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _06249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _11941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _05942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _06237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _12604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _26976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _05982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _12423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _12371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _12504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _26977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _06213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _10742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _06219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _26974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _05989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _12160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _11132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _03451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _26975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _05987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _12645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _04760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _01371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _05984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _12559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _12532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _26967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _06928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _26968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _26969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _26970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _26971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _11041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _03953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _26960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _26961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _06956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _26962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _07117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _26963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _26964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _26965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _26957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _06982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _10823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _07125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _26958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _26959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _06973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _07197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _10874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _06970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _10882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _07121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _10888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _10899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _06962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _07195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _06999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _10751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _06994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _10762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _07131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _26955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _10809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _26956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _09818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _09861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _07009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _26954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _10451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _10650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _07004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _10656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _26951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _26952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _26953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _07184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _07239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _09791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _09816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _07013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _06382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _26947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _07333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _07078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _07338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _07173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _07430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _07448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _11083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _22744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _24727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _24419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _11137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _24454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _11139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _24183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _11104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _22629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _26942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _24022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _11703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _24790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _26943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _26944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _26929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _10546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _10579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _08907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _09122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _10586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _10622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _08904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _00420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _08539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _27243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _07867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _09366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _09341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _27244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _09546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _11159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _24159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _11061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _26939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _11057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _26940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _26941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _11123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _10302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _09067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _10374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _10460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _08914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _09137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _26927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _26928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _08921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _10203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _09076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _10216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _26925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _08917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _09126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _26926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _03190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _27317_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _04628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _02967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _12045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _03197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _04575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _10902_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _27318_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _27319_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _27319_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _27319_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _27319_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _27320_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _27321_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _27322_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _27322_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _27322_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _27322_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _27322_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _27322_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _27322_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _27322_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10511_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10500_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10414_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10380_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10177_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _06433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _06437_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _06435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _06450_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _06459_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _06456_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _06465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _09941_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _09939_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _09907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _09892_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _09879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _09740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _09981_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _09762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09776_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _09932_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _09854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _09806_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _09937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _09935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _09852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _09950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _11650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _22647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _09078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _09242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _09188_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _09132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _09104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _11732_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _08562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _11447_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _11586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _08453_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _22649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _11534_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _08759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _22648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _11529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _08082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _11558_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _11460_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _11550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _11510_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _07624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _07604_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _07585_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _11523_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _07060_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _06907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _07039_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _07003_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _06955_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _22650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _07403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _11597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _06545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _06526_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _06503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _06483_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _22651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _06761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _06717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _11561_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _11382_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _11355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _11331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _05905_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _11811_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _11654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _11786_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _10963_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _10447_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _10424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _10401_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _10378_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _05929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _10980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _10777_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _10945_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _09994_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _09827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _09956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _09928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _09902_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _09875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _05998_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _10802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _09390_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _09369_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _09347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _09305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _06005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _09650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _09507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _10929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10185_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _09841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _06619_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _06900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _06894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _06911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _06908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _06909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _06918_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _06916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _06641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _03784_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _03390_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _04087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _05233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _04648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _04060_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _06116_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _10977_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _10001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _01918_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _04094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _06060_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _24831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _02094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _08256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _22691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _22677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _22702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _11603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _08935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12614_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _04110_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _12647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _12643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _06385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12568_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _04133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _12598_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _12596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _12594_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _12591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _25345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _06553_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12546_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12541_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _04135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _02153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _24756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _01337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _04534_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _04320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _22641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _22637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _22636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _22634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _07470_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _07467_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _07465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _03788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _07411_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _07409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _25886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02944_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _03815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _07360_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _07339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _07358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _07352_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _07347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _22633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _07327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _07325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _07323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _07320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _07316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _07314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _07249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _07277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _07275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _07273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _07255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02992_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _18587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _07206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _07219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _07217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _07213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _07211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _07208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _03002_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01259_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _22894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _22904_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _22901_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _22898_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _22747_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _22766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _22734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _22735_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _22736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _22751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _01186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _25649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _25645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _01269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _25686_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _25684_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _22757_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _01265_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _22752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _22754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _22819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _01184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _22639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _22640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _22851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _22638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _22879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _22831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _22859_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _01202_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _25563_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _25557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _25560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _01279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _22756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _22758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _22759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _25626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _22733_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _22732_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _22731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _22730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _22728_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _22727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _22726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _22725_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22724_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _25624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _22722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _22721_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _22635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _22720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _11753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _22719_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _22718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _22717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _22716_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _22715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _22714_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _22713_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _22712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _22711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01176_);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
