
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire [7:0] acc;
  input clk;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_pc;
  wire [7:0] psw;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [7:0] \uc8051golden_1.ACC ;
  wire [7:0] \uc8051golden_1.ACC_03 ;
  wire [7:0] \uc8051golden_1.ACC_13 ;
  wire [7:0] \uc8051golden_1.ACC_23 ;
  wire [7:0] \uc8051golden_1.ACC_33 ;
  wire [7:0] \uc8051golden_1.ACC_c4 ;
  wire [7:0] \uc8051golden_1.ACC_c6 ;
  wire [7:0] \uc8051golden_1.ACC_c7 ;
  wire [7:0] \uc8051golden_1.ACC_d6 ;
  wire [7:0] \uc8051golden_1.ACC_d7 ;
  wire [7:0] \uc8051golden_1.ACC_e6 ;
  wire [7:0] \uc8051golden_1.ACC_e7 ;
  wire [7:0] \uc8051golden_1.B ;
  wire [7:0] \uc8051golden_1.DPH ;
  wire [7:0] \uc8051golden_1.DPL ;
  wire [7:0] \uc8051golden_1.IE ;
  wire [7:0] \uc8051golden_1.IP ;
  wire [7:0] \uc8051golden_1.IRAM[0] ;
  wire [7:0] \uc8051golden_1.IRAM[100] ;
  wire [7:0] \uc8051golden_1.IRAM[101] ;
  wire [7:0] \uc8051golden_1.IRAM[102] ;
  wire [7:0] \uc8051golden_1.IRAM[103] ;
  wire [7:0] \uc8051golden_1.IRAM[104] ;
  wire [7:0] \uc8051golden_1.IRAM[105] ;
  wire [7:0] \uc8051golden_1.IRAM[106] ;
  wire [7:0] \uc8051golden_1.IRAM[107] ;
  wire [7:0] \uc8051golden_1.IRAM[108] ;
  wire [7:0] \uc8051golden_1.IRAM[109] ;
  wire [7:0] \uc8051golden_1.IRAM[10] ;
  wire [7:0] \uc8051golden_1.IRAM[110] ;
  wire [7:0] \uc8051golden_1.IRAM[111] ;
  wire [7:0] \uc8051golden_1.IRAM[112] ;
  wire [7:0] \uc8051golden_1.IRAM[113] ;
  wire [7:0] \uc8051golden_1.IRAM[114] ;
  wire [7:0] \uc8051golden_1.IRAM[115] ;
  wire [7:0] \uc8051golden_1.IRAM[116] ;
  wire [7:0] \uc8051golden_1.IRAM[117] ;
  wire [7:0] \uc8051golden_1.IRAM[118] ;
  wire [7:0] \uc8051golden_1.IRAM[119] ;
  wire [7:0] \uc8051golden_1.IRAM[11] ;
  wire [7:0] \uc8051golden_1.IRAM[120] ;
  wire [7:0] \uc8051golden_1.IRAM[121] ;
  wire [7:0] \uc8051golden_1.IRAM[122] ;
  wire [7:0] \uc8051golden_1.IRAM[123] ;
  wire [7:0] \uc8051golden_1.IRAM[124] ;
  wire [7:0] \uc8051golden_1.IRAM[125] ;
  wire [7:0] \uc8051golden_1.IRAM[126] ;
  wire [7:0] \uc8051golden_1.IRAM[127] ;
  wire [7:0] \uc8051golden_1.IRAM[128] ;
  wire [7:0] \uc8051golden_1.IRAM[129] ;
  wire [7:0] \uc8051golden_1.IRAM[12] ;
  wire [7:0] \uc8051golden_1.IRAM[130] ;
  wire [7:0] \uc8051golden_1.IRAM[131] ;
  wire [7:0] \uc8051golden_1.IRAM[132] ;
  wire [7:0] \uc8051golden_1.IRAM[133] ;
  wire [7:0] \uc8051golden_1.IRAM[134] ;
  wire [7:0] \uc8051golden_1.IRAM[135] ;
  wire [7:0] \uc8051golden_1.IRAM[136] ;
  wire [7:0] \uc8051golden_1.IRAM[137] ;
  wire [7:0] \uc8051golden_1.IRAM[138] ;
  wire [7:0] \uc8051golden_1.IRAM[139] ;
  wire [7:0] \uc8051golden_1.IRAM[13] ;
  wire [7:0] \uc8051golden_1.IRAM[140] ;
  wire [7:0] \uc8051golden_1.IRAM[141] ;
  wire [7:0] \uc8051golden_1.IRAM[142] ;
  wire [7:0] \uc8051golden_1.IRAM[143] ;
  wire [7:0] \uc8051golden_1.IRAM[144] ;
  wire [7:0] \uc8051golden_1.IRAM[145] ;
  wire [7:0] \uc8051golden_1.IRAM[146] ;
  wire [7:0] \uc8051golden_1.IRAM[147] ;
  wire [7:0] \uc8051golden_1.IRAM[148] ;
  wire [7:0] \uc8051golden_1.IRAM[149] ;
  wire [7:0] \uc8051golden_1.IRAM[14] ;
  wire [7:0] \uc8051golden_1.IRAM[150] ;
  wire [7:0] \uc8051golden_1.IRAM[151] ;
  wire [7:0] \uc8051golden_1.IRAM[152] ;
  wire [7:0] \uc8051golden_1.IRAM[153] ;
  wire [7:0] \uc8051golden_1.IRAM[154] ;
  wire [7:0] \uc8051golden_1.IRAM[155] ;
  wire [7:0] \uc8051golden_1.IRAM[156] ;
  wire [7:0] \uc8051golden_1.IRAM[157] ;
  wire [7:0] \uc8051golden_1.IRAM[158] ;
  wire [7:0] \uc8051golden_1.IRAM[159] ;
  wire [7:0] \uc8051golden_1.IRAM[15] ;
  wire [7:0] \uc8051golden_1.IRAM[160] ;
  wire [7:0] \uc8051golden_1.IRAM[161] ;
  wire [7:0] \uc8051golden_1.IRAM[162] ;
  wire [7:0] \uc8051golden_1.IRAM[163] ;
  wire [7:0] \uc8051golden_1.IRAM[164] ;
  wire [7:0] \uc8051golden_1.IRAM[165] ;
  wire [7:0] \uc8051golden_1.IRAM[166] ;
  wire [7:0] \uc8051golden_1.IRAM[167] ;
  wire [7:0] \uc8051golden_1.IRAM[168] ;
  wire [7:0] \uc8051golden_1.IRAM[169] ;
  wire [7:0] \uc8051golden_1.IRAM[16] ;
  wire [7:0] \uc8051golden_1.IRAM[170] ;
  wire [7:0] \uc8051golden_1.IRAM[171] ;
  wire [7:0] \uc8051golden_1.IRAM[172] ;
  wire [7:0] \uc8051golden_1.IRAM[173] ;
  wire [7:0] \uc8051golden_1.IRAM[174] ;
  wire [7:0] \uc8051golden_1.IRAM[175] ;
  wire [7:0] \uc8051golden_1.IRAM[176] ;
  wire [7:0] \uc8051golden_1.IRAM[177] ;
  wire [7:0] \uc8051golden_1.IRAM[178] ;
  wire [7:0] \uc8051golden_1.IRAM[179] ;
  wire [7:0] \uc8051golden_1.IRAM[17] ;
  wire [7:0] \uc8051golden_1.IRAM[180] ;
  wire [7:0] \uc8051golden_1.IRAM[181] ;
  wire [7:0] \uc8051golden_1.IRAM[182] ;
  wire [7:0] \uc8051golden_1.IRAM[183] ;
  wire [7:0] \uc8051golden_1.IRAM[184] ;
  wire [7:0] \uc8051golden_1.IRAM[185] ;
  wire [7:0] \uc8051golden_1.IRAM[186] ;
  wire [7:0] \uc8051golden_1.IRAM[187] ;
  wire [7:0] \uc8051golden_1.IRAM[188] ;
  wire [7:0] \uc8051golden_1.IRAM[189] ;
  wire [7:0] \uc8051golden_1.IRAM[18] ;
  wire [7:0] \uc8051golden_1.IRAM[190] ;
  wire [7:0] \uc8051golden_1.IRAM[191] ;
  wire [7:0] \uc8051golden_1.IRAM[192] ;
  wire [7:0] \uc8051golden_1.IRAM[193] ;
  wire [7:0] \uc8051golden_1.IRAM[194] ;
  wire [7:0] \uc8051golden_1.IRAM[195] ;
  wire [7:0] \uc8051golden_1.IRAM[196] ;
  wire [7:0] \uc8051golden_1.IRAM[197] ;
  wire [7:0] \uc8051golden_1.IRAM[198] ;
  wire [7:0] \uc8051golden_1.IRAM[199] ;
  wire [7:0] \uc8051golden_1.IRAM[19] ;
  wire [7:0] \uc8051golden_1.IRAM[1] ;
  wire [7:0] \uc8051golden_1.IRAM[200] ;
  wire [7:0] \uc8051golden_1.IRAM[201] ;
  wire [7:0] \uc8051golden_1.IRAM[202] ;
  wire [7:0] \uc8051golden_1.IRAM[203] ;
  wire [7:0] \uc8051golden_1.IRAM[204] ;
  wire [7:0] \uc8051golden_1.IRAM[205] ;
  wire [7:0] \uc8051golden_1.IRAM[206] ;
  wire [7:0] \uc8051golden_1.IRAM[207] ;
  wire [7:0] \uc8051golden_1.IRAM[208] ;
  wire [7:0] \uc8051golden_1.IRAM[209] ;
  wire [7:0] \uc8051golden_1.IRAM[20] ;
  wire [7:0] \uc8051golden_1.IRAM[210] ;
  wire [7:0] \uc8051golden_1.IRAM[211] ;
  wire [7:0] \uc8051golden_1.IRAM[212] ;
  wire [7:0] \uc8051golden_1.IRAM[213] ;
  wire [7:0] \uc8051golden_1.IRAM[214] ;
  wire [7:0] \uc8051golden_1.IRAM[215] ;
  wire [7:0] \uc8051golden_1.IRAM[216] ;
  wire [7:0] \uc8051golden_1.IRAM[217] ;
  wire [7:0] \uc8051golden_1.IRAM[218] ;
  wire [7:0] \uc8051golden_1.IRAM[219] ;
  wire [7:0] \uc8051golden_1.IRAM[21] ;
  wire [7:0] \uc8051golden_1.IRAM[220] ;
  wire [7:0] \uc8051golden_1.IRAM[221] ;
  wire [7:0] \uc8051golden_1.IRAM[222] ;
  wire [7:0] \uc8051golden_1.IRAM[223] ;
  wire [7:0] \uc8051golden_1.IRAM[224] ;
  wire [7:0] \uc8051golden_1.IRAM[225] ;
  wire [7:0] \uc8051golden_1.IRAM[226] ;
  wire [7:0] \uc8051golden_1.IRAM[227] ;
  wire [7:0] \uc8051golden_1.IRAM[228] ;
  wire [7:0] \uc8051golden_1.IRAM[229] ;
  wire [7:0] \uc8051golden_1.IRAM[22] ;
  wire [7:0] \uc8051golden_1.IRAM[230] ;
  wire [7:0] \uc8051golden_1.IRAM[231] ;
  wire [7:0] \uc8051golden_1.IRAM[232] ;
  wire [7:0] \uc8051golden_1.IRAM[233] ;
  wire [7:0] \uc8051golden_1.IRAM[234] ;
  wire [7:0] \uc8051golden_1.IRAM[235] ;
  wire [7:0] \uc8051golden_1.IRAM[236] ;
  wire [7:0] \uc8051golden_1.IRAM[237] ;
  wire [7:0] \uc8051golden_1.IRAM[238] ;
  wire [7:0] \uc8051golden_1.IRAM[239] ;
  wire [7:0] \uc8051golden_1.IRAM[23] ;
  wire [7:0] \uc8051golden_1.IRAM[240] ;
  wire [7:0] \uc8051golden_1.IRAM[241] ;
  wire [7:0] \uc8051golden_1.IRAM[242] ;
  wire [7:0] \uc8051golden_1.IRAM[243] ;
  wire [7:0] \uc8051golden_1.IRAM[244] ;
  wire [7:0] \uc8051golden_1.IRAM[245] ;
  wire [7:0] \uc8051golden_1.IRAM[246] ;
  wire [7:0] \uc8051golden_1.IRAM[247] ;
  wire [7:0] \uc8051golden_1.IRAM[248] ;
  wire [7:0] \uc8051golden_1.IRAM[249] ;
  wire [7:0] \uc8051golden_1.IRAM[24] ;
  wire [7:0] \uc8051golden_1.IRAM[250] ;
  wire [7:0] \uc8051golden_1.IRAM[251] ;
  wire [7:0] \uc8051golden_1.IRAM[252] ;
  wire [7:0] \uc8051golden_1.IRAM[253] ;
  wire [7:0] \uc8051golden_1.IRAM[254] ;
  wire [7:0] \uc8051golden_1.IRAM[255] ;
  wire [7:0] \uc8051golden_1.IRAM[25] ;
  wire [7:0] \uc8051golden_1.IRAM[26] ;
  wire [7:0] \uc8051golden_1.IRAM[27] ;
  wire [7:0] \uc8051golden_1.IRAM[28] ;
  wire [7:0] \uc8051golden_1.IRAM[29] ;
  wire [7:0] \uc8051golden_1.IRAM[2] ;
  wire [7:0] \uc8051golden_1.IRAM[30] ;
  wire [7:0] \uc8051golden_1.IRAM[31] ;
  wire [7:0] \uc8051golden_1.IRAM[32] ;
  wire [7:0] \uc8051golden_1.IRAM[33] ;
  wire [7:0] \uc8051golden_1.IRAM[34] ;
  wire [7:0] \uc8051golden_1.IRAM[35] ;
  wire [7:0] \uc8051golden_1.IRAM[36] ;
  wire [7:0] \uc8051golden_1.IRAM[37] ;
  wire [7:0] \uc8051golden_1.IRAM[38] ;
  wire [7:0] \uc8051golden_1.IRAM[39] ;
  wire [7:0] \uc8051golden_1.IRAM[3] ;
  wire [7:0] \uc8051golden_1.IRAM[40] ;
  wire [7:0] \uc8051golden_1.IRAM[41] ;
  wire [7:0] \uc8051golden_1.IRAM[42] ;
  wire [7:0] \uc8051golden_1.IRAM[43] ;
  wire [7:0] \uc8051golden_1.IRAM[44] ;
  wire [7:0] \uc8051golden_1.IRAM[45] ;
  wire [7:0] \uc8051golden_1.IRAM[46] ;
  wire [7:0] \uc8051golden_1.IRAM[47] ;
  wire [7:0] \uc8051golden_1.IRAM[48] ;
  wire [7:0] \uc8051golden_1.IRAM[49] ;
  wire [7:0] \uc8051golden_1.IRAM[4] ;
  wire [7:0] \uc8051golden_1.IRAM[50] ;
  wire [7:0] \uc8051golden_1.IRAM[51] ;
  wire [7:0] \uc8051golden_1.IRAM[52] ;
  wire [7:0] \uc8051golden_1.IRAM[53] ;
  wire [7:0] \uc8051golden_1.IRAM[54] ;
  wire [7:0] \uc8051golden_1.IRAM[55] ;
  wire [7:0] \uc8051golden_1.IRAM[56] ;
  wire [7:0] \uc8051golden_1.IRAM[57] ;
  wire [7:0] \uc8051golden_1.IRAM[58] ;
  wire [7:0] \uc8051golden_1.IRAM[59] ;
  wire [7:0] \uc8051golden_1.IRAM[5] ;
  wire [7:0] \uc8051golden_1.IRAM[60] ;
  wire [7:0] \uc8051golden_1.IRAM[61] ;
  wire [7:0] \uc8051golden_1.IRAM[62] ;
  wire [7:0] \uc8051golden_1.IRAM[63] ;
  wire [7:0] \uc8051golden_1.IRAM[64] ;
  wire [7:0] \uc8051golden_1.IRAM[65] ;
  wire [7:0] \uc8051golden_1.IRAM[66] ;
  wire [7:0] \uc8051golden_1.IRAM[67] ;
  wire [7:0] \uc8051golden_1.IRAM[68] ;
  wire [7:0] \uc8051golden_1.IRAM[69] ;
  wire [7:0] \uc8051golden_1.IRAM[6] ;
  wire [7:0] \uc8051golden_1.IRAM[70] ;
  wire [7:0] \uc8051golden_1.IRAM[71] ;
  wire [7:0] \uc8051golden_1.IRAM[72] ;
  wire [7:0] \uc8051golden_1.IRAM[73] ;
  wire [7:0] \uc8051golden_1.IRAM[74] ;
  wire [7:0] \uc8051golden_1.IRAM[75] ;
  wire [7:0] \uc8051golden_1.IRAM[76] ;
  wire [7:0] \uc8051golden_1.IRAM[77] ;
  wire [7:0] \uc8051golden_1.IRAM[78] ;
  wire [7:0] \uc8051golden_1.IRAM[79] ;
  wire [7:0] \uc8051golden_1.IRAM[7] ;
  wire [7:0] \uc8051golden_1.IRAM[80] ;
  wire [7:0] \uc8051golden_1.IRAM[81] ;
  wire [7:0] \uc8051golden_1.IRAM[82] ;
  wire [7:0] \uc8051golden_1.IRAM[83] ;
  wire [7:0] \uc8051golden_1.IRAM[84] ;
  wire [7:0] \uc8051golden_1.IRAM[85] ;
  wire [7:0] \uc8051golden_1.IRAM[86] ;
  wire [7:0] \uc8051golden_1.IRAM[87] ;
  wire [7:0] \uc8051golden_1.IRAM[88] ;
  wire [7:0] \uc8051golden_1.IRAM[89] ;
  wire [7:0] \uc8051golden_1.IRAM[8] ;
  wire [7:0] \uc8051golden_1.IRAM[90] ;
  wire [7:0] \uc8051golden_1.IRAM[91] ;
  wire [7:0] \uc8051golden_1.IRAM[92] ;
  wire [7:0] \uc8051golden_1.IRAM[93] ;
  wire [7:0] \uc8051golden_1.IRAM[94] ;
  wire [7:0] \uc8051golden_1.IRAM[95] ;
  wire [7:0] \uc8051golden_1.IRAM[96] ;
  wire [7:0] \uc8051golden_1.IRAM[97] ;
  wire [7:0] \uc8051golden_1.IRAM[98] ;
  wire [7:0] \uc8051golden_1.IRAM[99] ;
  wire [7:0] \uc8051golden_1.IRAM[9] ;
  wire [7:0] \uc8051golden_1.P0 ;
  wire [7:0] \uc8051golden_1.P1 ;
  wire [7:0] \uc8051golden_1.P2 ;
  wire [7:0] \uc8051golden_1.P3 ;
  wire [15:0] \uc8051golden_1.PC ;
  wire [7:0] \uc8051golden_1.PCON ;
  wire [7:0] \uc8051golden_1.PSW ;
  wire [7:0] \uc8051golden_1.PSW_0d ;
  wire [7:0] \uc8051golden_1.PSW_13 ;
  wire [7:0] \uc8051golden_1.PSW_24 ;
  wire [7:0] \uc8051golden_1.PSW_25 ;
  wire [7:0] \uc8051golden_1.PSW_26 ;
  wire [7:0] \uc8051golden_1.PSW_27 ;
  wire [7:0] \uc8051golden_1.PSW_28 ;
  wire [7:0] \uc8051golden_1.PSW_29 ;
  wire [7:0] \uc8051golden_1.PSW_2a ;
  wire [7:0] \uc8051golden_1.PSW_2b ;
  wire [7:0] \uc8051golden_1.PSW_2c ;
  wire [7:0] \uc8051golden_1.PSW_2d ;
  wire [7:0] \uc8051golden_1.PSW_2e ;
  wire [7:0] \uc8051golden_1.PSW_2f ;
  wire [7:0] \uc8051golden_1.PSW_33 ;
  wire [7:0] \uc8051golden_1.PSW_34 ;
  wire [7:0] \uc8051golden_1.PSW_35 ;
  wire [7:0] \uc8051golden_1.PSW_36 ;
  wire [7:0] \uc8051golden_1.PSW_37 ;
  wire [7:0] \uc8051golden_1.PSW_38 ;
  wire [7:0] \uc8051golden_1.PSW_39 ;
  wire [7:0] \uc8051golden_1.PSW_3a ;
  wire [7:0] \uc8051golden_1.PSW_3b ;
  wire [7:0] \uc8051golden_1.PSW_3c ;
  wire [7:0] \uc8051golden_1.PSW_3d ;
  wire [7:0] \uc8051golden_1.PSW_3e ;
  wire [7:0] \uc8051golden_1.PSW_3f ;
  wire [7:0] \uc8051golden_1.PSW_46 ;
  wire [7:0] \uc8051golden_1.PSW_65 ;
  wire [7:0] \uc8051golden_1.PSW_72 ;
  wire [7:0] \uc8051golden_1.PSW_82 ;
  wire [7:0] \uc8051golden_1.PSW_84 ;
  wire [7:0] \uc8051golden_1.PSW_94 ;
  wire [7:0] \uc8051golden_1.PSW_95 ;
  wire [7:0] \uc8051golden_1.PSW_96 ;
  wire [7:0] \uc8051golden_1.PSW_97 ;
  wire [7:0] \uc8051golden_1.PSW_98 ;
  wire [7:0] \uc8051golden_1.PSW_99 ;
  wire [7:0] \uc8051golden_1.PSW_9a ;
  wire [7:0] \uc8051golden_1.PSW_9b ;
  wire [7:0] \uc8051golden_1.PSW_9c ;
  wire [7:0] \uc8051golden_1.PSW_9d ;
  wire [7:0] \uc8051golden_1.PSW_9e ;
  wire [7:0] \uc8051golden_1.PSW_9f ;
  wire [7:0] \uc8051golden_1.PSW_a0 ;
  wire [7:0] \uc8051golden_1.PSW_a2 ;
  wire [7:0] \uc8051golden_1.PSW_a4 ;
  wire [7:0] \uc8051golden_1.PSW_b0 ;
  wire [7:0] \uc8051golden_1.PSW_b3 ;
  wire [7:0] \uc8051golden_1.PSW_b4 ;
  wire [7:0] \uc8051golden_1.PSW_b5 ;
  wire [7:0] \uc8051golden_1.PSW_b6 ;
  wire [7:0] \uc8051golden_1.PSW_b7 ;
  wire [7:0] \uc8051golden_1.PSW_b8 ;
  wire [7:0] \uc8051golden_1.PSW_b9 ;
  wire [7:0] \uc8051golden_1.PSW_ba ;
  wire [7:0] \uc8051golden_1.PSW_bb ;
  wire [7:0] \uc8051golden_1.PSW_bc ;
  wire [7:0] \uc8051golden_1.PSW_bd ;
  wire [7:0] \uc8051golden_1.PSW_be ;
  wire [7:0] \uc8051golden_1.PSW_bf ;
  wire [7:0] \uc8051golden_1.PSW_c0 ;
  wire [7:0] \uc8051golden_1.PSW_c3 ;
  wire [7:0] \uc8051golden_1.PSW_ce ;
  wire [7:0] \uc8051golden_1.PSW_d3 ;
  wire [7:0] \uc8051golden_1.PSW_d4 ;
  wire [7:0] \uc8051golden_1.SBUF ;
  wire [7:0] \uc8051golden_1.SCON ;
  wire [7:0] \uc8051golden_1.SP ;
  wire [7:0] \uc8051golden_1.TCON ;
  wire [7:0] \uc8051golden_1.TH0 ;
  wire [7:0] \uc8051golden_1.TH1 ;
  wire [7:0] \uc8051golden_1.TL0 ;
  wire [7:0] \uc8051golden_1.TL1 ;
  wire [7:0] \uc8051golden_1.TMOD ;
  wire \uc8051golden_1.clk ;
  wire [7:0] \uc8051golden_1.n0014 ;
  wire [1:0] \uc8051golden_1.n0109 ;
  wire [7:0] \uc8051golden_1.n0110 ;
  wire [7:0] \uc8051golden_1.n0112 ;
  wire [7:0] \uc8051golden_1.n0115 ;
  wire [7:0] \uc8051golden_1.n0117 ;
  wire [7:0] \uc8051golden_1.n0124 ;
  wire [7:0] \uc8051golden_1.n0128 ;
  wire [7:0] \uc8051golden_1.n0132 ;
  wire [7:0] \uc8051golden_1.n0136 ;
  wire \uc8051golden_1.n0139 ;
  wire \uc8051golden_1.n0140 ;
  wire [2:0] \uc8051golden_1.n0141 ;
  wire \uc8051golden_1.n0142 ;
  wire [1:0] \uc8051golden_1.n0143 ;
  wire [7:0] \uc8051golden_1.n0144 ;
  wire [7:0] \uc8051golden_1.n0146 ;
  wire [7:0] \uc8051golden_1.n0150 ;
  wire [8:0] \uc8051golden_1.n0223 ;
  wire [8:0] \uc8051golden_1.n0224 ;
  wire [7:0] \uc8051golden_1.n0225 ;
  wire \uc8051golden_1.n0226 ;
  wire [7:0] \uc8051golden_1.n0227 ;
  wire [7:0] \uc8051golden_1.n0266 ;
  wire [8:0] \uc8051golden_1.n0268 ;
  wire [3:0] \uc8051golden_1.n0274 ;
  wire [4:0] \uc8051golden_1.n0275 ;
  wire [8:0] \uc8051golden_1.n0282 ;
  wire [7:0] \uc8051golden_1.n0291 ;
  wire [7:0] \uc8051golden_1.n0359 ;
  wire [8:0] \uc8051golden_1.n0361 ;
  wire [3:0] \uc8051golden_1.n0365 ;
  wire [4:0] \uc8051golden_1.n0366 ;
  wire [8:0] \uc8051golden_1.n0370 ;
  wire [7:0] \uc8051golden_1.n0378 ;
  wire [8:0] \uc8051golden_1.n0380 ;
  wire [3:0] \uc8051golden_1.n0385 ;
  wire [4:0] \uc8051golden_1.n0386 ;
  wire [8:0] \uc8051golden_1.n0390 ;
  wire [7:0] \uc8051golden_1.n0398 ;
  wire [7:0] \uc8051golden_1.n0417 ;
  wire [7:0] \uc8051golden_1.n0436 ;
  wire [7:0] \uc8051golden_1.n0455 ;
  wire [7:0] \uc8051golden_1.n0474 ;
  wire [7:0] \uc8051golden_1.n0493 ;
  wire [7:0] \uc8051golden_1.n0513 ;
  wire [7:0] \uc8051golden_1.n0532 ;
  wire [7:0] \uc8051golden_1.n0551 ;
  wire [8:0] \uc8051golden_1.n0555 ;
  wire [8:0] \uc8051golden_1.n0556 ;
  wire [7:0] \uc8051golden_1.n0557 ;
  wire \uc8051golden_1.n0558 ;
  wire [7:0] \uc8051golden_1.n0559 ;
  wire [7:0] \uc8051golden_1.n0560 ;
  wire [8:0] \uc8051golden_1.n0563 ;
  wire [4:0] \uc8051golden_1.n0567 ;
  wire [7:0] \uc8051golden_1.n0578 ;
  wire [7:0] \uc8051golden_1.n0594 ;
  wire [7:0] \uc8051golden_1.n0610 ;
  wire [7:0] \uc8051golden_1.n0626 ;
  wire [7:0] \uc8051golden_1.n0642 ;
  wire [7:0] \uc8051golden_1.n0658 ;
  wire [7:0] \uc8051golden_1.n0674 ;
  wire [7:0] \uc8051golden_1.n0690 ;
  wire [7:0] \uc8051golden_1.n0706 ;
  wire [7:0] \uc8051golden_1.n0722 ;
  wire [7:0] \uc8051golden_1.n0738 ;
  wire [7:0] \uc8051golden_1.n0754 ;
  wire [6:0] \uc8051golden_1.n0934 ;
  wire [7:0] \uc8051golden_1.n0935 ;
  wire [15:0] \uc8051golden_1.n0936 ;
  wire [15:0] \uc8051golden_1.n0937 ;
  wire [7:0] \uc8051golden_1.n0962 ;
  wire [3:0] \uc8051golden_1.n0971 ;
  wire [7:0] \uc8051golden_1.n0973 ;
  wire [7:0] \uc8051golden_1.n1207 ;
  wire [7:0] \uc8051golden_1.n1223 ;
  wire [7:0] \uc8051golden_1.n1235 ;
  wire [7:0] \uc8051golden_1.n1248 ;
  wire [7:0] \uc8051golden_1.n1261 ;
  wire [7:0] \uc8051golden_1.n1274 ;
  wire [7:0] \uc8051golden_1.n1287 ;
  wire [7:0] \uc8051golden_1.n1300 ;
  wire [7:0] \uc8051golden_1.n1313 ;
  wire [7:0] \uc8051golden_1.n1326 ;
  wire [7:0] \uc8051golden_1.n1339 ;
  wire [7:0] \uc8051golden_1.n1352 ;
  wire [7:0] \uc8051golden_1.n1365 ;
  wire [7:0] \uc8051golden_1.n1378 ;
  wire [7:0] \uc8051golden_1.n1381 ;
  wire [7:0] \uc8051golden_1.n1382 ;
  wire [15:0] \uc8051golden_1.n1386 ;
  wire [7:0] \uc8051golden_1.n1393 ;
  wire [7:0] \uc8051golden_1.n1395 ;
  wire [7:0] \uc8051golden_1.n1411 ;
  wire [7:0] \uc8051golden_1.n1417 ;
  wire [7:0] \uc8051golden_1.n1423 ;
  wire [7:0] \uc8051golden_1.n1429 ;
  wire [7:0] \uc8051golden_1.n1436 ;
  wire [7:0] \uc8051golden_1.n1442 ;
  wire [7:0] \uc8051golden_1.n1448 ;
  wire [7:0] \uc8051golden_1.n1454 ;
  wire [7:0] \uc8051golden_1.n1460 ;
  wire [7:0] \uc8051golden_1.n1466 ;
  wire [7:0] \uc8051golden_1.n1473 ;
  wire [7:0] \uc8051golden_1.n1479 ;
  wire [7:0] \uc8051golden_1.n1485 ;
  wire [7:0] \uc8051golden_1.n1486 ;
  wire [3:0] \uc8051golden_1.n1487 ;
  wire [7:0] \uc8051golden_1.n1488 ;
  wire [7:0] \uc8051golden_1.n1544 ;
  wire [7:0] \uc8051golden_1.n1564 ;
  wire [7:0] \uc8051golden_1.n1568 ;
  wire [3:0] \uc8051golden_1.n1569 ;
  wire [7:0] \uc8051golden_1.n1570 ;
  wire [7:0] \uc8051golden_1.n1571 ;
  wire [3:0] \uc8051golden_1.n1572 ;
  wire [7:0] \uc8051golden_1.n1573 ;
  wire \uc8051golden_1.rst ;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [31:0] word_in;
  not _25368_ (_00000_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _25369_ (_00001_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _00000_);
  and _25370_ (_00002_, _00001_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _25371_ (_00003_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _00000_);
  and _25372_ (_00004_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _00000_);
  nor _25373_ (_00005_, _00004_, _00003_);
  and _25374_ (_00006_, _00005_, _00002_);
  not _25375_ (_00007_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _25376_ (_00008_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _00007_);
  not _25377_ (_00009_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _25378_ (_00011_, _00009_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nor _25379_ (_00013_, _00011_, _00008_);
  nand _25380_ (_00015_, _00013_, _00006_);
  not _25381_ (_25365_, rst);
  or _25382_ (_00018_, _00006_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _25383_ (_00020_, _00018_, _25365_);
  and _25384_ (_25272_, _00020_, _00015_);
  nor _25385_ (_00023_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _25386_ (_00025_, _00023_);
  and _25387_ (_00027_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _25388_ (_00029_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _25389_ (_00031_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _25390_ (_00033_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _25391_ (_00035_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _25392_ (_00037_, _00035_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _25393_ (_00039_, _00037_, _00033_);
  nor _25394_ (_00041_, _00039_, _00031_);
  nor _25395_ (_00043_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _25396_ (_00045_, _00043_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _25397_ (_00047_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _25398_ (_00049_, _00047_, _00041_);
  nor _25399_ (_00051_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _25400_ (_00053_, _00051_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _25401_ (_00055_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or _25402_ (_00057_, _00037_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _25403_ (_00059_, _00057_);
  and _25404_ (_00061_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _25405_ (_00063_, _00061_, _00055_);
  and _25406_ (_00065_, _00063_, _00049_);
  not _25407_ (_00067_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _25408_ (_00069_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _00067_);
  or _25409_ (_00070_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  not _25410_ (_00071_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _25411_ (_00072_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _00071_);
  and _25412_ (_00073_, _00072_, _00070_);
  or _25413_ (_00074_, _00073_, _00069_);
  nand _25414_ (_00075_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _00067_);
  or _25415_ (_00076_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _25416_ (_00077_, _00076_, _00074_);
  nand _25417_ (_00078_, _00051_, _00035_);
  or _25418_ (_00079_, _00078_, _00077_);
  and _25419_ (_00080_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _25420_ (_00081_, _00080_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _25421_ (_00082_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and _25422_ (_00083_, _00080_, _00033_);
  and _25423_ (_00084_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _25424_ (_00085_, _00084_, _00082_);
  and _25425_ (_00086_, _00085_, _00079_);
  and _25426_ (_00087_, _00086_, _00065_);
  not _25427_ (_00088_, _00087_);
  or _25428_ (_00089_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or _25429_ (_00090_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or _25430_ (_00091_, _00071_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and _25431_ (_00092_, _00091_, _00090_);
  or _25432_ (_00093_, _00092_, _00069_);
  or _25433_ (_00094_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _25434_ (_00095_, _00094_, _00093_);
  or _25435_ (_00096_, _00095_, _00089_);
  and _25436_ (_00097_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _25437_ (_00098_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not _25438_ (_00099_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _25439_ (_00100_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _25440_ (_00101_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _00100_);
  nor _25441_ (_00102_, _00101_, _00099_);
  nor _25442_ (_00103_, _00102_, _00098_);
  and _25443_ (_00104_, _00103_, _00096_);
  nand _25444_ (_00105_, _00104_, _00023_);
  not _25445_ (_00106_, _00008_);
  or _25446_ (_00107_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or _25447_ (_00108_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _00071_);
  and _25448_ (_00109_, _00108_, _00107_);
  or _25449_ (_00110_, _00109_, _00069_);
  or _25450_ (_00111_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _25451_ (_00112_, _00111_, _00110_);
  or _25452_ (_00113_, _00112_, _00089_);
  nand _25453_ (_00114_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not _25454_ (_00115_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _25455_ (_00116_, _00101_, _00115_);
  and _25456_ (_00117_, _00116_, _00114_);
  and _25457_ (_00118_, _00117_, _00113_);
  or _25458_ (_00119_, _00118_, _00106_);
  not _25459_ (_00120_, _00011_);
  or _25460_ (_00121_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or _25461_ (_00122_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _00071_);
  and _25462_ (_00123_, _00122_, _00121_);
  or _25463_ (_00124_, _00123_, _00069_);
  or _25464_ (_00125_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _25465_ (_00126_, _00125_, _00124_);
  or _25466_ (_00127_, _00126_, _00089_);
  nand _25467_ (_00128_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not _25468_ (_00129_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _25469_ (_00130_, _00101_, _00129_);
  and _25470_ (_00131_, _00130_, _00128_);
  and _25471_ (_00132_, _00131_, _00127_);
  or _25472_ (_00133_, _00132_, _00120_);
  and _25473_ (_00134_, _00133_, _00119_);
  or _25474_ (_00135_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or _25475_ (_00136_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _00071_);
  and _25476_ (_00137_, _00136_, _00135_);
  or _25477_ (_00138_, _00137_, _00069_);
  or _25478_ (_00139_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _25479_ (_00140_, _00139_, _00138_);
  or _25480_ (_00141_, _00140_, _00089_);
  nand _25481_ (_00142_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not _25482_ (_00143_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _25483_ (_00144_, _00101_, _00143_);
  and _25484_ (_00145_, _00144_, _00142_);
  nand _25485_ (_00146_, _00145_, _00141_);
  or _25486_ (_00147_, _00146_, _00007_);
  nand _25487_ (_00148_, _00147_, _00013_);
  nand _25488_ (_00149_, _00148_, _00134_);
  and _25489_ (_00150_, _00149_, _00105_);
  and _25490_ (_00151_, _00150_, _00088_);
  or _25491_ (_00152_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or _25492_ (_00153_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _00071_);
  and _25493_ (_00154_, _00153_, _00152_);
  or _25494_ (_00155_, _00154_, _00069_);
  or _25495_ (_00156_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _25496_ (_00157_, _00156_, _00155_);
  or _25497_ (_00158_, _00157_, _00089_);
  and _25498_ (_00159_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not _25499_ (_00160_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _25500_ (_00161_, _00101_, _00160_);
  nor _25501_ (_00162_, _00161_, _00159_);
  and _25502_ (_00163_, _00162_, _00158_);
  nand _25503_ (_00164_, _00163_, _00023_);
  or _25504_ (_00165_, _00077_, _00089_);
  nand _25505_ (_00166_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not _25506_ (_00167_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _25507_ (_00168_, _00101_, _00167_);
  and _25508_ (_00169_, _00168_, _00166_);
  and _25509_ (_00170_, _00169_, _00165_);
  or _25510_ (_00171_, _00170_, _00106_);
  or _25511_ (_00172_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or _25512_ (_00173_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _00071_);
  and _25513_ (_00174_, _00173_, _00172_);
  or _25514_ (_00175_, _00174_, _00069_);
  or _25515_ (_00176_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _25516_ (_00177_, _00176_, _00175_);
  or _25517_ (_00178_, _00177_, _00089_);
  nand _25518_ (_00179_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _25519_ (_00180_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _25520_ (_00181_, _00101_, _00180_);
  and _25521_ (_00182_, _00181_, _00179_);
  and _25522_ (_00183_, _00182_, _00178_);
  or _25523_ (_00184_, _00183_, _00120_);
  and _25524_ (_00185_, _00184_, _00171_);
  or _25525_ (_00186_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or _25526_ (_00187_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _00071_);
  and _25527_ (_00188_, _00187_, _00186_);
  or _25528_ (_00189_, _00188_, _00069_);
  or _25529_ (_00190_, _00075_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _25530_ (_00191_, _00190_, _00189_);
  or _25531_ (_00192_, _00191_, _00089_);
  nand _25532_ (_00193_, _00097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not _25533_ (_00194_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _25534_ (_00195_, _00101_, _00194_);
  and _25535_ (_00196_, _00195_, _00193_);
  nand _25536_ (_00197_, _00196_, _00192_);
  or _25537_ (_00198_, _00197_, _00007_);
  nand _25538_ (_00199_, _00198_, _00013_);
  nand _25539_ (_00200_, _00199_, _00185_);
  and _25540_ (_00201_, _00200_, _00164_);
  not _25541_ (_00202_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _25542_ (_00203_, _00039_, _00202_);
  nand _25543_ (_00204_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _25544_ (_00205_, _00204_, _00203_);
  nand _25545_ (_00206_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nand _25546_ (_00207_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _25547_ (_00208_, _00207_, _00206_);
  and _25548_ (_00209_, _00208_, _00205_);
  or _25549_ (_00210_, _00126_, _00078_);
  nand _25550_ (_00211_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nand _25551_ (_00212_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _25552_ (_00213_, _00212_, _00211_);
  and _25553_ (_00214_, _00213_, _00210_);
  and _25554_ (_00215_, _00214_, _00209_);
  not _25555_ (_00216_, _00215_);
  and _25556_ (_00217_, _00216_, _00201_);
  and _25557_ (_00218_, _00217_, _00151_);
  and _25558_ (_00219_, _00088_, _00201_);
  not _25559_ (_00220_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _25560_ (_00221_, _00039_, _00220_);
  and _25561_ (_00222_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _25562_ (_00223_, _00222_, _00221_);
  and _25563_ (_00224_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _25564_ (_00225_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _25565_ (_00226_, _00225_, _00224_);
  and _25566_ (_00227_, _00226_, _00223_);
  or _25567_ (_00228_, _00112_, _00078_);
  and _25568_ (_00229_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _25569_ (_00230_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _25570_ (_00231_, _00230_, _00229_);
  and _25571_ (_00232_, _00231_, _00228_);
  and _25572_ (_00233_, _00232_, _00227_);
  not _25573_ (_00234_, _00233_);
  and _25574_ (_00235_, _00234_, _00150_);
  nand _25575_ (_00236_, _00235_, _00219_);
  and _25576_ (_00237_, _00234_, _00201_);
  or _25577_ (_00238_, _00237_, _00151_);
  and _25578_ (_00239_, _00238_, _00236_);
  and _25579_ (_00240_, _00239_, _00218_);
  not _25580_ (_00241_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _25581_ (_00242_, _00039_, _00241_);
  and _25582_ (_00243_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _25583_ (_00244_, _00243_, _00242_);
  and _25584_ (_00245_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and _25585_ (_00246_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _25586_ (_00247_, _00246_, _00245_);
  and _25587_ (_00248_, _00247_, _00244_);
  or _25588_ (_00249_, _00078_, _00157_);
  and _25589_ (_00250_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _25590_ (_00251_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _25591_ (_00252_, _00251_, _00250_);
  and _25592_ (_00253_, _00252_, _00249_);
  and _25593_ (_00254_, _00253_, _00248_);
  or _25594_ (_00255_, _00254_, _00236_);
  not _25595_ (_00256_, _00254_);
  and _25596_ (_00257_, _00256_, _00201_);
  not _25597_ (_00258_, _00257_);
  nand _25598_ (_00259_, _00258_, _00236_);
  and _25599_ (_00260_, _00259_, _00255_);
  nand _25600_ (_00261_, _00260_, _00235_);
  or _25601_ (_00262_, _00257_, _00235_);
  and _25602_ (_00263_, _00262_, _00261_);
  nand _25603_ (_00264_, _00263_, _00240_);
  not _25604_ (_00265_, _00264_);
  not _25605_ (_00266_, _00255_);
  and _25606_ (_00267_, _00260_, _00235_);
  nand _25607_ (_00268_, _00149_, _00105_);
  or _25608_ (_00269_, _00254_, _00268_);
  nand _25609_ (_00270_, _00200_, _00164_);
  not _25610_ (_00271_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _25611_ (_00272_, _00039_, _00271_);
  and _25612_ (_00273_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _25613_ (_00274_, _00273_, _00272_);
  and _25614_ (_00275_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _25615_ (_00276_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _25616_ (_00277_, _00276_, _00275_);
  and _25617_ (_00278_, _00277_, _00274_);
  nor _25618_ (_00279_, _00095_, _00078_);
  and _25619_ (_00280_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _25620_ (_00281_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _25621_ (_00282_, _00281_, _00280_);
  not _25622_ (_00283_, _00282_);
  nor _25623_ (_00284_, _00283_, _00279_);
  and _25624_ (_00285_, _00284_, _00278_);
  or _25625_ (_00286_, _00285_, _00270_);
  or _25626_ (_00287_, _00286_, _00269_);
  nand _25627_ (_00288_, _00286_, _00269_);
  and _25628_ (_00289_, _00288_, _00287_);
  nand _25629_ (_00290_, _00289_, _00267_);
  or _25630_ (_00291_, _00289_, _00267_);
  and _25631_ (_00292_, _00291_, _00290_);
  nand _25632_ (_00293_, _00292_, _00266_);
  or _25633_ (_00294_, _00292_, _00266_);
  and _25634_ (_00295_, _00294_, _00293_);
  nand _25635_ (_00296_, _00295_, _00265_);
  or _25636_ (_00297_, _00295_, _00265_);
  nand _25637_ (_00298_, _00297_, _00296_);
  not _25638_ (_00299_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _25639_ (_00300_, _00039_, _00299_);
  nand _25640_ (_00301_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _25641_ (_00302_, _00301_, _00300_);
  nand _25642_ (_00303_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nand _25643_ (_00304_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _25644_ (_00305_, _00304_, _00303_);
  and _25645_ (_00306_, _00305_, _00302_);
  or _25646_ (_00307_, _00140_, _00078_);
  nand _25647_ (_00308_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand _25648_ (_00309_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _25649_ (_00310_, _00309_, _00308_);
  and _25650_ (_00311_, _00310_, _00307_);
  nand _25651_ (_00312_, _00311_, _00306_);
  and _25652_ (_00313_, _00312_, _00150_);
  nand _25653_ (_00314_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand _25654_ (_00315_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _25655_ (_00316_, _00315_, _00314_);
  not _25656_ (_00317_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _25657_ (_00318_, _00039_, _00317_);
  nand _25658_ (_00319_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _25659_ (_00320_, _00319_, _00318_);
  and _25660_ (_00321_, _00320_, _00316_);
  or _25661_ (_00322_, _00078_, _00177_);
  nand _25662_ (_00323_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand _25663_ (_00324_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _25664_ (_00325_, _00324_, _00323_);
  and _25665_ (_00326_, _00325_, _00322_);
  nand _25666_ (_00327_, _00326_, _00321_);
  and _25667_ (_00328_, _00327_, _00201_);
  and _25668_ (_00329_, _00328_, _00313_);
  not _25669_ (_00330_, _00329_);
  and _25670_ (_00331_, _00312_, _00201_);
  not _25671_ (_00332_, _00331_);
  and _25672_ (_00333_, _00327_, _00150_);
  and _25673_ (_00334_, _00333_, _00332_);
  nand _25674_ (_00335_, _00334_, _00217_);
  nand _25675_ (_00336_, _00335_, _00330_);
  not _25676_ (_00337_, _00218_);
  and _25677_ (_00338_, _00216_, _00150_);
  or _25678_ (_00339_, _00338_, _00219_);
  and _25679_ (_00340_, _00339_, _00337_);
  and _25680_ (_00341_, _00340_, _00336_);
  not _25681_ (_00342_, _00240_);
  or _25682_ (_00343_, _00239_, _00218_);
  and _25683_ (_00344_, _00343_, _00342_);
  and _25684_ (_00345_, _00344_, _00341_);
  or _25685_ (_00346_, _00263_, _00240_);
  and _25686_ (_00347_, _00346_, _00264_);
  nand _25687_ (_00348_, _00347_, _00345_);
  not _25688_ (_00349_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _25689_ (_00350_, _00039_, _00349_);
  and _25690_ (_00351_, _00045_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _25691_ (_00352_, _00351_, _00350_);
  and _25692_ (_00353_, _00053_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _25693_ (_00354_, _00059_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _25694_ (_00355_, _00354_, _00353_);
  and _25695_ (_00356_, _00355_, _00352_);
  nor _25696_ (_00357_, _00078_, _00191_);
  and _25697_ (_00358_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _25698_ (_00359_, _00081_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor _25699_ (_00360_, _00359_, _00358_);
  not _25700_ (_00361_, _00360_);
  nor _25701_ (_00362_, _00361_, _00357_);
  and _25702_ (_00363_, _00362_, _00356_);
  not _25703_ (_00364_, _00363_);
  and _25704_ (_00365_, _00364_, _00150_);
  and _25705_ (_00366_, _00365_, _00331_);
  or _25706_ (_00367_, _00328_, _00313_);
  and _25707_ (_00368_, _00367_, _00330_);
  and _25708_ (_00369_, _00368_, _00366_);
  or _25709_ (_00370_, _00334_, _00217_);
  and _25710_ (_00371_, _00370_, _00335_);
  nand _25711_ (_00372_, _00371_, _00369_);
  not _25712_ (_00373_, _00372_);
  nand _25713_ (_00374_, _00340_, _00336_);
  or _25714_ (_00375_, _00340_, _00336_);
  and _25715_ (_00376_, _00375_, _00374_);
  nand _25716_ (_00377_, _00376_, _00373_);
  nand _25717_ (_00378_, _00344_, _00341_);
  or _25718_ (_00379_, _00344_, _00341_);
  nand _25719_ (_00380_, _00379_, _00378_);
  or _25720_ (_00381_, _00380_, _00377_);
  or _25721_ (_00382_, _00347_, _00345_);
  nand _25722_ (_00383_, _00382_, _00348_);
  or _25723_ (_00384_, _00383_, _00381_);
  and _25724_ (_00385_, _00384_, _00348_);
  or _25725_ (_00386_, _00385_, _00298_);
  nand _25726_ (_00387_, _00386_, _00296_);
  not _25727_ (_00388_, _00285_);
  and _25728_ (_00389_, _00388_, _00150_);
  and _25729_ (_00390_, _00389_, _00258_);
  and _25730_ (_00391_, _00293_, _00290_);
  not _25731_ (_00392_, _00391_);
  nand _25732_ (_00393_, _00392_, _00390_);
  or _25733_ (_00394_, _00392_, _00390_);
  and _25734_ (_00395_, _00394_, _00393_);
  nand _25735_ (_00396_, _00395_, _00387_);
  and _25736_ (_00397_, _00393_, _00287_);
  nand _25737_ (_00398_, _00397_, _00396_);
  nand _25738_ (_00399_, _00398_, _00029_);
  or _25739_ (_00400_, _00398_, _00029_);
  nand _25740_ (_00401_, _00400_, _00399_);
  and _25741_ (_00402_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or _25742_ (_00403_, _00395_, _00387_);
  and _25743_ (_00404_, _00403_, _00396_);
  nand _25744_ (_00405_, _00404_, _00402_);
  or _25745_ (_00406_, _00405_, _00401_);
  nand _25746_ (_00407_, _00406_, _00399_);
  and _25747_ (_00408_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _25748_ (_00409_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _25749_ (_00410_, _00409_, _00408_);
  and _25750_ (_00411_, _00410_, _00407_);
  and _25751_ (_00412_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand _25752_ (_00413_, _00385_, _00298_);
  and _25753_ (_00414_, _00413_, _00386_);
  nand _25754_ (_00415_, _00414_, _00412_);
  or _25755_ (_00416_, _00414_, _00412_);
  nand _25756_ (_00417_, _00416_, _00415_);
  and _25757_ (_00418_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nand _25758_ (_00419_, _00383_, _00381_);
  and _25759_ (_00420_, _00419_, _00384_);
  nand _25760_ (_00421_, _00420_, _00418_);
  or _25761_ (_00422_, _00420_, _00418_);
  nand _25762_ (_00423_, _00422_, _00421_);
  and _25763_ (_00424_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nand _25764_ (_00425_, _00380_, _00377_);
  and _25765_ (_00426_, _00425_, _00381_);
  nand _25766_ (_00427_, _00426_, _00424_);
  or _25767_ (_00428_, _00426_, _00424_);
  nand _25768_ (_00429_, _00428_, _00427_);
  and _25769_ (_00430_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or _25770_ (_00431_, _00376_, _00373_);
  and _25771_ (_00432_, _00431_, _00377_);
  nand _25772_ (_00433_, _00432_, _00430_);
  and _25773_ (_00434_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or _25774_ (_00435_, _00371_, _00369_);
  and _25775_ (_00436_, _00435_, _00372_);
  nand _25776_ (_00437_, _00436_, _00434_);
  and _25777_ (_00438_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand _25778_ (_00439_, _00368_, _00366_);
  or _25779_ (_00440_, _00368_, _00366_);
  and _25780_ (_00441_, _00440_, _00439_);
  and _25781_ (_00442_, _00441_, _00438_);
  not _25782_ (_00443_, _00442_);
  or _25783_ (_00444_, _00436_, _00434_);
  nand _25784_ (_00445_, _00444_, _00437_);
  or _25785_ (_00446_, _00445_, _00443_);
  and _25786_ (_00447_, _00446_, _00437_);
  or _25787_ (_00448_, _00432_, _00430_);
  nand _25788_ (_00449_, _00448_, _00433_);
  or _25789_ (_00450_, _00449_, _00447_);
  and _25790_ (_00451_, _00450_, _00433_);
  or _25791_ (_00452_, _00451_, _00429_);
  and _25792_ (_00453_, _00452_, _00427_);
  or _25793_ (_00454_, _00453_, _00423_);
  and _25794_ (_00455_, _00454_, _00421_);
  or _25795_ (_00456_, _00455_, _00417_);
  and _25796_ (_00457_, _00456_, _00415_);
  and _25797_ (_00458_, _00400_, _00399_);
  or _25798_ (_00459_, _00404_, _00402_);
  and _25799_ (_00460_, _00459_, _00405_);
  and _25800_ (_00461_, _00460_, _00458_);
  nand _25801_ (_00462_, _00410_, _00461_);
  nor _25802_ (_00463_, _00462_, _00457_);
  or _25803_ (_00464_, _00463_, _00411_);
  and _25804_ (_00465_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _25805_ (_00466_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _25806_ (_00467_, _00466_, _00465_);
  and _25807_ (_00468_, _00467_, _00464_);
  nand _25808_ (_00469_, _00468_, _00027_);
  and _25809_ (_00470_, _00025_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _25810_ (_00471_, _00470_, _00469_);
  or _25811_ (_00472_, _00469_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _25812_ (_00473_, _00472_, _00471_);
  and _25813_ (_25273_, _00473_, _25365_);
  nor _25814_ (_00474_, _00006_, _00009_);
  and _25815_ (_00475_, _00006_, _00009_);
  or _25816_ (_00476_, _00475_, _00474_);
  and _25817_ (_02734_, _00476_, _25365_);
  and _25818_ (_00477_, _00364_, _00201_);
  and _25819_ (_02921_, _00477_, _25365_);
  nor _25820_ (_00478_, _00365_, _00331_);
  nor _25821_ (_00479_, _00478_, _00366_);
  and _25822_ (_03120_, _00479_, _25365_);
  nor _25823_ (_00480_, _00441_, _00438_);
  nor _25824_ (_00481_, _00480_, _00442_);
  and _25825_ (_03308_, _00481_, _25365_);
  and _25826_ (_00482_, _00445_, _00443_);
  not _25827_ (_00483_, _00482_);
  and _25828_ (_00484_, _00483_, _00446_);
  and _25829_ (_03499_, _00484_, _25365_);
  and _25830_ (_00485_, _00449_, _00447_);
  not _25831_ (_00486_, _00485_);
  and _25832_ (_00487_, _00486_, _00450_);
  and _25833_ (_03687_, _00487_, _25365_);
  and _25834_ (_00489_, _00451_, _00429_);
  not _25835_ (_00490_, _00489_);
  and _25836_ (_00492_, _00490_, _00452_);
  and _25837_ (_03875_, _00492_, _25365_);
  and _25838_ (_00494_, _00453_, _00423_);
  not _25839_ (_00495_, _00494_);
  and _25840_ (_00497_, _00495_, _00454_);
  and _25841_ (_04060_, _00497_, _25365_);
  and _25842_ (_00499_, _00455_, _00417_);
  not _25843_ (_00500_, _00499_);
  and _25844_ (_00502_, _00500_, _00456_);
  and _25845_ (_04243_, _00502_, _25365_);
  not _25846_ (_00504_, _00460_);
  or _25847_ (_00505_, _00504_, _00457_);
  not _25848_ (_00507_, _00505_);
  and _25849_ (_00508_, _00504_, _00457_);
  nor _25850_ (_00510_, _00508_, _00507_);
  and _25851_ (_04339_, _00510_, _25365_);
  and _25852_ (_00512_, _00505_, _00405_);
  or _25853_ (_00513_, _00512_, _00401_);
  and _25854_ (_00515_, _00512_, _00401_);
  not _25855_ (_00516_, _00515_);
  and _25856_ (_00518_, _00516_, _00513_);
  and _25857_ (_04433_, _00518_, _25365_);
  nand _25858_ (_00520_, _00513_, _00399_);
  nand _25859_ (_00521_, _00520_, _00408_);
  or _25860_ (_00523_, _00520_, _00408_);
  and _25861_ (_00524_, _00523_, _00521_);
  and _25862_ (_04522_, _00524_, _25365_);
  not _25863_ (_00526_, _00409_);
  and _25864_ (_00528_, _00526_, _00521_);
  nor _25865_ (_00529_, _00528_, _00464_);
  and _25866_ (_04613_, _00529_, _25365_);
  nand _25867_ (_00531_, _00465_, _00464_);
  or _25868_ (_00533_, _00465_, _00464_);
  and _25869_ (_00534_, _00533_, _00531_);
  and _25870_ (_04706_, _00534_, _25365_);
  not _25871_ (_00536_, _00466_);
  and _25872_ (_00537_, _00536_, _00531_);
  nor _25873_ (_00538_, _00537_, _00468_);
  and _25874_ (_04792_, _00538_, _25365_);
  or _25875_ (_00539_, _00468_, _00027_);
  and _25876_ (_00540_, _00539_, _00469_);
  and _25877_ (_04876_, _00540_, _25365_);
  and _25878_ (_00541_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _00000_);
  nor _25879_ (_00542_, _00541_, _00001_);
  not _25880_ (_00543_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _25881_ (_00544_, _00003_, _00543_);
  and _25882_ (_00545_, _00544_, _00542_);
  and _25883_ (_00546_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _25884_ (_00547_, _00546_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _25885_ (_00548_, _00546_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _25886_ (_00549_, _00548_, _00547_);
  and _25887_ (_00881_, _00549_, _25365_);
  and _25888_ (_00912_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _25365_);
  nor _25889_ (_00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _25890_ (_00551_, _00550_, _00285_);
  nor _25891_ (_00552_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor _25892_ (_00553_, _00552_, _00551_);
  not _25893_ (_00554_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _25894_ (_00555_, _00197_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _25895_ (_00556_, _00183_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _25896_ (_00557_, _00556_, _00555_);
  and _25897_ (_00558_, _00557_, _00554_);
  not _25898_ (_00559_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _25899_ (_00560_, _00170_, _00559_);
  and _25900_ (_00561_, _00163_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _25901_ (_00562_, _00561_, _00560_);
  nor _25902_ (_00563_, _00562_, _00554_);
  nor _25903_ (_00564_, _00563_, _00558_);
  not _25904_ (_00565_, _00564_);
  and _25905_ (_00566_, _00565_, _00553_);
  nor _25906_ (_00567_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and _25907_ (_00568_, _00550_, _00254_);
  nor _25908_ (_00569_, _00568_, _00567_);
  not _25909_ (_00570_, _00569_);
  and _25910_ (_00571_, _00145_, _00141_);
  or _25911_ (_00572_, _00571_, _00559_);
  and _25912_ (_00573_, _00572_, _00554_);
  and _25913_ (_00574_, _00132_, _00559_);
  and _25914_ (_00575_, _00118_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _25915_ (_00576_, _00575_, _00574_);
  nor _25916_ (_00577_, _00576_, _00554_);
  nor _25917_ (_00578_, _00577_, _00573_);
  nor _25918_ (_00579_, _00578_, _00570_);
  nor _25919_ (_00580_, _00565_, _00553_);
  nor _25920_ (_00581_, _00580_, _00566_);
  and _25921_ (_00582_, _00581_, _00579_);
  nor _25922_ (_00583_, _00582_, _00566_);
  and _25923_ (_00584_, _00578_, _00570_);
  nor _25924_ (_00585_, _00584_, _00579_);
  and _25925_ (_00586_, _00585_, _00581_);
  and _25926_ (_00587_, _00550_, _00233_);
  nor _25927_ (_00588_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor _25928_ (_00589_, _00588_, _00587_);
  not _25929_ (_00590_, _00589_);
  nand _25930_ (_00591_, _00197_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _25931_ (_00592_, _00591_, _00554_);
  and _25932_ (_00593_, _00183_, _00559_);
  and _25933_ (_00594_, _00170_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _25934_ (_00595_, _00594_, _00593_);
  nor _25935_ (_00596_, _00595_, _00554_);
  nor _25936_ (_00597_, _00596_, _00592_);
  nor _25937_ (_00598_, _00597_, _00590_);
  and _25938_ (_00599_, _00597_, _00590_);
  nor _25939_ (_00600_, _00599_, _00598_);
  or _25940_ (_00601_, _00146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _25941_ (_00602_, _00132_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _25942_ (_00603_, _00602_, _00601_);
  and _25943_ (_00604_, _00603_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _25944_ (_00605_, _00604_);
  nand _25945_ (_00606_, _00550_, _00087_);
  nor _25946_ (_00607_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _25947_ (_00608_, _00607_);
  and _25948_ (_00609_, _00608_, _00606_);
  nand _25949_ (_00610_, _00609_, _00605_);
  nor _25950_ (_00611_, _00557_, _00554_);
  not _25951_ (_00612_, _00611_);
  nor _25952_ (_00613_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _25953_ (_00614_, _00613_);
  nand _25954_ (_00615_, _00550_, _00215_);
  and _25955_ (_00616_, _00615_, _00614_);
  nand _25956_ (_00617_, _00616_, _00612_);
  or _25957_ (_00618_, _00616_, _00612_);
  nand _25958_ (_00619_, _00618_, _00617_);
  or _25959_ (_00620_, _00572_, _00554_);
  nor _25960_ (_00621_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _25961_ (_00622_, _00621_);
  not _25962_ (_00623_, _00550_);
  or _25963_ (_00624_, _00623_, _00327_);
  and _25964_ (_00625_, _00624_, _00622_);
  nand _25965_ (_00626_, _00625_, _00620_);
  nor _25966_ (_00627_, _00591_, _00554_);
  or _25967_ (_00628_, _00623_, _00312_);
  nor _25968_ (_00629_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _25969_ (_00630_, _00629_);
  nand _25970_ (_00631_, _00630_, _00628_);
  and _25971_ (_00632_, _00631_, _00627_);
  or _25972_ (_00633_, _00625_, _00620_);
  nand _25973_ (_00634_, _00633_, _00626_);
  or _25974_ (_00635_, _00634_, _00632_);
  and _25975_ (_00636_, _00635_, _00626_);
  or _25976_ (_00637_, _00636_, _00619_);
  and _25977_ (_00638_, _00637_, _00617_);
  or _25978_ (_00639_, _00609_, _00605_);
  nand _25979_ (_00640_, _00639_, _00610_);
  or _25980_ (_00641_, _00640_, _00638_);
  nand _25981_ (_00642_, _00641_, _00610_);
  and _25982_ (_00643_, _00642_, _00600_);
  or _25983_ (_00644_, _00643_, _00598_);
  nand _25984_ (_00645_, _00644_, _00586_);
  nand _25985_ (_00646_, _00645_, _00583_);
  nor _25986_ (_00647_, _00603_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _25987_ (_00648_, _00118_, _00559_);
  and _25988_ (_00649_, _00104_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _25989_ (_00650_, _00649_, _00648_);
  nor _25990_ (_00651_, _00650_, _00554_);
  nor _25991_ (_00652_, _00651_, _00647_);
  not _25992_ (_00653_, _00652_);
  and _25993_ (_00654_, _00104_, _00163_);
  nor _25994_ (_00655_, _00654_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _25995_ (_00656_, _00595_, _00562_);
  nor _25996_ (_00657_, _00650_, _00576_);
  and _25997_ (_00658_, _00657_, _00656_);
  nor _25998_ (_00659_, _00658_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _25999_ (_00660_, _00659_, _00655_);
  and _26000_ (_00661_, _00660_, _00653_);
  and _26001_ (_00662_, _00661_, _00646_);
  or _26002_ (_00663_, _00662_, _00553_);
  and _26003_ (_00664_, _00644_, _00585_);
  nor _26004_ (_00665_, _00664_, _00579_);
  or _26005_ (_00666_, _00665_, _00581_);
  nand _26006_ (_00667_, _00666_, _00662_);
  and _26007_ (_00668_, _00667_, _00663_);
  and _26008_ (_00669_, _00668_, _00653_);
  nor _26009_ (_00670_, _00668_, _00653_);
  nor _26010_ (_00671_, _00644_, _00585_);
  or _26011_ (_00672_, _00671_, _00664_);
  nand _26012_ (_00673_, _00672_, _00662_);
  or _26013_ (_00674_, _00662_, _00569_);
  and _26014_ (_00675_, _00674_, _00673_);
  nand _26015_ (_00676_, _00675_, _00565_);
  nor _26016_ (_00677_, _00676_, _00670_);
  nor _26017_ (_00678_, _00677_, _00669_);
  or _26018_ (_00679_, _00670_, _00669_);
  or _26019_ (_00680_, _00675_, _00565_);
  and _26020_ (_00681_, _00680_, _00676_);
  not _26021_ (_00682_, _00681_);
  or _26022_ (_00683_, _00682_, _00679_);
  not _26023_ (_00684_, _00578_);
  nand _26024_ (_00685_, _00661_, _00646_);
  nor _26025_ (_00686_, _00642_, _00600_);
  nor _26026_ (_00687_, _00686_, _00643_);
  or _26027_ (_00688_, _00687_, _00685_);
  or _26028_ (_00689_, _00662_, _00589_);
  and _26029_ (_00690_, _00689_, _00688_);
  and _26030_ (_00691_, _00690_, _00684_);
  not _26031_ (_00692_, _00597_);
  and _26032_ (_00693_, _00640_, _00638_);
  not _26033_ (_00694_, _00693_);
  and _26034_ (_00695_, _00694_, _00641_);
  or _26035_ (_00696_, _00695_, _00685_);
  or _26036_ (_00697_, _00662_, _00609_);
  and _26037_ (_00698_, _00697_, _00696_);
  and _26038_ (_00699_, _00698_, _00692_);
  not _26039_ (_00700_, _00699_);
  nor _26040_ (_00701_, _00690_, _00684_);
  or _26041_ (_00702_, _00701_, _00691_);
  nor _26042_ (_00703_, _00702_, _00700_);
  nor _26043_ (_00704_, _00703_, _00691_);
  or _26044_ (_00705_, _00704_, _00683_);
  and _26045_ (_00706_, _00705_, _00678_);
  and _26046_ (_00707_, _00636_, _00619_);
  not _26047_ (_00708_, _00707_);
  and _26048_ (_00709_, _00708_, _00637_);
  or _26049_ (_00710_, _00709_, _00685_);
  or _26050_ (_00711_, _00662_, _00616_);
  and _26051_ (_00712_, _00711_, _00710_);
  and _26052_ (_00713_, _00712_, _00605_);
  and _26053_ (_00714_, _00634_, _00632_);
  not _26054_ (_00715_, _00714_);
  and _26055_ (_00716_, _00715_, _00635_);
  or _26056_ (_00717_, _00716_, _00685_);
  or _26057_ (_00718_, _00662_, _00625_);
  and _26058_ (_00719_, _00718_, _00717_);
  nand _26059_ (_00720_, _00719_, _00612_);
  nand _26060_ (_00721_, _00711_, _00710_);
  and _26061_ (_00722_, _00721_, _00604_);
  or _26062_ (_00723_, _00713_, _00722_);
  nor _26063_ (_00724_, _00723_, _00720_);
  or _26064_ (_00725_, _00724_, _00713_);
  nor _26065_ (_00726_, _00662_, _00631_);
  not _26066_ (_00727_, _00627_);
  and _26067_ (_00728_, _00631_, _00727_);
  nor _26068_ (_00729_, _00631_, _00727_);
  nor _26069_ (_00730_, _00729_, _00728_);
  and _26070_ (_00731_, _00662_, _00730_);
  or _26071_ (_00732_, _00731_, _00726_);
  nand _26072_ (_00733_, _00732_, _00620_);
  or _26073_ (_00734_, _00732_, _00620_);
  nand _26074_ (_00735_, _00734_, _00733_);
  and _26075_ (_00736_, _00550_, _00363_);
  nor _26076_ (_00737_, _00550_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _26077_ (_00738_, _00737_, _00736_);
  nor _26078_ (_00739_, _00738_, _00727_);
  or _26079_ (_00740_, _00739_, _00735_);
  nand _26080_ (_00741_, _00740_, _00733_);
  or _26081_ (_00742_, _00719_, _00612_);
  and _26082_ (_00743_, _00742_, _00720_);
  nor _26083_ (_00744_, _00713_, _00722_);
  and _26084_ (_00745_, _00744_, _00743_);
  and _26085_ (_00746_, _00745_, _00741_);
  or _26086_ (_00747_, _00746_, _00725_);
  or _26087_ (_00748_, _00698_, _00692_);
  and _26088_ (_00749_, _00748_, _00700_);
  not _26089_ (_00750_, _00702_);
  nand _26090_ (_00751_, _00750_, _00749_);
  nor _26091_ (_00752_, _00751_, _00683_);
  nand _26092_ (_00753_, _00752_, _00747_);
  nand _26093_ (_00754_, _00753_, _00706_);
  and _26094_ (_00755_, _00754_, _00660_);
  or _26095_ (_00756_, _00755_, _00668_);
  nor _26096_ (_00757_, _00746_, _00725_);
  or _26097_ (_00758_, _00751_, _00757_);
  nand _26098_ (_00759_, _00758_, _00704_);
  nand _26099_ (_00760_, _00759_, _00681_);
  nand _26100_ (_00761_, _00760_, _00676_);
  nand _26101_ (_00762_, _00761_, _00679_);
  nand _26102_ (_00763_, _00762_, _00755_);
  and _26103_ (_00764_, _00763_, _00756_);
  and _26104_ (_00933_, _00764_, _25365_);
  and _26105_ (_02979_, _00755_, _25365_);
  and _26106_ (_02989_, _00662_, _25365_);
  and _26107_ (_03009_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _25365_);
  and _26108_ (_03028_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _25365_);
  and _26109_ (_03048_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _25365_);
  or _26110_ (_00765_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _26111_ (_00766_, _00546_, rst);
  and _26112_ (_03058_, _00766_, _00765_);
  nand _26113_ (_00767_, _00754_, _00660_);
  or _26114_ (_00768_, _00767_, _00727_);
  and _26115_ (_00769_, _00768_, _00738_);
  nor _26116_ (_00770_, _00768_, _00738_);
  or _26117_ (_00771_, _00770_, _00769_);
  and _26118_ (_03069_, _00771_, _25365_);
  and _26119_ (_00772_, _00739_, _00735_);
  not _26120_ (_00773_, _00772_);
  and _26121_ (_00774_, _00773_, _00740_);
  or _26122_ (_00775_, _00774_, _00767_);
  or _26123_ (_00776_, _00755_, _00732_);
  and _26124_ (_00777_, _00776_, _00775_);
  and _26125_ (_03079_, _00777_, _25365_);
  nand _26126_ (_00778_, _00743_, _00741_);
  or _26127_ (_00779_, _00743_, _00741_);
  nand _26128_ (_00780_, _00779_, _00778_);
  nand _26129_ (_00781_, _00780_, _00755_);
  or _26130_ (_00782_, _00755_, _00719_);
  and _26131_ (_00783_, _00782_, _00781_);
  and _26132_ (_03089_, _00783_, _25365_);
  and _26133_ (_00784_, _00778_, _00720_);
  or _26134_ (_00785_, _00784_, _00723_);
  nand _26135_ (_00786_, _00784_, _00723_);
  nand _26136_ (_00787_, _00786_, _00785_);
  nand _26137_ (_00788_, _00787_, _00755_);
  or _26138_ (_00789_, _00755_, _00712_);
  and _26139_ (_00790_, _00789_, _00788_);
  and _26140_ (_03100_, _00790_, _25365_);
  not _26141_ (_00791_, _00749_);
  or _26142_ (_00792_, _00791_, _00757_);
  or _26143_ (_00793_, _00749_, _00747_);
  nand _26144_ (_00794_, _00793_, _00792_);
  nand _26145_ (_00795_, _00794_, _00755_);
  or _26146_ (_00796_, _00755_, _00698_);
  and _26147_ (_00797_, _00796_, _00795_);
  and _26148_ (_03110_, _00797_, _25365_);
  and _26149_ (_00798_, _00792_, _00700_);
  nand _26150_ (_00799_, _00702_, _00798_);
  or _26151_ (_00800_, _00702_, _00798_);
  nand _26152_ (_00801_, _00800_, _00799_);
  nand _26153_ (_00802_, _00801_, _00755_);
  or _26154_ (_00803_, _00755_, _00690_);
  and _26155_ (_00804_, _00803_, _00802_);
  and _26156_ (_03121_, _00804_, _25365_);
  or _26157_ (_00805_, _00759_, _00681_);
  nand _26158_ (_00806_, _00805_, _00760_);
  nand _26159_ (_00807_, _00806_, _00755_);
  or _26160_ (_00808_, _00755_, _00675_);
  and _26161_ (_00809_, _00808_, _00807_);
  and _26162_ (_03131_, _00809_, _25365_);
  not _26163_ (_00810_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _26164_ (_00811_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _00000_);
  and _26165_ (_00812_, _00811_, _00810_);
  and _26166_ (_00813_, _00812_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _26167_ (_00814_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _26168_ (_00815_, _00814_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _26169_ (_00816_, _00814_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _26170_ (_00817_, _00816_, _00815_);
  and _26171_ (_00818_, _00817_, _00813_);
  nor _26172_ (_00819_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _26173_ (_00820_, _00819_, _00811_);
  and _26174_ (_00821_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _26175_ (_00822_, _00821_, _00818_);
  not _26176_ (_00823_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _26177_ (_00824_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _00000_);
  and _26178_ (_00825_, _00824_, _00823_);
  and _26179_ (_00826_, _00825_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _26180_ (_00827_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _26181_ (_00828_, _00825_, _00810_);
  and _26182_ (_00829_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  nor _26183_ (_00830_, _00819_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _26184_ (_00831_, _00830_, _00811_);
  and _26185_ (_00832_, _00831_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _26186_ (_00833_, _00832_, _00829_);
  nor _26187_ (_00834_, _00833_, _00827_);
  and _26188_ (_00835_, _00834_, _00822_);
  nor _26189_ (_00836_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _26190_ (_00837_, _00836_, _00814_);
  and _26191_ (_00838_, _00837_, _00813_);
  and _26192_ (_00839_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  nor _26193_ (_00840_, _00839_, _00838_);
  and _26194_ (_00841_, _00831_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  not _26195_ (_00842_, _00841_);
  and _26196_ (_00843_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _26197_ (_00844_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _26198_ (_00845_, _00844_, _00843_);
  and _26199_ (_00846_, _00845_, _00842_);
  and _26200_ (_00847_, _00846_, _00840_);
  and _26201_ (_00848_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and _26202_ (_00849_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _26203_ (_00850_, _00849_, _00848_);
  and _26204_ (_00851_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not _26205_ (_00852_, _00851_);
  not _26206_ (_00853_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _26207_ (_00854_, _00813_, _00853_);
  and _26208_ (_00855_, _00831_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _26209_ (_00856_, _00855_, _00854_);
  and _26210_ (_00857_, _00856_, _00852_);
  and _26211_ (_00858_, _00857_, _00850_);
  and _26212_ (_00859_, _00858_, _00847_);
  and _26213_ (_00860_, _00859_, _00835_);
  and _26214_ (_00861_, _00815_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _26215_ (_00862_, _00861_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _26216_ (_00863_, _00862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _26217_ (_00864_, _00863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _26218_ (_00865_, _00864_);
  not _26219_ (_00866_, _00813_);
  nor _26220_ (_00867_, _00863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _26221_ (_00868_, _00867_, _00866_);
  and _26222_ (_00869_, _00868_, _00865_);
  not _26223_ (_00870_, _00869_);
  and _26224_ (_00871_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _26225_ (_00872_, _00871_, _00811_);
  and _26226_ (_00873_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _26227_ (_00874_, _00873_, _00872_);
  and _26228_ (_00875_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _26229_ (_00876_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _26230_ (_00877_, _00876_, _00875_);
  and _26231_ (_00878_, _00877_, _00874_);
  and _26232_ (_00879_, _00878_, _00870_);
  nor _26233_ (_00880_, _00862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _26234_ (_00882_, _00880_);
  nor _26235_ (_00883_, _00863_, _00866_);
  and _26236_ (_00884_, _00883_, _00882_);
  not _26237_ (_00885_, _00884_);
  and _26238_ (_00886_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _26239_ (_00887_, _00886_, _00872_);
  and _26240_ (_00888_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _26241_ (_00889_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _26242_ (_00890_, _00889_, _00888_);
  and _26243_ (_00891_, _00890_, _00887_);
  and _26244_ (_00892_, _00891_, _00885_);
  nor _26245_ (_00893_, _00892_, _00879_);
  not _26246_ (_00894_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _26247_ (_00895_, _00864_, _00894_);
  and _26248_ (_00896_, _00864_, _00894_);
  nor _26249_ (_00897_, _00896_, _00895_);
  nor _26250_ (_00898_, _00897_, _00866_);
  not _26251_ (_00899_, _00898_);
  and _26252_ (_00900_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor _26253_ (_00901_, _00900_, _00872_);
  and _26254_ (_00902_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _26255_ (_00903_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor _26256_ (_00904_, _00903_, _00902_);
  and _26257_ (_00905_, _00904_, _00901_);
  and _26258_ (_00906_, _00905_, _00899_);
  not _26259_ (_00907_, _00906_);
  not _26260_ (_00908_, _00861_);
  nor _26261_ (_00909_, _00815_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _26262_ (_00910_, _00909_, _00866_);
  and _26263_ (_00911_, _00910_, _00908_);
  not _26264_ (_00913_, _00911_);
  and _26265_ (_00914_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and _26266_ (_00915_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _26267_ (_00916_, _00915_, _00914_);
  and _26268_ (_00917_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _26269_ (_00918_, _00831_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor _26270_ (_00919_, _00918_, _00917_);
  and _26271_ (_00920_, _00919_, _00916_);
  and _26272_ (_00921_, _00920_, _00913_);
  not _26273_ (_00922_, _00921_);
  and _26274_ (_00923_, _00820_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _26275_ (_00924_, _00923_, _00872_);
  and _26276_ (_00925_, _00826_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not _26277_ (_00926_, _00925_);
  and _26278_ (_00927_, _00926_, _00924_);
  nor _26279_ (_00928_, _00861_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _26280_ (_00929_, _00928_);
  nor _26281_ (_00930_, _00862_, _00866_);
  and _26282_ (_00931_, _00930_, _00929_);
  and _26283_ (_00932_, _00828_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and _26284_ (_00934_, _00831_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor _26285_ (_00935_, _00934_, _00932_);
  not _26286_ (_00936_, _00935_);
  nor _26287_ (_00937_, _00936_, _00931_);
  and _26288_ (_00938_, _00937_, _00927_);
  nor _26289_ (_00939_, _00938_, _00922_);
  and _26290_ (_00940_, _00939_, _00907_);
  and _26291_ (_00941_, _00940_, _00893_);
  nand _26292_ (_00942_, _00941_, _00860_);
  nand _26293_ (_00943_, _00764_, _00545_);
  nand _26294_ (_00944_, _00473_, _00006_);
  nor _26295_ (_00945_, _00233_, _00118_);
  and _26296_ (_00946_, _00233_, _00118_);
  nor _26297_ (_00947_, _00946_, _00945_);
  nor _26298_ (_00948_, _00087_, _00170_);
  and _26299_ (_00949_, _00087_, _00170_);
  nor _26300_ (_00950_, _00949_, _00948_);
  nor _26301_ (_00951_, _00215_, _00132_);
  and _26302_ (_00952_, _00215_, _00132_);
  nor _26303_ (_00953_, _00952_, _00951_);
  not _26304_ (_00954_, _00183_);
  and _26305_ (_00955_, _00327_, _00954_);
  nor _26306_ (_00956_, _00327_, _00954_);
  nor _26307_ (_00957_, _00956_, _00955_);
  not _26308_ (_00958_, _00957_);
  and _26309_ (_00959_, _00312_, _00146_);
  not _26310_ (_00960_, _00197_);
  nor _26311_ (_00961_, _00363_, _00960_);
  nor _26312_ (_00962_, _00312_, _00146_);
  nor _26313_ (_00963_, _00962_, _00959_);
  and _26314_ (_00964_, _00963_, _00961_);
  nor _26315_ (_00965_, _00964_, _00959_);
  nor _26316_ (_00966_, _00965_, _00958_);
  nor _26317_ (_00967_, _00966_, _00955_);
  nor _26318_ (_00968_, _00967_, _00953_);
  and _26319_ (_00969_, _00967_, _00953_);
  nor _26320_ (_00970_, _00969_, _00968_);
  nor _26321_ (_00971_, _00075_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not _26322_ (_00972_, _00971_);
  nor _26323_ (_00973_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _26324_ (_00974_, _00973_, _00073_);
  and _26325_ (_00975_, _00974_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not _26326_ (_00976_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _26327_ (_00977_, _00976_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _26328_ (_00978_, _00977_, _00154_);
  nor _26329_ (_00979_, _00976_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _26330_ (_00980_, _00979_, _00109_);
  and _26331_ (_00981_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _26332_ (_00982_, _00981_, _00092_);
  and _26333_ (_00983_, _00982_, _00980_);
  and _26334_ (_00984_, _00983_, _00978_);
  nand _26335_ (_00985_, _00984_, _00975_);
  not _26336_ (_00986_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _26337_ (_00987_, _00973_, _00188_);
  and _26338_ (_00988_, _00987_, _00986_);
  nand _26339_ (_00989_, _00981_, _00123_);
  nand _26340_ (_00990_, _00979_, _00137_);
  nand _26341_ (_00991_, _00977_, _00174_);
  and _26342_ (_00992_, _00991_, _00990_);
  and _26343_ (_00993_, _00992_, _00989_);
  nand _26344_ (_00994_, _00993_, _00988_);
  nand _26345_ (_00995_, _00994_, _00985_);
  nand _26346_ (_00996_, _00995_, _00075_);
  and _26347_ (_00997_, _00996_, _00972_);
  and _26348_ (_00998_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _26349_ (_00999_, _00998_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _26350_ (_01000_, _00999_);
  and _26351_ (_01001_, _01000_, _00997_);
  and _26352_ (_01002_, _01000_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _26353_ (_01003_, _01002_, _01001_);
  and _26354_ (_01004_, _00363_, _00960_);
  nor _26355_ (_01005_, _01004_, _00961_);
  not _26356_ (_01006_, _01005_);
  nor _26357_ (_01007_, _01006_, _01003_);
  and _26358_ (_01008_, _01007_, _00963_);
  and _26359_ (_01009_, _00965_, _00958_);
  nor _26360_ (_01010_, _01009_, _00966_);
  and _26361_ (_01011_, _01010_, _01008_);
  not _26362_ (_01012_, _01011_);
  nor _26363_ (_01013_, _01012_, _00970_);
  nor _26364_ (_01014_, _00967_, _00952_);
  or _26365_ (_01015_, _01014_, _00951_);
  or _26366_ (_01016_, _01015_, _01013_);
  and _26367_ (_01017_, _01016_, _00950_);
  and _26368_ (_01018_, _01017_, _00947_);
  nor _26369_ (_01019_, _00254_, _00163_);
  and _26370_ (_01020_, _00254_, _00163_);
  nor _26371_ (_01021_, _01020_, _01019_);
  not _26372_ (_01022_, _01021_);
  and _26373_ (_01023_, _00948_, _00947_);
  nor _26374_ (_01024_, _01023_, _00945_);
  nor _26375_ (_01025_, _01024_, _01022_);
  and _26376_ (_01026_, _01024_, _01022_);
  nor _26377_ (_01027_, _01026_, _01025_);
  and _26378_ (_01028_, _01027_, _01018_);
  nor _26379_ (_01029_, _01025_, _01019_);
  not _26380_ (_01030_, _01029_);
  nor _26381_ (_01031_, _01030_, _01028_);
  nor _26382_ (_01032_, _00285_, _00104_);
  and _26383_ (_01033_, _00285_, _00104_);
  nor _26384_ (_01034_, _01033_, _01032_);
  not _26385_ (_01035_, _01034_);
  and _26386_ (_01036_, _01035_, _01031_);
  nor _26387_ (_01037_, _01035_, _01031_);
  not _26388_ (_01038_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _26389_ (_01039_, _00541_, _01038_);
  and _26390_ (_01040_, _01039_, _00005_);
  not _26391_ (_01041_, _01040_);
  or _26392_ (_01042_, _01041_, _01037_);
  nor _26393_ (_01043_, _01042_, _01036_);
  not _26394_ (_01044_, _01043_);
  not _26395_ (_01045_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _26396_ (_01046_, _00001_, _01045_);
  and _26397_ (_01047_, _01046_, _00005_);
  not _26398_ (_01048_, _01047_);
  not _26399_ (_01049_, _00163_);
  nor _26400_ (_01050_, _00254_, _01049_);
  not _26401_ (_01051_, _00118_);
  nor _26402_ (_01052_, _00233_, _01051_);
  not _26403_ (_01053_, _00170_);
  and _26404_ (_01054_, _00087_, _01053_);
  nor _26405_ (_01055_, _01054_, _00947_);
  nor _26406_ (_01056_, _01055_, _01052_);
  nor _26407_ (_01057_, _01056_, _01021_);
  nor _26408_ (_01058_, _01057_, _01050_);
  and _26409_ (_01059_, _01056_, _01021_);
  nor _26410_ (_01060_, _01059_, _01057_);
  not _26411_ (_01061_, _01060_);
  and _26412_ (_01062_, _01054_, _00947_);
  nor _26413_ (_01063_, _01062_, _01055_);
  not _26414_ (_01064_, _01063_);
  not _26415_ (_01065_, _00950_);
  and _26416_ (_01066_, _00363_, _00197_);
  nor _26417_ (_01067_, _01066_, _00963_);
  and _26418_ (_01068_, _00312_, _00571_);
  nor _26419_ (_01069_, _01068_, _01067_);
  nor _26420_ (_01070_, _01069_, _00957_);
  and _26421_ (_01071_, _00327_, _00183_);
  nor _26422_ (_01072_, _01071_, _01070_);
  nor _26423_ (_01073_, _01072_, _00953_);
  and _26424_ (_01074_, _01072_, _00953_);
  nor _26425_ (_01075_, _01074_, _01073_);
  not _26426_ (_01076_, _01075_);
  and _26427_ (_01077_, _01069_, _00957_);
  nor _26428_ (_01078_, _01077_, _01070_);
  not _26429_ (_01079_, _01078_);
  and _26430_ (_01080_, _01066_, _00963_);
  nor _26431_ (_01081_, _01080_, _01067_);
  not _26432_ (_01082_, _01081_);
  nor _26433_ (_01083_, _01005_, _01003_);
  and _26434_ (_01084_, _01083_, _01082_);
  and _26435_ (_01085_, _01084_, _01079_);
  and _26436_ (_01086_, _01085_, _01076_);
  not _26437_ (_01087_, _00132_);
  or _26438_ (_01088_, _00215_, _01087_);
  and _26439_ (_01089_, _00215_, _01087_);
  or _26440_ (_01090_, _01072_, _01089_);
  and _26441_ (_01091_, _01090_, _01088_);
  or _26442_ (_01092_, _01091_, _01086_);
  and _26443_ (_01093_, _01092_, _01065_);
  and _26444_ (_01094_, _01093_, _01064_);
  and _26445_ (_01095_, _01094_, _01061_);
  nor _26446_ (_01096_, _01095_, _01058_);
  nor _26447_ (_01097_, _01096_, _01034_);
  and _26448_ (_01098_, _01096_, _01034_);
  nor _26449_ (_01099_, _01098_, _01097_);
  nor _26450_ (_01100_, _01099_, _01048_);
  and _26451_ (_01101_, _00004_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _26452_ (_01102_, _01101_, _01046_);
  not _26453_ (_01103_, _00312_);
  nor _26454_ (_01104_, _00363_, _01103_);
  and _26455_ (_01105_, _01104_, _00327_);
  and _26456_ (_01106_, _01105_, _00216_);
  and _26457_ (_01107_, _01106_, _00088_);
  and _26458_ (_01108_, _01107_, _00234_);
  and _26459_ (_01109_, _01108_, _00256_);
  and _26460_ (_01110_, _01109_, _01003_);
  not _26461_ (_01111_, _01003_);
  and _26462_ (_01112_, _00254_, _00233_);
  nor _26463_ (_01113_, _00327_, _00312_);
  and _26464_ (_01114_, _01113_, _00363_);
  and _26465_ (_01115_, _01114_, _00215_);
  and _26466_ (_01116_, _01115_, _00087_);
  and _26467_ (_01117_, _01116_, _01112_);
  and _26468_ (_01118_, _01117_, _01111_);
  nor _26469_ (_01119_, _01118_, _01110_);
  and _26470_ (_01120_, _01119_, _00285_);
  nor _26471_ (_01121_, _01119_, _00285_);
  nor _26472_ (_01122_, _01121_, _01120_);
  and _26473_ (_01123_, _01122_, _01102_);
  not _26474_ (_01124_, _00104_);
  nor _26475_ (_01125_, _01003_, _01124_);
  not _26476_ (_01126_, _01125_);
  and _26477_ (_01127_, _01003_, _00285_);
  and _26478_ (_01128_, _01101_, _00002_);
  not _26479_ (_01129_, _01128_);
  nor _26480_ (_01130_, _01129_, _01127_);
  and _26481_ (_01131_, _01130_, _01126_);
  nor _26482_ (_01132_, _01131_, _01123_);
  not _26483_ (_01133_, _01112_);
  and _26484_ (_01134_, _01039_, _00544_);
  nor _26485_ (_01135_, _01113_, _00215_);
  and _26486_ (_01136_, _01135_, _01134_);
  and _26487_ (_01137_, _01136_, _00088_);
  nor _26488_ (_01138_, _01137_, _01133_);
  nor _26489_ (_01139_, _01112_, _00285_);
  nor _26490_ (_01140_, _01139_, _01136_);
  and _26491_ (_01141_, _01140_, _01003_);
  nor _26492_ (_01142_, _01141_, _01138_);
  and _26493_ (_01143_, _01142_, _00388_);
  not _26494_ (_01144_, _01134_);
  nor _26495_ (_01145_, _01142_, _00388_);
  or _26496_ (_01146_, _01145_, _01144_);
  nor _26497_ (_01147_, _01146_, _01143_);
  not _26498_ (_01148_, _01147_);
  not _26499_ (_01149_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _26500_ (_01150_, _00004_, _01149_);
  and _26501_ (_01151_, _01150_, _01039_);
  not _26502_ (_01152_, _01151_);
  nor _26503_ (_01153_, _01152_, _01033_);
  and _26504_ (_01154_, _01150_, _00542_);
  and _26505_ (_01155_, _01154_, _01034_);
  nor _26506_ (_01156_, _01155_, _01153_);
  and _26507_ (_01157_, _01150_, _00001_);
  not _26508_ (_01158_, _01157_);
  nor _26509_ (_01159_, _01158_, _00254_);
  and _26510_ (_01160_, _01101_, _00542_);
  and _26511_ (_01161_, _01160_, _00364_);
  nor _26512_ (_01162_, _01161_, _01159_);
  and _26513_ (_01163_, _01101_, _01039_);
  and _26514_ (_01164_, _01163_, _01111_);
  and _26515_ (_01165_, _00544_, _00002_);
  and _26516_ (_01166_, _01165_, _01032_);
  and _26517_ (_01167_, _01046_, _00544_);
  and _26518_ (_01168_, _01167_, _00285_);
  nor _26519_ (_01169_, _01168_, _01166_);
  and _26520_ (_01170_, _00542_, _00005_);
  not _26521_ (_01171_, _01170_);
  nor _26522_ (_01172_, _01171_, _00285_);
  not _26523_ (_01173_, _01172_);
  nand _26524_ (_01174_, _01173_, _01169_);
  nor _26525_ (_01175_, _01174_, _01164_);
  and _26526_ (_01176_, _01175_, _01162_);
  and _26527_ (_01177_, _01176_, _01156_);
  and _26528_ (_01178_, _01177_, _01148_);
  and _26529_ (_01179_, _01178_, _01132_);
  not _26530_ (_01180_, _01179_);
  nor _26531_ (_01181_, _01180_, _01100_);
  and _26532_ (_01182_, _01181_, _01044_);
  and _26533_ (_01183_, _01182_, _00944_);
  nand _26534_ (_01184_, _01183_, _00943_);
  or _26535_ (_01185_, _01184_, _00942_);
  not _26536_ (_01186_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _26537_ (_01187_, \oc8051_top_1.oc8051_decoder1.wr , _00000_);
  not _26538_ (_01188_, _01187_);
  nor _26539_ (_01189_, _01188_, _00812_);
  and _26540_ (_01190_, _01189_, _01186_);
  not _26541_ (_01191_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _26542_ (_01192_, _00942_, _01191_);
  and _26543_ (_01193_, _01192_, _01190_);
  and _26544_ (_01194_, _01193_, _01185_);
  nor _26545_ (_01195_, _01189_, _01191_);
  nor _26546_ (_01197_, _01037_, _01032_);
  nor _26547_ (_01199_, _01197_, _01041_);
  not _26548_ (_01201_, _01199_);
  and _26549_ (_01203_, _00285_, _01124_);
  nor _26550_ (_01205_, _01203_, _01097_);
  nor _26551_ (_01207_, _01205_, _01048_);
  and _26552_ (_01209_, _01138_, _01003_);
  nor _26553_ (_01211_, _01209_, _01127_);
  not _26554_ (_01213_, _01138_);
  nor _26555_ (_01215_, _01003_, _00285_);
  and _26556_ (_01217_, _01215_, _01213_);
  nor _26557_ (_01219_, _01217_, _01144_);
  and _26558_ (_01221_, _01219_, _01211_);
  not _26559_ (_01223_, _01221_);
  nor _26560_ (_01225_, _01002_, _00997_);
  not _26561_ (_01227_, _01154_);
  nor _26562_ (_01229_, _01227_, _01001_);
  nor _26563_ (_01231_, _01229_, _01151_);
  nor _26564_ (_01233_, _01231_, _01225_);
  not _26565_ (_01235_, _01160_);
  nor _26566_ (_01237_, _01235_, _01001_);
  nor _26567_ (_01239_, _01237_, _01003_);
  nor _26568_ (_01241_, _01167_, _01111_);
  nor _26569_ (_01243_, _01241_, _01239_);
  nor _26570_ (_01245_, _01243_, _01233_);
  nor _26571_ (_01247_, _01171_, _01003_);
  not _26572_ (_01249_, _01247_);
  and _26573_ (_01251_, _00999_, _00997_);
  and _26574_ (_01253_, _01150_, _01046_);
  and _26575_ (_01255_, _01165_, _00997_);
  nor _26576_ (_01257_, _01255_, _01253_);
  nor _26577_ (_01259_, _01257_, _01251_);
  not _26578_ (_01261_, _01259_);
  and _26579_ (_01263_, _01150_, _00002_);
  not _26580_ (_01265_, _01263_);
  nor _26581_ (_01267_, _01265_, _00285_);
  not _26582_ (_01269_, _01267_);
  and _26583_ (_01271_, _01163_, _00364_);
  nor _26584_ (_01273_, _01271_, _01136_);
  and _26585_ (_01275_, _01273_, _01269_);
  and _26586_ (_01277_, _01275_, _01261_);
  and _26587_ (_01279_, _01277_, _01249_);
  and _26588_ (_01281_, _01279_, _01245_);
  and _26589_ (_01283_, _01281_, _01223_);
  not _26590_ (_01285_, _01283_);
  nor _26591_ (_01287_, _01285_, _01207_);
  and _26592_ (_01289_, _01287_, _01201_);
  not _26593_ (_01291_, _00835_);
  nor _26594_ (_01293_, _00858_, _00847_);
  and _26595_ (_01294_, _01293_, _01291_);
  and _26596_ (_01295_, _01294_, _00941_);
  nand _26597_ (_01296_, _01295_, _01289_);
  or _26598_ (_01297_, _01295_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _26599_ (_01298_, _01189_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _26600_ (_01299_, _01298_, _01297_);
  and _26601_ (_01300_, _01299_, _01296_);
  or _26602_ (_01301_, _01300_, _01195_);
  or _26603_ (_01302_, _01301_, _01194_);
  and _26604_ (_08893_, _01302_, _25365_);
  nand _26605_ (_01303_, _00771_, _00545_);
  and _26606_ (_01304_, _00510_, _00006_);
  and _26607_ (_01305_, _01006_, _01003_);
  nor _26608_ (_01306_, _01305_, _01007_);
  not _26609_ (_01307_, _01306_);
  nor _26610_ (_01308_, _01047_, _01040_);
  nor _26611_ (_01309_, _01308_, _01307_);
  nor _26612_ (_01310_, _01265_, _01003_);
  not _26613_ (_01311_, _01310_);
  nor _26614_ (_01312_, _01227_, _00961_);
  nor _26615_ (_01313_, _01312_, _01151_);
  or _26616_ (_01314_, _01313_, _01004_);
  and _26617_ (_01315_, _01101_, _01038_);
  and _26618_ (_01316_, _01315_, _00312_);
  and _26619_ (_01317_, _01253_, _00388_);
  nor _26620_ (_01318_, _01317_, _01316_);
  and _26621_ (_01319_, _01165_, _00961_);
  and _26622_ (_01320_, _01167_, _00363_);
  nor _26623_ (_01321_, _01320_, _01319_);
  and _26624_ (_01322_, _01128_, _00197_);
  and _26625_ (_01323_, _01102_, _00363_);
  nor _26626_ (_01324_, _01323_, _01322_);
  nor _26627_ (_01325_, _01170_, _01134_);
  nor _26628_ (_01326_, _01325_, _00363_);
  not _26629_ (_01327_, _01326_);
  and _26630_ (_01328_, _01327_, _01324_);
  and _26631_ (_01329_, _01328_, _01321_);
  and _26632_ (_01330_, _01329_, _01318_);
  and _26633_ (_01331_, _01330_, _01314_);
  and _26634_ (_01332_, _01331_, _01311_);
  not _26635_ (_01333_, _01332_);
  nor _26636_ (_01334_, _01333_, _01309_);
  not _26637_ (_01335_, _01334_);
  nor _26638_ (_01336_, _01335_, _01304_);
  nand _26639_ (_01337_, _01336_, _01303_);
  or _26640_ (_01338_, _01337_, _00942_);
  not _26641_ (_01339_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _26642_ (_01340_, _00942_, _01339_);
  and _26643_ (_01341_, _01340_, _01190_);
  and _26644_ (_01342_, _01341_, _01338_);
  nor _26645_ (_01343_, _01189_, _01339_);
  not _26646_ (_01344_, _01289_);
  or _26647_ (_01345_, _01344_, _00942_);
  and _26648_ (_01346_, _01340_, _01298_);
  and _26649_ (_01347_, _01346_, _01345_);
  or _26650_ (_01348_, _01347_, _01343_);
  or _26651_ (_01349_, _01348_, _01342_);
  and _26652_ (_10754_, _01349_, _25365_);
  nand _26653_ (_01350_, _00777_, _00545_);
  nand _26654_ (_01351_, _00518_, _00006_);
  nor _26655_ (_01352_, _00963_, _00961_);
  or _26656_ (_01353_, _01352_, _00964_);
  and _26657_ (_01354_, _01353_, _01007_);
  nor _26658_ (_01355_, _01353_, _01007_);
  or _26659_ (_01356_, _01355_, _01354_);
  and _26660_ (_01357_, _01356_, _01040_);
  nor _26661_ (_01358_, _01135_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _26662_ (_01359_, _01358_, _00312_);
  nor _26663_ (_01360_, _01358_, _00312_);
  nor _26664_ (_01361_, _01360_, _01359_);
  nor _26665_ (_01362_, _01361_, _01144_);
  nor _26666_ (_01363_, _01152_, _00962_);
  and _26667_ (_01364_, _01154_, _00963_);
  nor _26668_ (_01365_, _01364_, _01363_);
  and _26669_ (_01366_, _01165_, _00959_);
  and _26670_ (_01367_, _01167_, _01103_);
  nor _26671_ (_01368_, _01367_, _01366_);
  and _26672_ (_01369_, _01170_, _00312_);
  not _26673_ (_01370_, _01369_);
  and _26674_ (_01371_, _01315_, _00327_);
  nor _26675_ (_01372_, _01158_, _00363_);
  nor _26676_ (_01373_, _01372_, _01371_);
  and _26677_ (_01374_, _01373_, _01370_);
  and _26678_ (_01375_, _01374_, _01368_);
  and _26679_ (_01376_, _01375_, _01365_);
  not _26680_ (_01377_, _01376_);
  nor _26681_ (_01378_, _01377_, _01362_);
  not _26682_ (_01379_, _01378_);
  nor _26683_ (_01380_, _01379_, _01357_);
  and _26684_ (_01381_, _01128_, _00146_);
  not _26685_ (_01382_, _01381_);
  and _26686_ (_01383_, _00363_, _01103_);
  nor _26687_ (_01384_, _01383_, _01104_);
  and _26688_ (_01385_, _01384_, _01111_);
  or _26689_ (_01386_, _01384_, _01111_);
  nand _26690_ (_01387_, _01386_, _01102_);
  or _26691_ (_01388_, _01387_, _01385_);
  and _26692_ (_01389_, _01388_, _01382_);
  nor _26693_ (_01390_, _01083_, _01082_);
  nor _26694_ (_01391_, _01390_, _01084_);
  nor _26695_ (_01392_, _01391_, _01048_);
  not _26696_ (_01393_, _01392_);
  and _26697_ (_01394_, _01393_, _01389_);
  and _26698_ (_01395_, _01394_, _01380_);
  and _26699_ (_01396_, _01395_, _01351_);
  nand _26700_ (_01397_, _01396_, _01350_);
  or _26701_ (_01398_, _01397_, _00942_);
  not _26702_ (_01399_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _26703_ (_01400_, _00942_, _01399_);
  and _26704_ (_01401_, _01400_, _01190_);
  and _26705_ (_01402_, _01401_, _01398_);
  nor _26706_ (_01403_, _01189_, _01399_);
  nand _26707_ (_01404_, _00941_, _00835_);
  not _26708_ (_01405_, _00858_);
  and _26709_ (_01406_, _01405_, _00847_);
  not _26710_ (_01407_, _01406_);
  nor _26711_ (_01408_, _01407_, _01404_);
  nand _26712_ (_01409_, _01408_, _01289_);
  or _26713_ (_01410_, _01408_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _26714_ (_01411_, _01410_, _01298_);
  and _26715_ (_01412_, _01411_, _01409_);
  or _26716_ (_01413_, _01412_, _01403_);
  or _26717_ (_01414_, _01413_, _01402_);
  and _26718_ (_10762_, _01414_, _25365_);
  nand _26719_ (_01415_, _00524_, _00006_);
  nand _26720_ (_01416_, _00783_, _00545_);
  nor _26721_ (_01417_, _01129_, _00183_);
  or _26722_ (_01418_, _01383_, _01003_);
  or _26723_ (_01419_, _01104_, _01111_);
  and _26724_ (_01420_, _01419_, _01418_);
  or _26725_ (_01421_, _01420_, _00327_);
  nand _26726_ (_01422_, _01420_, _00327_);
  and _26727_ (_01423_, _01422_, _01421_);
  and _26728_ (_01424_, _01423_, _01102_);
  nor _26729_ (_01425_, _01424_, _01417_);
  nor _26730_ (_01426_, _01084_, _01079_);
  nor _26731_ (_01427_, _01426_, _01085_);
  nor _26732_ (_01428_, _01427_, _01048_);
  not _26733_ (_01429_, _01428_);
  not _26734_ (_01430_, _01315_);
  nor _26735_ (_01431_, _01430_, _00215_);
  and _26736_ (_01432_, _01165_, _00955_);
  not _26737_ (_01433_, _00327_);
  and _26738_ (_01434_, _01167_, _01433_);
  nor _26739_ (_01435_, _01434_, _01432_);
  nor _26740_ (_01436_, _01152_, _00956_);
  and _26741_ (_01437_, _01154_, _00957_);
  nor _26742_ (_01438_, _01437_, _01436_);
  and _26743_ (_01439_, _01170_, _00327_);
  and _26744_ (_01440_, _01157_, _00312_);
  nor _26745_ (_01441_, _01440_, _01439_);
  and _26746_ (_01442_, _01441_, _01438_);
  nand _26747_ (_01443_, _01442_, _01435_);
  nor _26748_ (_01444_, _01443_, _01431_);
  and _26749_ (_01445_, _01444_, _01429_);
  nor _26750_ (_01446_, _01010_, _01008_);
  nor _26751_ (_01447_, _01446_, _01041_);
  and _26752_ (_01448_, _01447_, _01012_);
  nor _26753_ (_01449_, _01360_, _01433_);
  and _26754_ (_01450_, _01113_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _26755_ (_01451_, _01450_, _01449_);
  nor _26756_ (_01452_, _01451_, _01144_);
  nor _26757_ (_01453_, _01452_, _01448_);
  and _26758_ (_01454_, _01453_, _01445_);
  and _26759_ (_01455_, _01454_, _01425_);
  and _26760_ (_01456_, _01455_, _01416_);
  nand _26761_ (_01457_, _01456_, _01415_);
  or _26762_ (_01458_, _01457_, _00942_);
  not _26763_ (_01459_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _26764_ (_01460_, _00942_, _01459_);
  and _26765_ (_01461_, _01460_, _01190_);
  and _26766_ (_01462_, _01461_, _01458_);
  nor _26767_ (_01463_, _01189_, _01459_);
  or _26768_ (_01464_, _01293_, _01404_);
  and _26769_ (_01465_, _01464_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _26770_ (_01466_, _00847_);
  and _26771_ (_01467_, _00835_, _00858_);
  and _26772_ (_01468_, _01467_, _01466_);
  not _26773_ (_01469_, _01468_);
  nor _26774_ (_01470_, _01469_, _01289_);
  and _26775_ (_01471_, _00835_, _00847_);
  and _26776_ (_01472_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _26777_ (_01473_, _01472_, _01470_);
  and _26778_ (_01474_, _01473_, _00941_);
  or _26779_ (_01475_, _01474_, _01465_);
  and _26780_ (_01476_, _01475_, _01298_);
  or _26781_ (_01477_, _01476_, _01463_);
  or _26782_ (_01478_, _01477_, _01462_);
  and _26783_ (_10770_, _01478_, _25365_);
  nand _26784_ (_01479_, _00529_, _00006_);
  nand _26785_ (_01480_, _00790_, _00545_);
  and _26786_ (_01481_, _01012_, _00970_);
  or _26787_ (_01482_, _01481_, _01041_);
  nor _26788_ (_01483_, _01482_, _01013_);
  not _26789_ (_01484_, _01483_);
  nor _26790_ (_01485_, _01085_, _01076_);
  nor _26791_ (_01486_, _01485_, _01086_);
  nor _26792_ (_01487_, _01486_, _01048_);
  not _26793_ (_01488_, _01487_);
  nor _26794_ (_01489_, _01129_, _00132_);
  or _26795_ (_01490_, _01114_, _01003_);
  or _26796_ (_01491_, _01105_, _01111_);
  nand _26797_ (_01492_, _01491_, _01490_);
  and _26798_ (_01493_, _01492_, _00215_);
  or _26799_ (_01494_, _01492_, _00215_);
  nand _26800_ (_01495_, _01494_, _01102_);
  nor _26801_ (_01496_, _01495_, _01493_);
  nor _26802_ (_01497_, _01496_, _01489_);
  not _26803_ (_01498_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _26804_ (_01499_, _01113_, _01498_);
  nor _26805_ (_01500_, _01499_, _00216_);
  or _26806_ (_01501_, _01500_, _01144_);
  nor _26807_ (_01502_, _01501_, _01135_);
  not _26808_ (_01503_, _01502_);
  nor _26809_ (_01504_, _01152_, _00952_);
  and _26810_ (_01505_, _01154_, _00953_);
  nor _26811_ (_01506_, _01505_, _01504_);
  and _26812_ (_01507_, _01165_, _00951_);
  and _26813_ (_01508_, _01167_, _00215_);
  nor _26814_ (_01509_, _01508_, _01507_);
  nor _26815_ (_01510_, _01171_, _00215_);
  and _26816_ (_01511_, _01157_, _00327_);
  nor _26817_ (_01512_, _01430_, _00087_);
  or _26818_ (_01513_, _01512_, _01511_);
  nor _26819_ (_01514_, _01513_, _01510_);
  and _26820_ (_01515_, _01514_, _01509_);
  and _26821_ (_01516_, _01515_, _01506_);
  and _26822_ (_01517_, _01516_, _01503_);
  and _26823_ (_01518_, _01517_, _01497_);
  and _26824_ (_01519_, _01518_, _01488_);
  and _26825_ (_01520_, _01519_, _01484_);
  and _26826_ (_01521_, _01520_, _01480_);
  nand _26827_ (_01522_, _01521_, _01479_);
  or _26828_ (_01523_, _01522_, _00942_);
  not _26829_ (_01524_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _26830_ (_01525_, _00942_, _01524_);
  and _26831_ (_01526_, _01525_, _01190_);
  and _26832_ (_01527_, _01526_, _01523_);
  nor _26833_ (_01528_, _01189_, _01524_);
  and _26834_ (_01529_, _01404_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _26835_ (_01530_, _01293_, _00835_);
  and _26836_ (_01531_, _01530_, _01344_);
  or _26837_ (_01532_, _01293_, _01291_);
  nor _26838_ (_01533_, _01532_, _01524_);
  or _26839_ (_01534_, _01533_, _01531_);
  and _26840_ (_01535_, _01534_, _00941_);
  or _26841_ (_01536_, _01535_, _01529_);
  and _26842_ (_01537_, _01536_, _01298_);
  or _26843_ (_01538_, _01537_, _01528_);
  or _26844_ (_01539_, _01538_, _01527_);
  and _26845_ (_10777_, _01539_, _25365_);
  nand _26846_ (_01540_, _00797_, _00545_);
  nand _26847_ (_01541_, _00534_, _00006_);
  nor _26848_ (_01542_, _01016_, _00950_);
  nor _26849_ (_01543_, _01542_, _01017_);
  and _26850_ (_01544_, _01543_, _01040_);
  not _26851_ (_01545_, _01544_);
  nor _26852_ (_01546_, _01092_, _00950_);
  and _26853_ (_01547_, _01092_, _00950_);
  nor _26854_ (_01548_, _01547_, _01546_);
  and _26855_ (_01549_, _01548_, _01047_);
  and _26856_ (_01550_, _01003_, _00088_);
  nor _26857_ (_01551_, _01003_, _00170_);
  or _26858_ (_01552_, _01551_, _01550_);
  and _26859_ (_01553_, _01552_, _01128_);
  and _26860_ (_01554_, _01106_, _01003_);
  and _26861_ (_01555_, _01115_, _01111_);
  nor _26862_ (_01556_, _01555_, _01554_);
  nor _26863_ (_01557_, _01556_, _00087_);
  not _26864_ (_01558_, _01557_);
  not _26865_ (_01559_, _01102_);
  and _26866_ (_01560_, _01556_, _00087_);
  nor _26867_ (_01561_, _01560_, _01559_);
  and _26868_ (_01562_, _01561_, _01558_);
  nor _26869_ (_01563_, _01562_, _01553_);
  nor _26870_ (_01564_, _01136_, _00088_);
  not _26871_ (_01565_, _01564_);
  nor _26872_ (_01566_, _01137_, _01144_);
  and _26873_ (_01567_, _01566_, _01565_);
  not _26874_ (_01568_, _01567_);
  and _26875_ (_01569_, _01154_, _00950_);
  and _26876_ (_01570_, _01165_, _00948_);
  nor _26877_ (_01571_, _01152_, _00949_);
  and _26878_ (_01572_, _01167_, _00087_);
  or _26879_ (_01573_, _01572_, _01571_);
  or _26880_ (_01574_, _01573_, _01570_);
  nor _26881_ (_01575_, _01574_, _01569_);
  nor _26882_ (_01576_, _01171_, _00087_);
  not _26883_ (_01577_, _01576_);
  nor _26884_ (_01578_, _01430_, _00233_);
  nor _26885_ (_01579_, _01158_, _00215_);
  nor _26886_ (_01580_, _01579_, _01578_);
  and _26887_ (_01581_, _01580_, _01577_);
  and _26888_ (_01582_, _01581_, _01575_);
  and _26889_ (_01583_, _01582_, _01568_);
  and _26890_ (_01584_, _01583_, _01563_);
  not _26891_ (_01585_, _01584_);
  nor _26892_ (_01586_, _01585_, _01549_);
  and _26893_ (_01587_, _01586_, _01545_);
  and _26894_ (_01588_, _01587_, _01541_);
  nand _26895_ (_01589_, _01588_, _01540_);
  or _26896_ (_01590_, _01589_, _00942_);
  not _26897_ (_01591_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _26898_ (_01592_, _00942_, _01591_);
  and _26899_ (_01593_, _01592_, _01190_);
  and _26900_ (_01594_, _01593_, _01590_);
  nor _26901_ (_01595_, _01189_, _01591_);
  not _26902_ (_01596_, _00941_);
  and _26903_ (_01597_, _00859_, _01291_);
  nor _26904_ (_01598_, _00859_, _01291_);
  nor _26905_ (_01599_, _01598_, _01597_);
  or _26906_ (_01600_, _01599_, _01596_);
  and _26907_ (_01601_, _01600_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _26908_ (_01602_, _01597_, _01344_);
  and _26909_ (_01603_, _01598_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _26910_ (_01604_, _01603_, _01602_);
  and _26911_ (_01605_, _01604_, _00941_);
  or _26912_ (_01606_, _01605_, _01601_);
  and _26913_ (_01607_, _01606_, _01298_);
  or _26914_ (_01608_, _01607_, _01595_);
  or _26915_ (_01609_, _01608_, _01594_);
  and _26916_ (_10786_, _01609_, _25365_);
  nand _26917_ (_01610_, _00804_, _00545_);
  nand _26918_ (_01611_, _00538_, _00006_);
  nor _26919_ (_01612_, _01093_, _01064_);
  nor _26920_ (_01613_, _01612_, _01094_);
  nor _26921_ (_01614_, _01613_, _01048_);
  not _26922_ (_01615_, _01614_);
  nor _26923_ (_01616_, _00948_, _00947_);
  or _26924_ (_01617_, _01616_, _01023_);
  and _26925_ (_01618_, _01617_, _01017_);
  nor _26926_ (_01619_, _01617_, _01017_);
  or _26927_ (_01620_, _01619_, _01618_);
  and _26928_ (_01621_, _01620_, _01040_);
  nor _26929_ (_01622_, _01003_, _00118_);
  and _26930_ (_01623_, _01003_, _00234_);
  nor _26931_ (_01624_, _01623_, _01622_);
  nor _26932_ (_01626_, _01624_, _01129_);
  nor _26933_ (_01627_, _01107_, _01111_);
  nor _26934_ (_01629_, _01116_, _01003_);
  nor _26935_ (_01630_, _01629_, _01627_);
  and _26936_ (_01632_, _01630_, _00234_);
  nor _26937_ (_01633_, _01630_, _00234_);
  or _26938_ (_01635_, _01633_, _01559_);
  nor _26939_ (_01636_, _01635_, _01632_);
  nor _26940_ (_01638_, _01636_, _01626_);
  nor _26941_ (_01639_, _01137_, _00234_);
  not _26942_ (_01641_, _01141_);
  and _26943_ (_01642_, _01641_, _01639_);
  nor _26944_ (_01644_, _01141_, _01137_);
  nor _26945_ (_01645_, _01644_, _00233_);
  nor _26946_ (_01647_, _01645_, _01642_);
  nor _26947_ (_01648_, _01647_, _01144_);
  nor _26948_ (_01650_, _01152_, _00946_);
  and _26949_ (_01651_, _01154_, _00947_);
  nor _26950_ (_01653_, _01651_, _01650_);
  and _26951_ (_01654_, _01165_, _00945_);
  and _26952_ (_01656_, _01167_, _00233_);
  nor _26953_ (_01657_, _01656_, _01654_);
  nor _26954_ (_01658_, _01430_, _00254_);
  not _26955_ (_01659_, _01658_);
  nor _26956_ (_01660_, _01171_, _00233_);
  nor _26957_ (_01661_, _01158_, _00087_);
  nor _26958_ (_01662_, _01661_, _01660_);
  and _26959_ (_01663_, _01662_, _01659_);
  and _26960_ (_01664_, _01663_, _01657_);
  and _26961_ (_01665_, _01664_, _01653_);
  not _26962_ (_01666_, _01665_);
  nor _26963_ (_01667_, _01666_, _01648_);
  and _26964_ (_01668_, _01667_, _01638_);
  not _26965_ (_01669_, _01668_);
  nor _26966_ (_01670_, _01669_, _01621_);
  and _26967_ (_01671_, _01670_, _01615_);
  and _26968_ (_01672_, _01671_, _01611_);
  nand _26969_ (_01673_, _01672_, _01610_);
  or _26970_ (_01674_, _01673_, _00942_);
  not _26971_ (_01675_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _26972_ (_01676_, _00942_, _01675_);
  and _26973_ (_01677_, _01676_, _01190_);
  and _26974_ (_01678_, _01677_, _01674_);
  nor _26975_ (_01679_, _01189_, _01675_);
  and _26976_ (_01680_, _01406_, _01291_);
  and _26977_ (_01681_, _01680_, _00941_);
  nand _26978_ (_01682_, _01681_, _01289_);
  or _26979_ (_01683_, _01681_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _26980_ (_01684_, _01683_, _01298_);
  and _26981_ (_01685_, _01684_, _01682_);
  or _26982_ (_01686_, _01685_, _01679_);
  or _26983_ (_01687_, _01686_, _01678_);
  and _26984_ (_10793_, _01687_, _25365_);
  nand _26985_ (_01688_, _00809_, _00545_);
  nand _26986_ (_01689_, _00540_, _00006_);
  nor _26987_ (_01690_, _01094_, _01061_);
  nor _26988_ (_01691_, _01690_, _01095_);
  nor _26989_ (_01692_, _01691_, _01048_);
  not _26990_ (_01693_, _01692_);
  nor _26991_ (_01694_, _01027_, _01018_);
  not _26992_ (_01695_, _01694_);
  nor _26993_ (_01696_, _01041_, _01028_);
  and _26994_ (_01697_, _01696_, _01695_);
  and _26995_ (_01698_, _01003_, _00256_);
  nor _26996_ (_01699_, _01003_, _00163_);
  or _26997_ (_01700_, _01699_, _01698_);
  and _26998_ (_01701_, _01700_, _01128_);
  nor _26999_ (_01702_, _01003_, _00234_);
  nand _27000_ (_01703_, _01702_, _01116_);
  nand _27001_ (_01704_, _01108_, _01003_);
  and _27002_ (_01705_, _01704_, _01703_);
  nor _27003_ (_01706_, _01705_, _00254_);
  and _27004_ (_01707_, _01705_, _00254_);
  or _27005_ (_01708_, _01707_, _01559_);
  nor _27006_ (_01709_, _01708_, _01706_);
  nor _27007_ (_01710_, _01709_, _01701_);
  nor _27008_ (_01711_, _01642_, _00254_);
  and _27009_ (_01712_, _01642_, _00254_);
  nor _27010_ (_01713_, _01712_, _01711_);
  nor _27011_ (_01714_, _01713_, _01144_);
  and _27012_ (_01715_, _01154_, _01021_);
  nor _27013_ (_01716_, _01152_, _01020_);
  not _27014_ (_01717_, _01716_);
  and _27015_ (_01718_, _01165_, _01019_);
  and _27016_ (_01719_, _01167_, _00254_);
  nor _27017_ (_01720_, _01719_, _01718_);
  nand _27018_ (_01721_, _01720_, _01717_);
  nor _27019_ (_01722_, _01721_, _01715_);
  nor _27020_ (_01723_, _01430_, _00285_);
  not _27021_ (_01724_, _01723_);
  nor _27022_ (_01725_, _01171_, _00254_);
  nor _27023_ (_01726_, _01158_, _00233_);
  nor _27024_ (_01727_, _01726_, _01725_);
  and _27025_ (_01728_, _01727_, _01724_);
  and _27026_ (_01729_, _01728_, _01722_);
  not _27027_ (_01730_, _01729_);
  nor _27028_ (_01731_, _01730_, _01714_);
  and _27029_ (_01732_, _01731_, _01710_);
  not _27030_ (_01733_, _01732_);
  nor _27031_ (_01734_, _01733_, _01697_);
  and _27032_ (_01735_, _01734_, _01693_);
  and _27033_ (_01736_, _01735_, _01689_);
  nand _27034_ (_01737_, _01736_, _01688_);
  or _27035_ (_01738_, _01737_, _00942_);
  not _27036_ (_01739_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _27037_ (_01740_, _00942_, _01739_);
  and _27038_ (_01741_, _01740_, _01190_);
  and _27039_ (_01742_, _01741_, _01738_);
  nor _27040_ (_01743_, _01189_, _01739_);
  nor _27041_ (_01744_, _00835_, _00847_);
  and _27042_ (_01745_, _01744_, _00858_);
  and _27043_ (_01746_, _01745_, _00941_);
  nand _27044_ (_01747_, _01746_, _01289_);
  or _27045_ (_01748_, _01746_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _27046_ (_01749_, _01748_, _01298_);
  and _27047_ (_01750_, _01749_, _01747_);
  or _27048_ (_01751_, _01750_, _01743_);
  or _27049_ (_01752_, _01751_, _01742_);
  and _27050_ (_10801_, _01752_, _25365_);
  and _27051_ (_01753_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _27052_ (_01754_, _01753_);
  nor _27053_ (_01755_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or _27054_ (_01756_, _01755_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _27055_ (_01757_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _27056_ (_01758_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _27057_ (_01759_, _01758_, _01757_);
  and _27058_ (_01760_, _01755_, _00000_);
  and _27059_ (_01761_, _01760_, _01759_);
  and _27060_ (_01762_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _27061_ (_01763_, _01762_);
  not _27062_ (_01764_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _27063_ (_01765_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _27064_ (_01766_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _27065_ (_01767_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _27066_ (_01768_, _01767_);
  not _27067_ (_01769_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _27068_ (_01770_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _27069_ (_01771_, _01770_, _01769_);
  nand _27070_ (_01772_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not _27071_ (_01773_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _27072_ (_01774_, _01773_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _27073_ (_01775_, _01774_, _01769_);
  nand _27074_ (_01776_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _27075_ (_01777_, _01776_, _01772_);
  nor _27076_ (_01778_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _27077_ (_01779_, _01778_, _01769_);
  nand _27078_ (_01780_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _27079_ (_01781_, _01778_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _27080_ (_01782_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _27081_ (_01783_, _01782_, _01780_);
  and _27082_ (_01784_, _01778_, _01769_);
  nand _27083_ (_01785_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not _27084_ (_01786_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  not _27085_ (_01787_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _27086_ (_01788_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _01787_);
  nand _27087_ (_01789_, _01788_, _01769_);
  or _27088_ (_01790_, _01789_, _01786_);
  and _27089_ (_01791_, _01790_, _01785_);
  and _27090_ (_01792_, _01791_, _01783_);
  nand _27091_ (_01793_, _01792_, _01777_);
  and _27092_ (_01794_, _01793_, _01768_);
  and _27093_ (_01795_, _01794_, _01766_);
  or _27094_ (_01796_, _01795_, _01765_);
  nand _27095_ (_01797_, _01796_, _01764_);
  and _27096_ (_01798_, _01797_, _01763_);
  nand _27097_ (_01799_, _01798_, _01761_);
  not _27098_ (_01800_, _01759_);
  nor _27099_ (_01801_, _01760_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _27100_ (_01802_, _01801_, _01800_);
  and _27101_ (_01803_, _01802_, _01799_);
  and _27102_ (_01804_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not _27103_ (_01805_, _01804_);
  and _27104_ (_01806_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nand _27105_ (_01807_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _27106_ (_01808_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _27107_ (_01809_, _01808_, _01807_);
  nand _27108_ (_01810_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not _27109_ (_01811_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _27110_ (_01812_, _01789_, _01811_);
  and _27111_ (_01813_, _01812_, _01810_);
  nand _27112_ (_01814_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _27113_ (_01815_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _27114_ (_01816_, _01815_, _01814_);
  and _27115_ (_01817_, _01816_, _01813_);
  and _27116_ (_01818_, _01817_, _01809_);
  or _27117_ (_01819_, _01767_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _27118_ (_01820_, _01819_, _01818_);
  or _27119_ (_01821_, _01820_, _01806_);
  nand _27120_ (_01822_, _01821_, _01764_);
  and _27121_ (_01823_, _01822_, _01805_);
  nand _27122_ (_01824_, _01823_, _01761_);
  nor _27123_ (_01825_, _01760_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _27124_ (_01826_, _01825_, _01800_);
  and _27125_ (_01827_, _01826_, _01824_);
  and _27126_ (_01828_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _27127_ (_01829_, _01828_);
  and _27128_ (_01830_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand _27129_ (_01831_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _27130_ (_01832_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _27131_ (_01833_, _01832_, _01831_);
  nand _27132_ (_01834_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not _27133_ (_01835_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _27134_ (_01836_, _01789_, _01835_);
  and _27135_ (_01837_, _01836_, _01834_);
  nand _27136_ (_01838_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _27137_ (_01839_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _27138_ (_01840_, _01839_, _01838_);
  and _27139_ (_01841_, _01840_, _01837_);
  and _27140_ (_01842_, _01841_, _01833_);
  nor _27141_ (_01843_, _01842_, _01819_);
  or _27142_ (_01844_, _01843_, _01830_);
  nand _27143_ (_01845_, _01844_, _01764_);
  and _27144_ (_01846_, _01845_, _01829_);
  nand _27145_ (_01847_, _01846_, _01761_);
  nor _27146_ (_01848_, _01760_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _27147_ (_01849_, _01848_, _01800_);
  and _27148_ (_01850_, _01849_, _01847_);
  nor _27149_ (_01851_, _01850_, _01827_);
  and _27150_ (_01852_, _01851_, _01803_);
  and _27151_ (_01853_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _27152_ (_01854_, _01853_);
  and _27153_ (_01855_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand _27154_ (_01856_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand _27155_ (_01857_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _27156_ (_01858_, _01857_, _01856_);
  nand _27157_ (_01859_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _27158_ (_01860_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _27159_ (_01861_, _01860_, _01859_);
  nand _27160_ (_01862_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _27161_ (_01863_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _27162_ (_01864_, _01789_, _01863_);
  and _27163_ (_01865_, _01864_, _01862_);
  and _27164_ (_01866_, _01865_, _01861_);
  nand _27165_ (_01867_, _01866_, _01858_);
  nand _27166_ (_01868_, _01867_, _01768_);
  nor _27167_ (_01869_, _01868_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _27168_ (_01870_, _01869_, _01855_);
  nand _27169_ (_01871_, _01870_, _01764_);
  and _27170_ (_01872_, _01871_, _01854_);
  nand _27171_ (_01873_, _01872_, _01761_);
  nor _27172_ (_01874_, _01760_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _27173_ (_01875_, _01874_, _01800_);
  and _27174_ (_01876_, _01875_, _01873_);
  not _27175_ (_01877_, _01876_);
  not _27176_ (_01878_, _01761_);
  nand _27177_ (_01879_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _27178_ (_01880_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand _27179_ (_01881_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _27180_ (_01882_, _01881_, _01880_);
  and _27181_ (_01883_, _01882_, _01879_);
  nand _27182_ (_01884_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nand _27183_ (_01885_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _27184_ (_01886_, _01885_, _01884_);
  not _27185_ (_01887_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _27186_ (_01888_, _01789_, _01887_);
  and _27187_ (_01889_, _01888_, _01768_);
  and _27188_ (_01890_, _01889_, _01886_);
  nand _27189_ (_01891_, _01890_, _01883_);
  nor _27190_ (_01892_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _27191_ (_01893_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _01766_);
  or _27192_ (_01894_, _01893_, _01892_);
  nand _27193_ (_01895_, _01894_, _01764_);
  nor _27194_ (_01896_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _01764_);
  not _27195_ (_01897_, _01896_);
  and _27196_ (_01898_, _01897_, _01895_);
  or _27197_ (_01899_, _01898_, _01878_);
  nor _27198_ (_01900_, _01760_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _27199_ (_01901_, _01900_, _01800_);
  and _27200_ (_01902_, _01901_, _01899_);
  and _27201_ (_01903_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _27202_ (_01904_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _27203_ (_01905_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _27204_ (_01906_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _27205_ (_01907_, _01906_, _01905_);
  not _27206_ (_01908_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _27207_ (_01909_, _01789_, _01908_);
  nand _27208_ (_01910_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _27209_ (_01911_, _01910_, _01909_);
  nand _27210_ (_01912_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand _27211_ (_01913_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _27212_ (_01914_, _01913_, _01912_);
  nand _27213_ (_01915_, _01914_, _01911_);
  nor _27214_ (_01916_, _01915_, _01907_);
  or _27215_ (_01917_, _01916_, _01819_);
  and _27216_ (_01918_, _01917_, _01904_);
  nor _27217_ (_01919_, _01918_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _27218_ (_01920_, _01919_, _01903_);
  or _27219_ (_01921_, _01920_, _01878_);
  nor _27220_ (_01922_, _01760_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _27221_ (_01923_, _01922_, _01800_);
  and _27222_ (_01924_, _01923_, _01921_);
  and _27223_ (_01925_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _27224_ (_01926_, _01925_);
  nand _27225_ (_01927_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand _27226_ (_01928_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _27227_ (_01929_, _01928_, _01927_);
  nand _27228_ (_01930_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _27229_ (_01931_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _27230_ (_01932_, _01931_, _01930_);
  nand _27231_ (_01933_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  not _27232_ (_01934_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _27233_ (_01935_, _01789_, _01934_);
  and _27234_ (_01936_, _01935_, _01933_);
  and _27235_ (_01937_, _01936_, _01932_);
  nand _27236_ (_01938_, _01937_, _01929_);
  nand _27237_ (_01939_, _01938_, _01768_);
  nand _27238_ (_01940_, _01939_, _01766_);
  nor _27239_ (_01941_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _01766_);
  nor _27240_ (_01942_, _01941_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _27241_ (_01943_, _01942_, _01940_);
  and _27242_ (_01944_, _01943_, _01926_);
  nand _27243_ (_01945_, _01944_, _01761_);
  nor _27244_ (_01946_, _01760_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _27245_ (_01947_, _01946_, _01800_);
  and _27246_ (_01948_, _01947_, _01945_);
  nor _27247_ (_01949_, _01948_, _01924_);
  and _27248_ (_01950_, _01949_, _01902_);
  and _27249_ (_01951_, _01950_, _01877_);
  and _27250_ (_01952_, _01951_, _01852_);
  not _27251_ (_01953_, _01948_);
  and _27252_ (_01954_, _01953_, _01924_);
  not _27253_ (_01955_, _01902_);
  and _27254_ (_01956_, _01955_, _01876_);
  and _27255_ (_01957_, _01956_, _01954_);
  nand _27256_ (_01958_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nand _27257_ (_01959_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _27258_ (_01960_, _01959_, _01958_);
  not _27259_ (_01961_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _27260_ (_01962_, _01789_, _01961_);
  and _27261_ (_01963_, _01962_, _01768_);
  and _27262_ (_01964_, _01963_, _01960_);
  nand _27263_ (_01965_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nand _27264_ (_01966_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand _27265_ (_01967_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _27266_ (_01968_, _01967_, _01966_);
  and _27267_ (_01969_, _01968_, _01965_);
  nand _27268_ (_01970_, _01969_, _01964_);
  nor _27269_ (_01971_, _01970_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _27270_ (_01972_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _01766_);
  or _27271_ (_01973_, _01972_, _01971_);
  nand _27272_ (_01974_, _01973_, _01764_);
  nor _27273_ (_01975_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _01764_);
  not _27274_ (_01976_, _01975_);
  and _27275_ (_01977_, _01976_, _01974_);
  or _27276_ (_01978_, _01977_, _01878_);
  nor _27277_ (_01979_, _01760_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _27278_ (_01980_, _01979_, _01800_);
  and _27279_ (_01981_, _01980_, _01978_);
  not _27280_ (_01982_, _01850_);
  and _27281_ (_01983_, _01982_, _01827_);
  and _27282_ (_01984_, _01983_, _01981_);
  and _27283_ (_01985_, _01984_, _01957_);
  nor _27284_ (_01986_, _01985_, _01952_);
  not _27285_ (_01987_, _01981_);
  and _27286_ (_01988_, _01850_, _01827_);
  and _27287_ (_01989_, _01988_, _01803_);
  and _27288_ (_01990_, _01989_, _01987_);
  and _27289_ (_01991_, _01990_, _01957_);
  not _27290_ (_01992_, _01827_);
  and _27291_ (_01993_, _01850_, _01992_);
  and _27292_ (_01994_, _01993_, _01803_);
  and _27293_ (_01995_, _01994_, _01987_);
  and _27294_ (_01996_, _01995_, _01950_);
  nor _27295_ (_01997_, _01902_, _01876_);
  and _27296_ (_01998_, _01997_, _01949_);
  not _27297_ (_01999_, _01803_);
  and _27298_ (_02000_, _01988_, _01999_);
  and _27299_ (_02001_, _02000_, _01998_);
  or _27300_ (_02002_, _02001_, _01996_);
  nor _27301_ (_02003_, _02002_, _01991_);
  and _27302_ (_02004_, _02003_, _01986_);
  and _27303_ (_02005_, _01983_, _01999_);
  and _27304_ (_02006_, _02005_, _01987_);
  and _27305_ (_02007_, _02006_, _01957_);
  and _27306_ (_02008_, _02005_, _01981_);
  and _27307_ (_02009_, _02008_, _01951_);
  nor _27308_ (_02010_, _02009_, _02007_);
  and _27309_ (_02011_, _01983_, _01803_);
  and _27310_ (_02012_, _02011_, _01987_);
  and _27311_ (_02013_, _02012_, _01948_);
  nand _27312_ (_02014_, _01851_, _01999_);
  nor _27313_ (_02015_, _02014_, _01981_);
  and _27314_ (_02016_, _02015_, _01957_);
  not _27315_ (_02017_, _02016_);
  and _27316_ (_02018_, _01954_, _01902_);
  nand _27317_ (_02019_, _02018_, _02012_);
  nand _27318_ (_02020_, _02019_, _02017_);
  nor _27319_ (_02021_, _02020_, _02013_);
  and _27320_ (_02022_, _02021_, _02010_);
  and _27321_ (_02023_, _01995_, _01957_);
  and _27322_ (_02024_, _02000_, _01987_);
  and _27323_ (_02025_, _02024_, _01957_);
  or _27324_ (_02026_, _02025_, _02023_);
  and _27325_ (_02027_, _01981_, _01852_);
  nand _27326_ (_02028_, _02027_, _01998_);
  not _27327_ (_02029_, _01998_);
  or _27328_ (_02030_, _02014_, _01987_);
  or _27329_ (_02031_, _02030_, _02029_);
  and _27330_ (_02032_, _02031_, _02028_);
  and _27331_ (_02033_, _01987_, _01852_);
  and _27332_ (_02034_, _02033_, _01998_);
  not _27333_ (_02035_, _02034_);
  and _27334_ (_02036_, _02035_, _02032_);
  not _27335_ (_02037_, _02036_);
  nor _27336_ (_02038_, _02037_, _02026_);
  and _27337_ (_02039_, _02038_, _02022_);
  and _27338_ (_02040_, _02039_, _02004_);
  and _27339_ (_02041_, _02000_, _01981_);
  and _27340_ (_02042_, _02041_, _01957_);
  not _27341_ (_02043_, _01957_);
  nor _27342_ (_02044_, _02030_, _02043_);
  nor _27343_ (_02045_, _02044_, _02042_);
  and _27344_ (_02046_, _01993_, _01999_);
  and _27345_ (_02047_, _02046_, _01987_);
  and _27346_ (_02048_, _02047_, _01957_);
  and _27347_ (_02049_, _01998_, _02011_);
  nor _27348_ (_02050_, _02049_, _02048_);
  and _27349_ (_02051_, _02050_, _02045_);
  and _27350_ (_02052_, _02011_, _01981_);
  nand _27351_ (_02053_, _02052_, _01951_);
  nand _27352_ (_02054_, _02024_, _01951_);
  and _27353_ (_02055_, _02054_, _02053_);
  and _27354_ (_02056_, _02047_, _01950_);
  not _27355_ (_02057_, _02056_);
  and _27356_ (_02058_, _01994_, _01981_);
  nand _27357_ (_02059_, _02058_, _01951_);
  and _27358_ (_02060_, _02059_, _02057_);
  and _27359_ (_02061_, _02060_, _02055_);
  and _27360_ (_02062_, _02061_, _02051_);
  and _27361_ (_02063_, _02041_, _01951_);
  and _27362_ (_02064_, _02012_, _01951_);
  nor _27363_ (_02065_, _02064_, _02063_);
  and _27364_ (_02066_, _02046_, _01981_);
  or _27365_ (_02067_, _02066_, _01852_);
  and _27366_ (_02068_, _02067_, _01957_);
  and _27367_ (_02069_, _02066_, _01950_);
  and _27368_ (_02070_, _02006_, _01951_);
  or _27369_ (_02071_, _02070_, _02069_);
  nor _27370_ (_02072_, _02071_, _02068_);
  and _27371_ (_02073_, _02072_, _02065_);
  and _27372_ (_02074_, _02073_, _02062_);
  nand _27373_ (_02075_, _02074_, _02040_);
  nand _27374_ (_02076_, _02075_, _01756_);
  not _27375_ (_02077_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _27376_ (_02078_, _00000_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _27377_ (_02079_, _02078_, _02077_);
  and _27378_ (_02080_, _01998_, _01993_);
  and _27379_ (_02081_, _02080_, _02079_);
  and _27380_ (_02082_, \oc8051_top_1.oc8051_decoder1.state [0], _00000_);
  and _27381_ (_02083_, _02082_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _27382_ (_02084_, _02083_, _01952_);
  nor _27383_ (_02085_, _02084_, _02081_);
  nand _27384_ (_02086_, _02085_, _02076_);
  nand _27385_ (_02087_, _02086_, _00000_);
  and _27386_ (_02088_, _02087_, _01754_);
  not _27387_ (_02089_, _02088_);
  and _27388_ (_02090_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _27389_ (_02091_, _02090_);
  and _27390_ (_02092_, _02079_, _01998_);
  and _27391_ (_02093_, _02092_, _01994_);
  and _27392_ (_02094_, _02018_, _02000_);
  and _27393_ (_02095_, _01924_, _01902_);
  and _27394_ (_02096_, _01981_, _01953_);
  and _27395_ (_02097_, _02096_, _02095_);
  and _27396_ (_02098_, _02097_, _02005_);
  or _27397_ (_02099_, _02098_, _02094_);
  and _27398_ (_02100_, _02097_, _02011_);
  not _27399_ (_02101_, _02014_);
  and _27400_ (_02102_, _02018_, _02101_);
  nor _27401_ (_02103_, _02102_, _02100_);
  and _27402_ (_02104_, _02046_, _02097_);
  and _27403_ (_02105_, _02018_, _01852_);
  or _27404_ (_02106_, _02105_, _02104_);
  not _27405_ (_02107_, _02106_);
  nand _27406_ (_02108_, _02107_, _02103_);
  and _27407_ (_02109_, _01950_, _01876_);
  and _27408_ (_02110_, _02012_, _02109_);
  and _27409_ (_02111_, _02058_, _02109_);
  and _27410_ (_02112_, _02109_, _02005_);
  and _27411_ (_02113_, _02112_, _01981_);
  or _27412_ (_02114_, _02113_, _02111_);
  or _27413_ (_02115_, _02114_, _02110_);
  and _27414_ (_02116_, _02041_, _01998_);
  nor _27415_ (_02117_, _01981_, _01948_);
  and _27416_ (_02118_, _02117_, _02095_);
  and _27417_ (_02119_, _02118_, _02005_);
  or _27418_ (_02120_, _02119_, _02116_);
  and _27419_ (_02121_, _02046_, _02118_);
  and _27420_ (_02122_, _02118_, _01989_);
  or _27421_ (_02123_, _02122_, _02121_);
  and _27422_ (_02124_, _01949_, _01877_);
  and _27423_ (_02125_, _02124_, _01902_);
  and _27424_ (_02126_, _02125_, _01852_);
  and _27425_ (_02127_, _02118_, _01994_);
  or _27426_ (_02128_, _02127_, _02126_);
  or _27427_ (_02129_, _02128_, _02123_);
  or _27428_ (_02130_, _02129_, _02120_);
  or _27429_ (_02131_, _02130_, _02115_);
  or _27430_ (_02132_, _02131_, _02108_);
  or _27431_ (_02133_, _02132_, _02099_);
  or _27432_ (_02134_, _02084_, _01756_);
  and _27433_ (_02135_, _02134_, _02133_);
  or _27434_ (_02136_, _02135_, _02093_);
  nand _27435_ (_02137_, _02136_, _00000_);
  and _27436_ (_02138_, _02137_, _02091_);
  and _27437_ (_02139_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _27438_ (_02140_, _01756_);
  not _27439_ (_02141_, _02109_);
  nor _27440_ (_02142_, _02058_, _02008_);
  nor _27441_ (_02143_, _02142_, _02141_);
  nor _27442_ (_02144_, _02143_, _02110_);
  nor _27443_ (_02145_, _02144_, _02140_);
  not _27444_ (_02146_, _02081_);
  and _27445_ (_02147_, _01997_, _01954_);
  and _27446_ (_02148_, _02147_, _02006_);
  and _27447_ (_02149_, _02147_, _02012_);
  nor _27448_ (_02150_, _02149_, _02148_);
  and _27449_ (_02151_, _02150_, _02146_);
  not _27450_ (_02152_, _02151_);
  nor _27451_ (_02153_, _02152_, _02145_);
  nor _27452_ (_02154_, _02153_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _27453_ (_02155_, _02154_, _02139_);
  nand _27454_ (_02156_, _02155_, _25365_);
  nor _27455_ (_06146_, _02156_, _02138_);
  and _27456_ (_11184_, _06146_, _02089_);
  and _27457_ (_02157_, _01190_, _00921_);
  and _27458_ (_02158_, _02157_, _00835_);
  and _27459_ (_02159_, _00938_, _00892_);
  not _27460_ (_02160_, _00879_);
  nor _27461_ (_02161_, _02160_, _00906_);
  and _27462_ (_02162_, _02161_, _02159_);
  and _27463_ (_02163_, _02162_, _01406_);
  and _27464_ (_02164_, _02163_, _02158_);
  nor _27465_ (_02165_, _02164_, _00894_);
  not _27466_ (_02166_, _02164_);
  and _27467_ (_02167_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or _27468_ (_02168_, _00545_, _00006_);
  and _27469_ (_02169_, _01039_, _00543_);
  or _27470_ (_02170_, _01170_, _01157_);
  or _27471_ (_02171_, _02170_, _02169_);
  or _27472_ (_02172_, _02171_, _02168_);
  nor _27473_ (_02173_, _02172_, _01315_);
  nor _27474_ (_02174_, _02173_, _00254_);
  not _27475_ (_02175_, _02174_);
  and _27476_ (_02176_, _02175_, _01722_);
  and _27477_ (_02177_, _02176_, _01710_);
  nor _27478_ (_02178_, _02177_, _02166_);
  nor _27479_ (_02179_, _02178_, _02167_);
  and _27480_ (_02180_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _27481_ (_02182_, _02173_, _00233_);
  not _27482_ (_02184_, _02182_);
  and _27483_ (_02186_, _02184_, _01657_);
  and _27484_ (_02188_, _02186_, _01653_);
  and _27485_ (_02190_, _02188_, _01638_);
  nor _27486_ (_02192_, _02190_, _02166_);
  nor _27487_ (_02194_, _02192_, _02180_);
  and _27488_ (_02196_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _27489_ (_02198_, _02173_, _00087_);
  not _27490_ (_02200_, _02198_);
  and _27491_ (_02202_, _02200_, _01575_);
  and _27492_ (_02204_, _02202_, _01563_);
  nor _27493_ (_02206_, _02204_, _02166_);
  nor _27494_ (_02208_, _02206_, _02196_);
  and _27495_ (_02210_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _27496_ (_02212_, _02173_, _00215_);
  not _27497_ (_02214_, _02212_);
  and _27498_ (_02216_, _02214_, _01509_);
  and _27499_ (_02218_, _02216_, _01506_);
  nand _27500_ (_02220_, _02218_, _01497_);
  and _27501_ (_02222_, _02220_, _02164_);
  nor _27502_ (_02224_, _02222_, _02210_);
  and _27503_ (_02226_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _27504_ (_02228_, _02173_, _01433_);
  not _27505_ (_02230_, _02228_);
  and _27506_ (_02232_, _02230_, _01435_);
  and _27507_ (_02234_, _02232_, _01438_);
  nand _27508_ (_02236_, _02234_, _01425_);
  and _27509_ (_02238_, _02236_, _02164_);
  nor _27510_ (_02240_, _02238_, _02226_);
  and _27511_ (_02242_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _27512_ (_02244_, _02173_, _01103_);
  not _27513_ (_02246_, _02244_);
  and _27514_ (_02248_, _02246_, _01368_);
  and _27515_ (_02250_, _02248_, _01365_);
  nand _27516_ (_02251_, _02250_, _01389_);
  and _27517_ (_02252_, _02251_, _02164_);
  nor _27518_ (_02253_, _02252_, _02242_);
  nor _27519_ (_02254_, _02164_, _00853_);
  nor _27520_ (_02255_, _02173_, _00363_);
  not _27521_ (_02256_, _02255_);
  and _27522_ (_02257_, _02256_, _01324_);
  and _27523_ (_02258_, _02257_, _01321_);
  and _27524_ (_02259_, _02258_, _01314_);
  not _27525_ (_02260_, _02259_);
  and _27526_ (_02261_, _02260_, _02164_);
  nor _27527_ (_02262_, _02261_, _02254_);
  and _27528_ (_02263_, _02262_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _27529_ (_02264_, _02263_, _02253_);
  and _27530_ (_02265_, _02264_, _02240_);
  and _27531_ (_02266_, _02265_, _02224_);
  and _27532_ (_02267_, _02266_, _02208_);
  and _27533_ (_02268_, _02267_, _02194_);
  and _27534_ (_02269_, _02268_, _02179_);
  nand _27535_ (_02270_, _02269_, _02165_);
  or _27536_ (_02271_, _02269_, _02165_);
  and _27537_ (_02272_, _02271_, _00866_);
  nand _27538_ (_02273_, _02272_, _02270_);
  nor _27539_ (_02274_, _02164_, _00898_);
  and _27540_ (_02275_, _02274_, _02273_);
  nor _27541_ (_02276_, _02173_, _00285_);
  not _27542_ (_02277_, _02276_);
  and _27543_ (_02278_, _02277_, _01169_);
  and _27544_ (_02279_, _02278_, _01156_);
  and _27545_ (_02280_, _02279_, _01132_);
  and _27546_ (_02281_, _02280_, _02164_);
  nor _27547_ (_02282_, _02281_, _02275_);
  and _27548_ (_11198_, _02282_, _25365_);
  not _27549_ (_02283_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _27550_ (_02284_, _02262_, _02283_);
  nor _27551_ (_02285_, _02262_, _02283_);
  nor _27552_ (_02286_, _02285_, _02284_);
  and _27553_ (_02287_, _02286_, _00866_);
  nor _27554_ (_02288_, _02287_, _00854_);
  nor _27555_ (_02289_, _02288_, _02164_);
  nor _27556_ (_02290_, _02289_, _02261_);
  nand _27557_ (_11985_, _02290_, _25365_);
  nor _27558_ (_02291_, _02263_, _02253_);
  nor _27559_ (_02292_, _02291_, _02264_);
  nor _27560_ (_02293_, _02292_, _00813_);
  nor _27561_ (_02294_, _02293_, _00838_);
  nor _27562_ (_02295_, _02294_, _02164_);
  nor _27563_ (_02296_, _02295_, _02252_);
  nand _27564_ (_11994_, _02296_, _25365_);
  nor _27565_ (_02297_, _02264_, _02240_);
  nor _27566_ (_02298_, _02297_, _02265_);
  nor _27567_ (_02299_, _02298_, _00813_);
  nor _27568_ (_02300_, _02299_, _00818_);
  nor _27569_ (_02301_, _02300_, _02164_);
  nor _27570_ (_02302_, _02301_, _02238_);
  nand _27571_ (_12002_, _02302_, _25365_);
  nor _27572_ (_02303_, _02265_, _02224_);
  nor _27573_ (_02304_, _02303_, _02266_);
  nor _27574_ (_02305_, _02304_, _00813_);
  nor _27575_ (_02306_, _02305_, _00911_);
  nor _27576_ (_02307_, _02306_, _02164_);
  nor _27577_ (_02308_, _02307_, _02222_);
  nor _27578_ (_12009_, _02308_, rst);
  nor _27579_ (_02309_, _02266_, _02208_);
  nor _27580_ (_02310_, _02309_, _02267_);
  nor _27581_ (_02311_, _02310_, _00813_);
  nor _27582_ (_02312_, _02311_, _00931_);
  nor _27583_ (_02313_, _02312_, _02164_);
  nor _27584_ (_02314_, _02313_, _02206_);
  nor _27585_ (_12018_, _02314_, rst);
  nor _27586_ (_02315_, _02267_, _02194_);
  nor _27587_ (_02316_, _02315_, _02268_);
  nor _27588_ (_02317_, _02316_, _00813_);
  nor _27589_ (_02318_, _02317_, _00884_);
  nor _27590_ (_02319_, _02318_, _02164_);
  nor _27591_ (_02320_, _02319_, _02192_);
  nor _27592_ (_12026_, _02320_, rst);
  nor _27593_ (_02321_, _02268_, _02179_);
  nor _27594_ (_02322_, _02321_, _02269_);
  nor _27595_ (_02323_, _02322_, _00813_);
  nor _27596_ (_02324_, _02323_, _00869_);
  nor _27597_ (_02325_, _02324_, _02164_);
  nor _27598_ (_02326_, _02325_, _02178_);
  nor _27599_ (_12034_, _02326_, rst);
  and _27600_ (_02327_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _00000_);
  and _27601_ (_02328_, _02327_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  nor _27602_ (_02329_, _01171_, _00104_);
  nor _27603_ (_02330_, _01265_, _00215_);
  and _27604_ (_02331_, _01003_, _00118_);
  not _27605_ (_02332_, _02331_);
  and _27606_ (_02333_, _01109_, _00388_);
  and _27607_ (_02334_, _02333_, _00197_);
  and _27608_ (_02335_, _02334_, _00146_);
  and _27609_ (_02336_, _02335_, _00954_);
  and _27610_ (_02337_, _02336_, _01087_);
  nor _27611_ (_02338_, _02337_, _01111_);
  and _27612_ (_02339_, _01003_, _00170_);
  nor _27613_ (_02340_, _02339_, _02338_);
  and _27614_ (_02341_, _02340_, _02332_);
  and _27615_ (_02342_, _01117_, _00285_);
  and _27616_ (_02343_, _00132_, _00183_);
  nor _27617_ (_02344_, _00146_, _00197_);
  and _27618_ (_02345_, _02344_, _02343_);
  and _27619_ (_02346_, _02345_, _02342_);
  and _27620_ (_02347_, _00118_, _00170_);
  and _27621_ (_02348_, _02347_, _02346_);
  nor _27622_ (_02349_, _02348_, _01003_);
  not _27623_ (_02350_, _02349_);
  and _27624_ (_02351_, _02350_, _02341_);
  and _27625_ (_02352_, _01003_, _00163_);
  nor _27626_ (_02353_, _02352_, _01699_);
  and _27627_ (_02354_, _02353_, _02351_);
  and _27628_ (_02355_, _02354_, _01124_);
  nor _27629_ (_02356_, _02354_, _01124_);
  nor _27630_ (_02357_, _02356_, _02355_);
  and _27631_ (_02358_, _02357_, _01102_);
  and _27632_ (_02359_, _01003_, _01124_);
  nor _27633_ (_02360_, _02359_, _01215_);
  nor _27634_ (_02361_, _02360_, _01129_);
  or _27635_ (_02362_, _02361_, _02358_);
  or _27636_ (_02363_, _02362_, _02330_);
  and _27637_ (_02364_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor _27638_ (_02365_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _27639_ (_02366_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _27640_ (_02367_, _02366_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27641_ (_02368_, _02367_, _02365_);
  nor _27642_ (_02369_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _27643_ (_02370_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _27644_ (_02371_, _02370_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27645_ (_02372_, _02371_, _02369_);
  nor _27646_ (_02373_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _27647_ (_02374_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _27648_ (_02375_, _02374_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27649_ (_02376_, _02375_, _02373_);
  not _27650_ (_02377_, _02376_);
  nor _27651_ (_02378_, _02377_, _01197_);
  nor _27652_ (_02379_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _27653_ (_02380_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _27654_ (_02381_, _02380_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27655_ (_02382_, _02381_, _02379_);
  and _27656_ (_02383_, _02382_, _02378_);
  nor _27657_ (_02384_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _27658_ (_02385_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _27659_ (_02386_, _02385_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27660_ (_02387_, _02386_, _02384_);
  and _27661_ (_02388_, _02387_, _02383_);
  and _27662_ (_02389_, _02388_, _02372_);
  nor _27663_ (_02390_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _27664_ (_02391_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _27665_ (_02392_, _02391_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27666_ (_02393_, _02392_, _02390_);
  and _27667_ (_02394_, _02393_, _02389_);
  and _27668_ (_02395_, _02394_, _02368_);
  nor _27669_ (_02396_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _27670_ (_02397_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _27671_ (_02398_, _02397_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27672_ (_02399_, _02398_, _02396_);
  and _27673_ (_02400_, _02399_, _02395_);
  nor _27674_ (_02401_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _27675_ (_02402_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _27676_ (_02403_, _02402_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _27677_ (_02404_, _02403_, _02401_);
  nor _27678_ (_02405_, _02404_, _02400_);
  and _27679_ (_02406_, _02404_, _02400_);
  or _27680_ (_02407_, _02406_, _02405_);
  nor _27681_ (_02408_, _02407_, _01041_);
  and _27682_ (_02409_, _00502_, _00006_);
  or _27683_ (_02410_, _02409_, _02408_);
  or _27684_ (_02411_, _02410_, _02364_);
  or _27685_ (_02412_, _02411_, _02363_);
  or _27686_ (_02413_, _02412_, _02329_);
  and _27687_ (_02414_, _02413_, _02328_);
  not _27688_ (_02415_, _02328_);
  and _27689_ (_02416_, _02162_, _01530_);
  and _27690_ (_02417_, _02416_, _02157_);
  or _27691_ (_02418_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _27692_ (_02419_, _02418_, _02415_);
  not _27693_ (_02420_, _02417_);
  or _27694_ (_02421_, _02420_, _01184_);
  and _27695_ (_02422_, _02421_, _02419_);
  or _27696_ (_02423_, _02422_, _02414_);
  and _27697_ (_15457_, _02423_, _25365_);
  and _27698_ (_02424_, _02162_, _01468_);
  and _27699_ (_02425_, _02424_, _02157_);
  nor _27700_ (_02426_, _02425_, _02328_);
  or _27701_ (_02427_, _02426_, _01184_);
  not _27702_ (_02428_, _02426_);
  or _27703_ (_02429_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _27704_ (_02430_, _02429_, _25365_);
  and _27705_ (_15472_, _02430_, _02427_);
  and _27706_ (_02431_, _01170_, _00197_);
  nor _27707_ (_02432_, _01265_, _00087_);
  nor _27708_ (_02433_, _01215_, _01127_);
  not _27709_ (_02434_, _02433_);
  nor _27710_ (_02435_, _02434_, _01119_);
  nor _27711_ (_02436_, _02435_, _00197_);
  and _27712_ (_02437_, _02435_, _00197_);
  nor _27713_ (_02438_, _02437_, _02436_);
  and _27714_ (_02439_, _02438_, _01102_);
  nor _27715_ (_02440_, _01129_, _00363_);
  or _27716_ (_02441_, _02440_, _02439_);
  or _27717_ (_02442_, _02441_, _02432_);
  and _27718_ (_02443_, _00755_, _00545_);
  and _27719_ (_02444_, _02377_, _01197_);
  nor _27720_ (_02445_, _02444_, _02378_);
  and _27721_ (_02446_, _02445_, _01040_);
  and _27722_ (_02447_, _00477_, _00006_);
  or _27723_ (_02448_, _02447_, _02446_);
  or _27724_ (_02449_, _02448_, _02443_);
  or _27725_ (_02450_, _02449_, _02442_);
  or _27726_ (_02451_, _02450_, _02431_);
  and _27727_ (_02452_, _02451_, _02328_);
  or _27728_ (_02453_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _27729_ (_02454_, _02453_, _02415_);
  or _27730_ (_02455_, _02420_, _01337_);
  and _27731_ (_02456_, _02455_, _02454_);
  or _27732_ (_02457_, _02456_, _02452_);
  and _27733_ (_16111_, _02457_, _25365_);
  nor _27734_ (_02458_, _02382_, _02378_);
  nor _27735_ (_02459_, _02458_, _02383_);
  and _27736_ (_02460_, _02459_, _01040_);
  not _27737_ (_02461_, _02460_);
  and _27738_ (_02462_, _00662_, _00545_);
  not _27739_ (_02463_, _02462_);
  and _27740_ (_02464_, _01170_, _00146_);
  nor _27741_ (_02465_, _02334_, _01111_);
  and _27742_ (_02466_, _02342_, _00960_);
  nor _27743_ (_02467_, _02466_, _01003_);
  or _27744_ (_02468_, _02467_, _02465_);
  nor _27745_ (_02469_, _02468_, _00571_);
  and _27746_ (_02470_, _02468_, _00571_);
  or _27747_ (_02471_, _02470_, _01559_);
  nor _27748_ (_02472_, _02471_, _02469_);
  and _27749_ (_02473_, _00479_, _00006_);
  nor _27750_ (_02474_, _01265_, _00233_);
  and _27751_ (_02475_, _01128_, _00312_);
  or _27752_ (_02476_, _02475_, _02474_);
  or _27753_ (_02477_, _02476_, _02473_);
  or _27754_ (_02478_, _02477_, _02472_);
  nor _27755_ (_02479_, _02478_, _02464_);
  and _27756_ (_02480_, _02479_, _02463_);
  and _27757_ (_02481_, _02480_, _02461_);
  nor _27758_ (_02482_, _02481_, _02415_);
  or _27759_ (_02483_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _27760_ (_02484_, _02483_, _02415_);
  or _27761_ (_02485_, _02420_, _01397_);
  and _27762_ (_02486_, _02485_, _02484_);
  or _27763_ (_02487_, _02486_, _02482_);
  and _27764_ (_16119_, _02487_, _25365_);
  nor _27765_ (_02488_, _02387_, _02383_);
  nor _27766_ (_02489_, _02488_, _02388_);
  and _27767_ (_02490_, _02489_, _01040_);
  not _27768_ (_02491_, _02490_);
  and _27769_ (_02492_, _02466_, _00571_);
  and _27770_ (_02493_, _02492_, _01111_);
  and _27771_ (_02494_, _02335_, _01003_);
  nor _27772_ (_02495_, _02494_, _02493_);
  and _27773_ (_02496_, _02495_, _00183_);
  nor _27774_ (_02497_, _02495_, _00183_);
  nor _27775_ (_02498_, _02497_, _02496_);
  and _27776_ (_02499_, _02498_, _01102_);
  and _27777_ (_02500_, _01128_, _00327_);
  and _27778_ (_02501_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _27779_ (_02502_, _02501_, _02500_);
  and _27780_ (_02503_, _00481_, _00006_);
  nor _27781_ (_02504_, _01265_, _00254_);
  nor _27782_ (_02505_, _01171_, _00183_);
  or _27783_ (_02506_, _02505_, _02504_);
  nor _27784_ (_02507_, _02506_, _02503_);
  and _27785_ (_02508_, _02507_, _02502_);
  not _27786_ (_02509_, _02508_);
  nor _27787_ (_02510_, _02509_, _02499_);
  and _27788_ (_02511_, _02510_, _02491_);
  nor _27789_ (_02512_, _02511_, _02415_);
  or _27790_ (_02513_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _27791_ (_02514_, _02513_, _02415_);
  or _27792_ (_02515_, _02420_, _01457_);
  and _27793_ (_02516_, _02515_, _02514_);
  or _27794_ (_02517_, _02516_, _02512_);
  and _27795_ (_16127_, _02517_, _25365_);
  nor _27796_ (_02518_, _02388_, _02372_);
  nor _27797_ (_02519_, _02518_, _02389_);
  and _27798_ (_02520_, _02519_, _01040_);
  not _27799_ (_02521_, _02520_);
  nor _27800_ (_02522_, _02336_, _01087_);
  not _27801_ (_02523_, _02522_);
  and _27802_ (_02524_, _02523_, _02338_);
  and _27803_ (_02525_, _02492_, _00183_);
  nor _27804_ (_02526_, _02525_, _00132_);
  nor _27805_ (_02527_, _02526_, _02346_);
  nor _27806_ (_02528_, _02527_, _01003_);
  nor _27807_ (_02529_, _02528_, _02524_);
  nor _27808_ (_02530_, _02529_, _01559_);
  nor _27809_ (_02531_, _01171_, _00132_);
  or _27810_ (_02532_, _02531_, _01267_);
  nor _27811_ (_02533_, _02532_, _02530_);
  and _27812_ (_02534_, _00484_, _00006_);
  nor _27813_ (_02535_, _01129_, _00215_);
  and _27814_ (_02536_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _27815_ (_02537_, _02536_, _02535_);
  nor _27816_ (_02538_, _02537_, _02534_);
  and _27817_ (_02539_, _02538_, _02533_);
  and _27818_ (_02540_, _02539_, _02521_);
  nor _27819_ (_02541_, _02540_, _02415_);
  or _27820_ (_02542_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _27821_ (_02543_, _02542_, _02415_);
  or _27822_ (_02544_, _02420_, _01522_);
  and _27823_ (_02545_, _02544_, _02543_);
  or _27824_ (_02546_, _02545_, _02541_);
  and _27825_ (_16135_, _02546_, _25365_);
  nor _27826_ (_02547_, _02393_, _02389_);
  not _27827_ (_02548_, _02547_);
  nor _27828_ (_02549_, _02394_, _01041_);
  and _27829_ (_02550_, _02549_, _02548_);
  not _27830_ (_02551_, _02550_);
  and _27831_ (_02552_, _00487_, _00006_);
  not _27832_ (_02553_, _02552_);
  nor _27833_ (_02554_, _02346_, _01003_);
  nor _27834_ (_02555_, _02554_, _02338_);
  nor _27835_ (_02556_, _02555_, _01053_);
  and _27836_ (_02557_, _02555_, _01053_);
  nor _27837_ (_02558_, _02557_, _02556_);
  and _27838_ (_02559_, _02558_, _01102_);
  and _27839_ (_02560_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _27840_ (_02561_, _01003_, _00088_);
  or _27841_ (_02562_, _02561_, _01129_);
  nor _27842_ (_02563_, _02562_, _02339_);
  nor _27843_ (_02564_, _01265_, _00363_);
  nor _27844_ (_02565_, _01171_, _00170_);
  or _27845_ (_02566_, _02565_, _02564_);
  or _27846_ (_02567_, _02566_, _02563_);
  nor _27847_ (_02568_, _02567_, _02560_);
  not _27848_ (_02569_, _02568_);
  nor _27849_ (_02570_, _02569_, _02559_);
  and _27850_ (_02571_, _02570_, _02553_);
  and _27851_ (_02572_, _02571_, _02551_);
  nor _27852_ (_02573_, _02572_, _02415_);
  or _27853_ (_02574_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _27854_ (_02575_, _02574_, _02415_);
  or _27855_ (_02576_, _02420_, _01589_);
  and _27856_ (_02577_, _02576_, _02575_);
  or _27857_ (_02578_, _02577_, _02573_);
  and _27858_ (_16143_, _02578_, _25365_);
  nor _27859_ (_02579_, _02394_, _02368_);
  nor _27860_ (_02580_, _02579_, _02395_);
  and _27861_ (_02581_, _02580_, _01040_);
  not _27862_ (_02582_, _02581_);
  and _27863_ (_02583_, _00492_, _00006_);
  and _27864_ (_02584_, _02346_, _00170_);
  nor _27865_ (_02585_, _02584_, _01003_);
  not _27866_ (_02586_, _02585_);
  and _27867_ (_02587_, _02586_, _02340_);
  and _27868_ (_02588_, _02587_, _00118_);
  nor _27869_ (_02589_, _02587_, _00118_);
  nor _27870_ (_02590_, _02589_, _02588_);
  nor _27871_ (_02591_, _02590_, _01559_);
  and _27872_ (_02592_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _27873_ (_02593_, _01702_, _01129_);
  and _27874_ (_02594_, _02593_, _02332_);
  and _27875_ (_02595_, _01263_, _00312_);
  nor _27876_ (_02596_, _01171_, _00118_);
  or _27877_ (_02597_, _02596_, _02595_);
  or _27878_ (_02598_, _02597_, _02594_);
  nor _27879_ (_02599_, _02598_, _02592_);
  not _27880_ (_02600_, _02599_);
  nor _27881_ (_02601_, _02600_, _02591_);
  not _27882_ (_02602_, _02601_);
  nor _27883_ (_02603_, _02602_, _02583_);
  and _27884_ (_02604_, _02603_, _02582_);
  nor _27885_ (_02605_, _02604_, _02415_);
  or _27886_ (_02606_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _27887_ (_02607_, _02606_, _02415_);
  or _27888_ (_02608_, _02420_, _01673_);
  and _27889_ (_02609_, _02608_, _02607_);
  or _27890_ (_02610_, _02609_, _02605_);
  and _27891_ (_16150_, _02610_, _25365_);
  nor _27892_ (_02611_, _02399_, _02395_);
  not _27893_ (_02612_, _02611_);
  nor _27894_ (_02613_, _02400_, _01041_);
  and _27895_ (_02614_, _02613_, _02612_);
  not _27896_ (_02615_, _02614_);
  and _27897_ (_02616_, _00497_, _00006_);
  nor _27898_ (_02617_, _02351_, _00163_);
  and _27899_ (_02618_, _02351_, _00163_);
  nor _27900_ (_02619_, _02618_, _02617_);
  nor _27901_ (_02620_, _02619_, _01559_);
  and _27902_ (_02621_, _00545_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _27903_ (_02622_, _01003_, _00256_);
  or _27904_ (_02623_, _02622_, _01129_);
  nor _27905_ (_02624_, _02623_, _02352_);
  and _27906_ (_02625_, _01263_, _00327_);
  nor _27907_ (_02626_, _01171_, _00163_);
  or _27908_ (_02627_, _02626_, _02625_);
  or _27909_ (_02628_, _02627_, _02624_);
  nor _27910_ (_02629_, _02628_, _02621_);
  not _27911_ (_02630_, _02629_);
  nor _27912_ (_02631_, _02630_, _02620_);
  not _27913_ (_02632_, _02631_);
  nor _27914_ (_02633_, _02632_, _02616_);
  and _27915_ (_02634_, _02633_, _02615_);
  nor _27916_ (_02635_, _02634_, _02415_);
  or _27917_ (_02636_, _02417_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _27918_ (_02637_, _02636_, _02415_);
  or _27919_ (_02638_, _02420_, _01737_);
  and _27920_ (_02639_, _02638_, _02637_);
  or _27921_ (_02640_, _02639_, _02635_);
  and _27922_ (_16159_, _02640_, _25365_);
  or _27923_ (_02641_, _02426_, _01337_);
  or _27924_ (_02642_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _27925_ (_02643_, _02642_, _25365_);
  and _27926_ (_16166_, _02643_, _02641_);
  or _27927_ (_02644_, _02426_, _01397_);
  or _27928_ (_02645_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _27929_ (_02646_, _02645_, _25365_);
  and _27930_ (_16175_, _02646_, _02644_);
  or _27931_ (_02647_, _02426_, _01457_);
  or _27932_ (_02648_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _27933_ (_02649_, _02648_, _25365_);
  and _27934_ (_16182_, _02649_, _02647_);
  or _27935_ (_02650_, _02426_, _01522_);
  or _27936_ (_02651_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _27937_ (_02652_, _02651_, _25365_);
  and _27938_ (_16190_, _02652_, _02650_);
  or _27939_ (_02653_, _02426_, _01589_);
  or _27940_ (_02654_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _27941_ (_02655_, _02654_, _25365_);
  and _27942_ (_16198_, _02655_, _02653_);
  or _27943_ (_02656_, _02426_, _01673_);
  or _27944_ (_02657_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _27945_ (_02658_, _02657_, _25365_);
  and _27946_ (_16206_, _02658_, _02656_);
  or _27947_ (_02660_, _02426_, _01737_);
  or _27948_ (_02661_, _02428_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _27949_ (_02662_, _02661_, _25365_);
  and _27950_ (_16214_, _02662_, _02660_);
  not _27951_ (_02663_, _00892_);
  nor _27952_ (_02664_, _02663_, _00879_);
  and _27953_ (_02665_, _02664_, _01298_);
  and _27954_ (_02666_, _02665_, _00940_);
  not _27955_ (_02667_, _01294_);
  nor _27956_ (_02669_, _02667_, _01289_);
  not _27957_ (_02670_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _27958_ (_02671_, _01294_, _02670_);
  or _27959_ (_02672_, _02671_, _02669_);
  and _27960_ (_02673_, _02672_, _02666_);
  nor _27961_ (_02674_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _27962_ (_02675_, _02674_);
  nand _27963_ (_02676_, _02675_, _01289_);
  and _27964_ (_02677_, _02674_, _02670_);
  nor _27965_ (_02678_, _02677_, _02666_);
  and _27966_ (_02679_, _02678_, _02676_);
  nor _27967_ (_02680_, _00938_, _02663_);
  nor _27968_ (_02681_, _00879_, _00906_);
  and _27969_ (_02682_, _02157_, _00860_);
  and _27970_ (_02683_, _02682_, _02681_);
  and _27971_ (_02684_, _02683_, _02680_);
  or _27972_ (_02685_, _02684_, _02679_);
  or _27973_ (_02686_, _02685_, _02673_);
  nand _27974_ (_02687_, _02684_, _02280_);
  and _27975_ (_02688_, _02687_, _25365_);
  and _27976_ (_17600_, _02688_, _02686_);
  and _27977_ (_02689_, _01406_, _00835_);
  and _27978_ (_02690_, _02666_, _02689_);
  nand _27979_ (_02691_, _02690_, _01289_);
  not _27980_ (_02692_, _02684_);
  or _27981_ (_02693_, _02690_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _27982_ (_02694_, _02693_, _02692_);
  and _27983_ (_02695_, _02694_, _02691_);
  and _27984_ (_02696_, _02684_, _02251_);
  or _27985_ (_02697_, _02696_, _02695_);
  and _27986_ (_19908_, _02697_, _25365_);
  or _27987_ (_02698_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _27988_ (_02699_, _00518_, _00510_);
  or _27989_ (_02700_, _02699_, _00524_);
  or _27990_ (_02701_, _02700_, _00529_);
  or _27991_ (_02702_, _00538_, _00534_);
  or _27992_ (_02703_, _00540_, _00473_);
  or _27993_ (_02704_, _02703_, _02702_);
  or _27994_ (_02705_, _02704_, _02701_);
  and _27995_ (_02706_, _02705_, _00006_);
  or _27996_ (_02707_, _01205_, _01096_);
  not _27997_ (_02708_, _01203_);
  nand _27998_ (_02709_, _02708_, _01096_);
  and _27999_ (_02710_, _02709_, _01047_);
  and _28000_ (_02711_, _02710_, _02707_);
  not _28001_ (_02712_, _01032_);
  nand _28002_ (_02713_, _01031_, _02712_);
  or _28003_ (_02714_, _01033_, _01031_);
  and _28004_ (_02715_, _01040_, _02714_);
  and _28005_ (_02716_, _02715_, _02713_);
  and _28006_ (_02717_, _02347_, _00654_);
  and _28007_ (_02718_, _02345_, _00545_);
  nand _28008_ (_02719_, _02718_, _02717_);
  nand _28009_ (_02720_, _02719_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _28010_ (_02721_, _02720_, _02716_);
  or _28011_ (_02722_, _02721_, _02711_);
  or _28012_ (_02723_, _02722_, _02706_);
  and _28013_ (_02724_, _02723_, _02698_);
  or _28014_ (_02725_, _02724_, _02666_);
  not _28015_ (_02726_, _02666_);
  and _28016_ (_02727_, _01469_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _28017_ (_02728_, _02727_, _01470_);
  or _28018_ (_02729_, _02728_, _02726_);
  and _28019_ (_02730_, _02729_, _02725_);
  or _28020_ (_02731_, _02730_, _02684_);
  or _28021_ (_02732_, _02692_, _02236_);
  and _28022_ (_02733_, _02732_, _25365_);
  and _28023_ (_19919_, _02733_, _02731_);
  and _28024_ (_02735_, _02666_, _01530_);
  nand _28025_ (_02736_, _02735_, _01289_);
  or _28026_ (_02737_, _02735_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _28027_ (_02738_, _02737_, _02692_);
  and _28028_ (_02739_, _02738_, _02736_);
  and _28029_ (_02740_, _02684_, _02220_);
  or _28030_ (_02741_, _02740_, _02739_);
  and _28031_ (_19930_, _02741_, _25365_);
  or _28032_ (_02742_, _02726_, _01599_);
  and _28033_ (_02743_, _02680_, _02681_);
  and _28034_ (_02744_, _02743_, _02682_);
  not _28035_ (_02745_, _02744_);
  and _28036_ (_02746_, _02745_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _28037_ (_02747_, _02745_, _02204_);
  nor _28038_ (_02748_, _02747_, _02746_);
  nor _28039_ (_06114_, _02748_, rst);
  and _28040_ (_02749_, _06114_, _02742_);
  and _28041_ (_02750_, _01598_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _28042_ (_02751_, _02750_, _01602_);
  nor _28043_ (_02752_, _02684_, rst);
  and _28044_ (_02753_, _02752_, _02666_);
  and _28045_ (_02754_, _02753_, _02751_);
  or _28046_ (_19941_, _02754_, _02749_);
  and _28047_ (_02755_, _02666_, _01680_);
  nand _28048_ (_02756_, _02755_, _01289_);
  or _28049_ (_02757_, _02755_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _28050_ (_02758_, _02757_, _02692_);
  and _28051_ (_02759_, _02758_, _02756_);
  nor _28052_ (_02760_, _02692_, _02190_);
  or _28053_ (_02761_, _02760_, _02759_);
  and _28054_ (_19952_, _02761_, _25365_);
  and _28055_ (_02762_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _28056_ (_02763_, _02762_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _28057_ (_02764_, _01092_, _01047_);
  and _28058_ (_02765_, _01040_, _01016_);
  nand _28059_ (_02766_, _01170_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _28060_ (_02767_, _02766_, _02762_);
  or _28061_ (_02768_, _02767_, _02765_);
  or _28062_ (_02769_, _02768_, _02764_);
  and _28063_ (_02770_, _02769_, _02763_);
  or _28064_ (_02771_, _02770_, _02666_);
  not _28065_ (_02772_, _01745_);
  nor _28066_ (_02773_, _02772_, _01289_);
  or _28067_ (_02774_, _01745_, _01498_);
  nand _28068_ (_02775_, _02774_, _02666_);
  or _28069_ (_02776_, _02775_, _02773_);
  and _28070_ (_02777_, _02776_, _02771_);
  or _28071_ (_02778_, _02777_, _02684_);
  nand _28072_ (_02779_, _02684_, _02177_);
  and _28073_ (_02780_, _02779_, _25365_);
  and _28074_ (_19963_, _02780_, _02778_);
  nor _28075_ (_02781_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _28076_ (_02782_, _02781_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _28077_ (_02783_, _00860_, _00921_);
  and _28078_ (_02784_, _00938_, _02663_);
  and _28079_ (_02785_, _02784_, _02681_);
  and _28080_ (_02786_, _02785_, _02783_);
  and _28081_ (_02787_, _02786_, _01190_);
  nor _28082_ (_02788_, _02787_, _02782_);
  not _28083_ (_02789_, _02788_);
  nand _28084_ (_02790_, _02789_, _01184_);
  not _28085_ (_02791_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _28086_ (_02792_, _02327_, _02791_);
  and _28087_ (_02793_, _00938_, _00921_);
  and _28088_ (_02794_, _02793_, _00893_);
  not _28089_ (_02795_, _01298_);
  nor _28090_ (_02796_, _02795_, _00906_);
  and _28091_ (_02797_, _02796_, _02794_);
  and _28092_ (_02798_, _02797_, _01294_);
  and _28093_ (_02799_, _02798_, _01289_);
  nor _28094_ (_02800_, _02798_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _28095_ (_02801_, _02800_);
  not _28096_ (_02802_, _02792_);
  and _28097_ (_02803_, _02802_, _02788_);
  and _28098_ (_02804_, _02803_, _02801_);
  not _28099_ (_02805_, _02804_);
  nor _28100_ (_02806_, _02805_, _02799_);
  nor _28101_ (_02807_, _02806_, _02792_);
  nand _28102_ (_02808_, _02807_, _02790_);
  or _28103_ (_02809_, _02802_, _02413_);
  and _28104_ (_02810_, _02809_, _02808_);
  and _28105_ (_20533_, _02810_, _25365_);
  nand _28106_ (_02811_, _02789_, _01337_);
  and _28107_ (_02812_, _02797_, _00860_);
  and _28108_ (_02813_, _02812_, _01289_);
  nor _28109_ (_02814_, _02812_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not _28110_ (_02815_, _02814_);
  and _28111_ (_02816_, _02815_, _02803_);
  not _28112_ (_02817_, _02816_);
  nor _28113_ (_02818_, _02817_, _02813_);
  nor _28114_ (_02819_, _02818_, _02792_);
  nand _28115_ (_02820_, _02819_, _02811_);
  or _28116_ (_02821_, _02802_, _02451_);
  and _28117_ (_02822_, _02821_, _02820_);
  and _28118_ (_22204_, _02822_, _25365_);
  and _28119_ (_02823_, _02792_, _02481_);
  not _28120_ (_02824_, _02823_);
  nand _28121_ (_02825_, _02789_, _01397_);
  and _28122_ (_02826_, _02797_, _02689_);
  and _28123_ (_02827_, _02826_, _01289_);
  nor _28124_ (_02828_, _02826_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not _28125_ (_02829_, _02828_);
  and _28126_ (_02830_, _02829_, _02803_);
  not _28127_ (_02831_, _02830_);
  nor _28128_ (_02832_, _02831_, _02827_);
  nor _28129_ (_02833_, _02832_, _02792_);
  nand _28130_ (_02834_, _02833_, _02825_);
  and _28131_ (_02835_, _02834_, _02824_);
  and _28132_ (_22213_, _02835_, _25365_);
  nand _28133_ (_02836_, _02789_, _01457_);
  and _28134_ (_02837_, _02797_, _01468_);
  and _28135_ (_02838_, _02837_, _01289_);
  nor _28136_ (_02839_, _02837_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _28137_ (_02840_, _02839_);
  and _28138_ (_02841_, _02840_, _02803_);
  not _28139_ (_02842_, _02841_);
  nor _28140_ (_02843_, _02842_, _02838_);
  nor _28141_ (_02844_, _02843_, _02792_);
  nand _28142_ (_02845_, _02844_, _02836_);
  and _28143_ (_02846_, _02792_, _02511_);
  not _28144_ (_02847_, _02846_);
  and _28145_ (_02848_, _02847_, _02845_);
  and _28146_ (_22214_, _02848_, _25365_);
  nand _28147_ (_02849_, _02789_, _01522_);
  not _28148_ (_02850_, _02797_);
  and _28149_ (_02851_, _02803_, _02850_);
  and _28150_ (_02852_, _02851_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _28151_ (_02853_, _01530_, _00129_);
  nor _28152_ (_02854_, _02853_, _01531_);
  and _28153_ (_02855_, _02797_, _02802_);
  not _28154_ (_02856_, _02855_);
  nor _28155_ (_02857_, _02856_, _02854_);
  and _28156_ (_02858_, _02857_, _02803_);
  nor _28157_ (_02859_, _02858_, _02852_);
  and _28158_ (_02860_, _02859_, _02802_);
  and _28159_ (_02861_, _02860_, _02849_);
  and _28160_ (_02862_, _02792_, _02540_);
  nor _28161_ (_02863_, _02862_, _02861_);
  and _28162_ (_22222_, _02863_, _25365_);
  nand _28163_ (_02864_, _02789_, _01589_);
  and _28164_ (_02865_, _02797_, _01597_);
  and _28165_ (_02866_, _02865_, _01289_);
  nor _28166_ (_02867_, _02865_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not _28167_ (_02868_, _02867_);
  and _28168_ (_02869_, _02868_, _02803_);
  not _28169_ (_02870_, _02869_);
  nor _28170_ (_02871_, _02870_, _02866_);
  nor _28171_ (_02872_, _02871_, _02792_);
  nand _28172_ (_02873_, _02872_, _02864_);
  and _28173_ (_02874_, _02792_, _02572_);
  not _28174_ (_02875_, _02874_);
  and _28175_ (_02876_, _02875_, _02873_);
  and _28176_ (_22233_, _02876_, _25365_);
  nand _28177_ (_02877_, _02789_, _01673_);
  and _28178_ (_02878_, _02797_, _01680_);
  and _28179_ (_02879_, _02878_, _01289_);
  nor _28180_ (_02880_, _02878_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not _28181_ (_02881_, _02880_);
  and _28182_ (_02882_, _02881_, _02803_);
  not _28183_ (_02883_, _02882_);
  nor _28184_ (_02884_, _02883_, _02879_);
  nor _28185_ (_02885_, _02884_, _02792_);
  nand _28186_ (_02886_, _02885_, _02877_);
  and _28187_ (_02887_, _02792_, _02604_);
  not _28188_ (_02888_, _02887_);
  and _28189_ (_02889_, _02888_, _02886_);
  and _28190_ (_22243_, _02889_, _25365_);
  nand _28191_ (_02890_, _02789_, _01737_);
  and _28192_ (_02891_, _02797_, _01745_);
  and _28193_ (_02892_, _02891_, _01289_);
  nor _28194_ (_02893_, _02891_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not _28195_ (_02894_, _02893_);
  and _28196_ (_02895_, _02894_, _02803_);
  not _28197_ (_02896_, _02895_);
  nor _28198_ (_02897_, _02896_, _02892_);
  nor _28199_ (_02898_, _02897_, _02792_);
  nand _28200_ (_02899_, _02898_, _02890_);
  and _28201_ (_02900_, _02792_, _02634_);
  not _28202_ (_02901_, _02900_);
  and _28203_ (_02902_, _02901_, _02899_);
  and _28204_ (_22254_, _02902_, _25365_);
  and _28205_ (_02903_, _00892_, _00879_);
  and _28206_ (_02904_, _02793_, _00907_);
  and _28207_ (_02905_, _02904_, _02903_);
  and _28208_ (_02906_, _02905_, _01294_);
  nand _28209_ (_02907_, _02906_, _01289_);
  or _28210_ (_02908_, _02906_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _28211_ (_02909_, _02908_, _01298_);
  and _28212_ (_02910_, _02909_, _02907_);
  and _28213_ (_02911_, _02162_, _02783_);
  nand _28214_ (_02912_, _02911_, _02280_);
  or _28215_ (_02913_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _28216_ (_02914_, _02913_, _01190_);
  and _28217_ (_02915_, _02914_, _02912_);
  not _28218_ (_02916_, _01189_);
  and _28219_ (_02917_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _28220_ (_02918_, _02917_, rst);
  or _28221_ (_02919_, _02918_, _02915_);
  or _28222_ (_25274_, _02919_, _02910_);
  and _28223_ (_02920_, _02903_, _00940_);
  and _28224_ (_02922_, _02920_, _01294_);
  nand _28225_ (_02923_, _02922_, _01289_);
  or _28226_ (_02924_, _02922_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _28227_ (_02925_, _02924_, _01298_);
  and _28228_ (_02926_, _02925_, _02923_);
  and _28229_ (_02927_, _02680_, _02161_);
  and _28230_ (_02928_, _02927_, _02783_);
  nand _28231_ (_02929_, _02928_, _02280_);
  or _28232_ (_02930_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _28233_ (_02931_, _02930_, _01190_);
  and _28234_ (_02932_, _02931_, _02929_);
  and _28235_ (_02933_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _28236_ (_02934_, _02933_, rst);
  or _28237_ (_02935_, _02934_, _02932_);
  or _28238_ (_25275_, _02935_, _02926_);
  and _28239_ (_02936_, _02663_, _00879_);
  and _28240_ (_02937_, _02936_, _02904_);
  and _28241_ (_02938_, _02937_, _01294_);
  nand _28242_ (_02939_, _02938_, _01289_);
  or _28243_ (_02940_, _02938_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _28244_ (_02941_, _02940_, _01298_);
  and _28245_ (_02942_, _02941_, _02939_);
  and _28246_ (_02943_, _02784_, _02161_);
  and _28247_ (_02944_, _02943_, _02783_);
  not _28248_ (_02945_, _02944_);
  nor _28249_ (_02946_, _02945_, _02280_);
  and _28250_ (_02947_, _02945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _28251_ (_02948_, _02947_, _02946_);
  and _28252_ (_02949_, _02948_, _01190_);
  and _28253_ (_02950_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _28254_ (_02951_, _02950_, rst);
  or _28255_ (_02952_, _02951_, _02949_);
  or _28256_ (_25276_, _02952_, _02942_);
  and _28257_ (_02953_, _02936_, _00940_);
  and _28258_ (_02954_, _02953_, _01294_);
  nand _28259_ (_02955_, _02954_, _01289_);
  or _28260_ (_02956_, _02954_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _28261_ (_02957_, _02956_, _01298_);
  and _28262_ (_02958_, _02957_, _02955_);
  nor _28263_ (_02959_, _00938_, _00892_);
  and _28264_ (_02960_, _02161_, _02959_);
  and _28265_ (_02961_, _02960_, _02783_);
  not _28266_ (_02962_, _02961_);
  nor _28267_ (_02963_, _02962_, _02280_);
  and _28268_ (_02964_, _02962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _28269_ (_02965_, _02964_, _02963_);
  and _28270_ (_02966_, _02965_, _01190_);
  and _28271_ (_02967_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _28272_ (_02968_, _02967_, rst);
  or _28273_ (_02969_, _02968_, _02966_);
  or _28274_ (_25277_, _02969_, _02958_);
  or _28275_ (_02970_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _28276_ (_02971_, _02970_, _01298_);
  nand _28277_ (_02972_, _02911_, _01289_);
  and _28278_ (_02973_, _02972_, _02971_);
  nand _28279_ (_02974_, _02911_, _02259_);
  and _28280_ (_02975_, _02974_, _01190_);
  and _28281_ (_02976_, _02975_, _02970_);
  not _28282_ (_02977_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _28283_ (_02978_, _01189_, _02977_);
  or _28284_ (_02980_, _02978_, rst);
  or _28285_ (_02981_, _02980_, _02976_);
  or _28286_ (_25278_, _02981_, _02973_);
  and _28287_ (_02982_, _02689_, _00921_);
  and _28288_ (_02983_, _02982_, _02162_);
  nand _28289_ (_02984_, _02983_, _01289_);
  or _28290_ (_02985_, _02983_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _28291_ (_02986_, _02985_, _01298_);
  and _28292_ (_02987_, _02986_, _02984_);
  not _28293_ (_02988_, _02911_);
  or _28294_ (_02990_, _02988_, _02251_);
  or _28295_ (_02991_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _28296_ (_02992_, _02991_, _01190_);
  and _28297_ (_02993_, _02992_, _02990_);
  not _28298_ (_02994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor _28299_ (_02995_, _01189_, _02994_);
  or _28300_ (_02996_, _02995_, rst);
  or _28301_ (_02997_, _02996_, _02993_);
  or _28302_ (_25279_, _02997_, _02987_);
  not _28303_ (_02998_, _01532_);
  nand _28304_ (_02999_, _02905_, _02998_);
  and _28305_ (_03000_, _02999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _28306_ (_03001_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _28307_ (_03002_, _03001_, _01470_);
  and _28308_ (_03003_, _03002_, _02905_);
  or _28309_ (_03004_, _03003_, _03000_);
  and _28310_ (_03005_, _03004_, _01298_);
  or _28311_ (_03006_, _02988_, _02236_);
  or _28312_ (_03007_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _28313_ (_03008_, _03007_, _01190_);
  and _28314_ (_03010_, _03008_, _03006_);
  and _28315_ (_03011_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _28316_ (_03012_, _03011_, rst);
  or _28317_ (_03013_, _03012_, _03010_);
  or _28318_ (_25280_, _03013_, _03005_);
  nand _28319_ (_03014_, _02905_, _00835_);
  and _28320_ (_03015_, _03014_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _28321_ (_03016_, _02998_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _28322_ (_03017_, _03016_, _01531_);
  and _28323_ (_03018_, _03017_, _02905_);
  or _28324_ (_03019_, _03018_, _03015_);
  and _28325_ (_03020_, _03019_, _01298_);
  or _28326_ (_03021_, _02988_, _02220_);
  or _28327_ (_03022_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _28328_ (_03023_, _03022_, _01190_);
  and _28329_ (_03024_, _03023_, _03021_);
  and _28330_ (_03025_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _28331_ (_03026_, _03025_, rst);
  or _28332_ (_03027_, _03026_, _03024_);
  or _28333_ (_25281_, _03027_, _03020_);
  not _28334_ (_03029_, _02905_);
  or _28335_ (_03030_, _03029_, _01599_);
  and _28336_ (_03031_, _03030_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _28337_ (_03032_, _01598_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _28338_ (_03033_, _03032_, _01602_);
  and _28339_ (_03034_, _03033_, _02905_);
  or _28340_ (_03035_, _03034_, _03031_);
  and _28341_ (_03036_, _03035_, _01298_);
  nand _28342_ (_03037_, _02911_, _02204_);
  or _28343_ (_03038_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _28344_ (_03039_, _03038_, _01190_);
  and _28345_ (_03040_, _03039_, _03037_);
  and _28346_ (_03041_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _28347_ (_03042_, _03041_, rst);
  or _28348_ (_03043_, _03042_, _03040_);
  or _28349_ (_25282_, _03043_, _03036_);
  and _28350_ (_03044_, _02905_, _01680_);
  nand _28351_ (_03045_, _03044_, _01289_);
  or _28352_ (_03046_, _03044_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _28353_ (_03047_, _03046_, _01298_);
  and _28354_ (_03049_, _03047_, _03045_);
  nand _28355_ (_03050_, _02911_, _02190_);
  or _28356_ (_03051_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _28357_ (_03052_, _03051_, _01190_);
  and _28358_ (_03053_, _03052_, _03050_);
  and _28359_ (_03054_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _28360_ (_03055_, _03054_, rst);
  or _28361_ (_03056_, _03055_, _03053_);
  or _28362_ (_25283_, _03056_, _03049_);
  and _28363_ (_03057_, _02905_, _01745_);
  nand _28364_ (_03059_, _03057_, _01289_);
  or _28365_ (_03060_, _03057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _28366_ (_03061_, _03060_, _01298_);
  and _28367_ (_03062_, _03061_, _03059_);
  nand _28368_ (_03063_, _02911_, _02177_);
  or _28369_ (_03064_, _02911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _28370_ (_03065_, _03064_, _01190_);
  and _28371_ (_03066_, _03065_, _03063_);
  not _28372_ (_03067_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _28373_ (_03068_, _01189_, _03067_);
  or _28374_ (_03070_, _03068_, rst);
  or _28375_ (_03071_, _03070_, _03066_);
  or _28376_ (_25284_, _03071_, _03062_);
  and _28377_ (_03072_, _02920_, _00860_);
  nand _28378_ (_03073_, _03072_, _01289_);
  or _28379_ (_03074_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _28380_ (_03075_, _03074_, _01298_);
  and _28381_ (_03076_, _03075_, _03073_);
  nand _28382_ (_03077_, _02928_, _02259_);
  and _28383_ (_03078_, _03077_, _01190_);
  and _28384_ (_03080_, _03078_, _03074_);
  not _28385_ (_03081_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _28386_ (_03082_, _01189_, _03081_);
  or _28387_ (_03083_, _03082_, rst);
  or _28388_ (_03084_, _03083_, _03080_);
  or _28389_ (_25285_, _03084_, _03076_);
  and _28390_ (_03085_, _02920_, _02689_);
  nand _28391_ (_03086_, _03085_, _01289_);
  or _28392_ (_03087_, _03085_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _28393_ (_03088_, _03087_, _01298_);
  and _28394_ (_03090_, _03088_, _03086_);
  not _28395_ (_03091_, _02928_);
  or _28396_ (_03092_, _03091_, _02251_);
  or _28397_ (_03093_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _28398_ (_03094_, _03093_, _01190_);
  and _28399_ (_03095_, _03094_, _03092_);
  not _28400_ (_03096_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor _28401_ (_03097_, _01189_, _03096_);
  or _28402_ (_03098_, _03097_, rst);
  or _28403_ (_03099_, _03098_, _03095_);
  or _28404_ (_25286_, _03099_, _03090_);
  and _28405_ (_03101_, _02920_, _01468_);
  nand _28406_ (_03102_, _03101_, _01289_);
  or _28407_ (_03103_, _03101_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _28408_ (_03104_, _03103_, _01298_);
  and _28409_ (_03105_, _03104_, _03102_);
  or _28410_ (_03106_, _03091_, _02236_);
  or _28411_ (_03107_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _28412_ (_03108_, _03107_, _01190_);
  and _28413_ (_03109_, _03108_, _03106_);
  and _28414_ (_03111_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _28415_ (_03112_, _03111_, rst);
  or _28416_ (_03113_, _03112_, _03109_);
  or _28417_ (_25287_, _03113_, _03105_);
  and _28418_ (_03114_, _02920_, _01530_);
  nand _28419_ (_03115_, _03114_, _01289_);
  or _28420_ (_03116_, _03114_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _28421_ (_03117_, _03116_, _01298_);
  and _28422_ (_03118_, _03117_, _03115_);
  or _28423_ (_03119_, _03091_, _02220_);
  or _28424_ (_03122_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _28425_ (_03123_, _03122_, _01190_);
  and _28426_ (_03124_, _03123_, _03119_);
  and _28427_ (_03125_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _28428_ (_03126_, _03125_, rst);
  or _28429_ (_03127_, _03126_, _03124_);
  or _28430_ (_25288_, _03127_, _03118_);
  and _28431_ (_03128_, _02920_, _01597_);
  nand _28432_ (_03129_, _03128_, _01289_);
  or _28433_ (_03130_, _03128_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _28434_ (_03132_, _03130_, _01298_);
  and _28435_ (_03133_, _03132_, _03129_);
  nand _28436_ (_03134_, _02928_, _02204_);
  or _28437_ (_03135_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _28438_ (_03136_, _03135_, _01190_);
  and _28439_ (_03137_, _03136_, _03134_);
  and _28440_ (_03138_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _28441_ (_03139_, _03138_, rst);
  or _28442_ (_03140_, _03139_, _03137_);
  or _28443_ (_25289_, _03140_, _03133_);
  and _28444_ (_03141_, _02920_, _01680_);
  nand _28445_ (_03142_, _03141_, _01289_);
  or _28446_ (_03143_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _28447_ (_03144_, _03143_, _01298_);
  and _28448_ (_03145_, _03144_, _03142_);
  nand _28449_ (_03146_, _02928_, _02190_);
  or _28450_ (_03147_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _28451_ (_03148_, _03147_, _01190_);
  and _28452_ (_03149_, _03148_, _03146_);
  and _28453_ (_03150_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _28454_ (_03151_, _03150_, rst);
  or _28455_ (_03152_, _03151_, _03149_);
  or _28456_ (_25290_, _03152_, _03145_);
  and _28457_ (_03153_, _02920_, _01745_);
  nand _28458_ (_03154_, _03153_, _01289_);
  or _28459_ (_03155_, _03153_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _28460_ (_03156_, _03155_, _01298_);
  and _28461_ (_03157_, _03156_, _03154_);
  nand _28462_ (_03158_, _02928_, _02177_);
  or _28463_ (_03159_, _02928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _28464_ (_03160_, _03159_, _01190_);
  and _28465_ (_03161_, _03160_, _03158_);
  not _28466_ (_03162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _28467_ (_03163_, _01189_, _03162_);
  or _28468_ (_03164_, _03163_, rst);
  or _28469_ (_03165_, _03164_, _03161_);
  or _28470_ (_25291_, _03165_, _03157_);
  and _28471_ (_03166_, _02937_, _00860_);
  nand _28472_ (_03167_, _03166_, _01289_);
  or _28473_ (_03168_, _03166_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _28474_ (_03169_, _03168_, _01298_);
  and _28475_ (_03170_, _03169_, _03167_);
  and _28476_ (_03171_, _02944_, _02260_);
  not _28477_ (_03172_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _28478_ (_03173_, _02944_, _03172_);
  or _28479_ (_03174_, _03173_, _03171_);
  and _28480_ (_03175_, _03174_, _01190_);
  nor _28481_ (_03176_, _01189_, _03172_);
  or _28482_ (_03177_, _03176_, rst);
  or _28483_ (_03178_, _03177_, _03175_);
  or _28484_ (_25292_, _03178_, _03170_);
  and _28485_ (_03179_, _02937_, _02689_);
  nand _28486_ (_03180_, _03179_, _01289_);
  or _28487_ (_03181_, _03179_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _28488_ (_03182_, _03181_, _01298_);
  and _28489_ (_03183_, _03182_, _03180_);
  and _28490_ (_03184_, _02944_, _02251_);
  not _28491_ (_03185_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor _28492_ (_03186_, _02944_, _03185_);
  or _28493_ (_03187_, _03186_, _03184_);
  and _28494_ (_03188_, _03187_, _01190_);
  nor _28495_ (_03189_, _01189_, _03185_);
  or _28496_ (_03190_, _03189_, rst);
  or _28497_ (_03191_, _03190_, _03188_);
  or _28498_ (_25293_, _03191_, _03183_);
  and _28499_ (_03192_, _02937_, _01468_);
  nand _28500_ (_03193_, _03192_, _01289_);
  or _28501_ (_03194_, _03192_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _28502_ (_03195_, _03194_, _01298_);
  and _28503_ (_03196_, _03195_, _03193_);
  and _28504_ (_03197_, _02944_, _02236_);
  and _28505_ (_03198_, _02945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _28506_ (_03199_, _03198_, _03197_);
  and _28507_ (_03200_, _03199_, _01190_);
  and _28508_ (_03201_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _28509_ (_03202_, _03201_, rst);
  or _28510_ (_03203_, _03202_, _03200_);
  or _28511_ (_25294_, _03203_, _03196_);
  and _28512_ (_03204_, _02937_, _01530_);
  nand _28513_ (_03205_, _03204_, _01289_);
  or _28514_ (_03206_, _03204_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _28515_ (_03207_, _03206_, _01298_);
  and _28516_ (_03208_, _03207_, _03205_);
  and _28517_ (_03209_, _02944_, _02220_);
  and _28518_ (_03210_, _02945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _28519_ (_03211_, _03210_, _03209_);
  and _28520_ (_03212_, _03211_, _01190_);
  and _28521_ (_03213_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _28522_ (_03214_, _03213_, rst);
  or _28523_ (_03215_, _03214_, _03212_);
  or _28524_ (_25295_, _03215_, _03208_);
  and _28525_ (_03216_, _02937_, _01597_);
  nand _28526_ (_03217_, _03216_, _01289_);
  or _28527_ (_03218_, _03216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _28528_ (_03219_, _03218_, _01298_);
  and _28529_ (_03220_, _03219_, _03217_);
  nor _28530_ (_03221_, _02945_, _02204_);
  and _28531_ (_03222_, _02945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _28532_ (_03223_, _03222_, _03221_);
  and _28533_ (_03224_, _03223_, _01190_);
  and _28534_ (_03225_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _28535_ (_03226_, _03225_, rst);
  or _28536_ (_03227_, _03226_, _03224_);
  or _28537_ (_25296_, _03227_, _03220_);
  and _28538_ (_03228_, _02937_, _01680_);
  nand _28539_ (_03229_, _03228_, _01289_);
  or _28540_ (_03230_, _03228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _28541_ (_03231_, _03230_, _01298_);
  and _28542_ (_03232_, _03231_, _03229_);
  nor _28543_ (_03233_, _02945_, _02190_);
  and _28544_ (_03234_, _02945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _28545_ (_03235_, _03234_, _03233_);
  and _28546_ (_03236_, _03235_, _01190_);
  and _28547_ (_03237_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _28548_ (_03238_, _03237_, rst);
  or _28549_ (_03239_, _03238_, _03236_);
  or _28550_ (_25297_, _03239_, _03232_);
  and _28551_ (_03240_, _02937_, _01745_);
  nand _28552_ (_03241_, _03240_, _01289_);
  or _28553_ (_03242_, _03240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _28554_ (_03243_, _03242_, _01298_);
  and _28555_ (_03244_, _03243_, _03241_);
  nor _28556_ (_03245_, _02945_, _02177_);
  not _28557_ (_03246_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor _28558_ (_03247_, _02944_, _03246_);
  or _28559_ (_03248_, _03247_, _03245_);
  and _28560_ (_03249_, _03248_, _01190_);
  nor _28561_ (_03250_, _01189_, _03246_);
  or _28562_ (_03251_, _03250_, rst);
  or _28563_ (_03252_, _03251_, _03249_);
  or _28564_ (_25298_, _03252_, _03244_);
  and _28565_ (_03253_, _02953_, _00860_);
  nand _28566_ (_03254_, _03253_, _01289_);
  or _28567_ (_03255_, _03253_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _28568_ (_03256_, _03255_, _01298_);
  and _28569_ (_03257_, _03256_, _03254_);
  and _28570_ (_03258_, _02961_, _02260_);
  not _28571_ (_03259_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _28572_ (_03260_, _02961_, _03259_);
  or _28573_ (_03261_, _03260_, _03258_);
  and _28574_ (_03262_, _03261_, _01190_);
  nor _28575_ (_03263_, _01189_, _03259_);
  or _28576_ (_03264_, _03263_, rst);
  or _28577_ (_03265_, _03264_, _03262_);
  or _28578_ (_25299_, _03265_, _03257_);
  and _28579_ (_03266_, _02953_, _02689_);
  nand _28580_ (_03267_, _03266_, _01289_);
  or _28581_ (_03268_, _03266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _28582_ (_03269_, _03268_, _01298_);
  and _28583_ (_03270_, _03269_, _03267_);
  and _28584_ (_03271_, _02961_, _02251_);
  not _28585_ (_03272_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor _28586_ (_03273_, _02961_, _03272_);
  or _28587_ (_03274_, _03273_, _03271_);
  and _28588_ (_03275_, _03274_, _01190_);
  nor _28589_ (_03276_, _01189_, _03272_);
  or _28590_ (_03277_, _03276_, rst);
  or _28591_ (_03278_, _03277_, _03275_);
  or _28592_ (_25300_, _03278_, _03270_);
  and _28593_ (_03279_, _02953_, _01468_);
  nand _28594_ (_03280_, _03279_, _01289_);
  or _28595_ (_03281_, _03279_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _28596_ (_03282_, _03281_, _01298_);
  and _28597_ (_03283_, _03282_, _03280_);
  and _28598_ (_03284_, _02961_, _02236_);
  and _28599_ (_03285_, _02962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _28600_ (_03286_, _03285_, _03284_);
  and _28601_ (_03287_, _03286_, _01190_);
  and _28602_ (_03288_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _28603_ (_03289_, _03288_, rst);
  or _28604_ (_03290_, _03289_, _03287_);
  or _28605_ (_25301_, _03290_, _03283_);
  and _28606_ (_03291_, _02953_, _01530_);
  nand _28607_ (_03292_, _03291_, _01289_);
  or _28608_ (_03293_, _03291_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _28609_ (_03294_, _03293_, _01298_);
  and _28610_ (_03295_, _03294_, _03292_);
  and _28611_ (_03296_, _02961_, _02220_);
  and _28612_ (_03297_, _02962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _28613_ (_03298_, _03297_, _03296_);
  and _28614_ (_03299_, _03298_, _01190_);
  and _28615_ (_03300_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _28616_ (_03301_, _03300_, rst);
  or _28617_ (_03302_, _03301_, _03299_);
  or _28618_ (_25302_, _03302_, _03295_);
  and _28619_ (_03303_, _02953_, _01597_);
  nand _28620_ (_03304_, _03303_, _01289_);
  or _28621_ (_03305_, _03303_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _28622_ (_03306_, _03305_, _01298_);
  and _28623_ (_03307_, _03306_, _03304_);
  nor _28624_ (_03309_, _02962_, _02204_);
  and _28625_ (_03310_, _02962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _28626_ (_03311_, _03310_, _03309_);
  and _28627_ (_03312_, _03311_, _01190_);
  and _28628_ (_03313_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _28629_ (_03314_, _03313_, rst);
  or _28630_ (_03315_, _03314_, _03312_);
  or _28631_ (_25303_, _03315_, _03307_);
  and _28632_ (_03316_, _02953_, _01680_);
  nand _28633_ (_03317_, _03316_, _01289_);
  or _28634_ (_03318_, _03316_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _28635_ (_03319_, _03318_, _01298_);
  and _28636_ (_03320_, _03319_, _03317_);
  nor _28637_ (_03321_, _02962_, _02190_);
  and _28638_ (_03322_, _02962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _28639_ (_03323_, _03322_, _03321_);
  and _28640_ (_03324_, _03323_, _01190_);
  and _28641_ (_03325_, _02916_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _28642_ (_03326_, _03325_, rst);
  or _28643_ (_03327_, _03326_, _03324_);
  or _28644_ (_25304_, _03327_, _03320_);
  and _28645_ (_03328_, _02953_, _01745_);
  nand _28646_ (_03329_, _03328_, _01289_);
  or _28647_ (_03330_, _03328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _28648_ (_03331_, _03330_, _01298_);
  and _28649_ (_03332_, _03331_, _03329_);
  nor _28650_ (_03333_, _02962_, _02177_);
  not _28651_ (_03334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _28652_ (_03335_, _02961_, _03334_);
  or _28653_ (_03336_, _03335_, _03333_);
  and _28654_ (_03337_, _03336_, _01190_);
  nor _28655_ (_03338_, _01189_, _03334_);
  or _28656_ (_03339_, _03338_, rst);
  or _28657_ (_03340_, _03339_, _03337_);
  or _28658_ (_25305_, _03340_, _03332_);
  and _28659_ (_25306_, t0_i, _25365_);
  and _28660_ (_25307_, t1_i, _25365_);
  not _28661_ (_03341_, _01190_);
  nor _28662_ (_03342_, _03341_, _00921_);
  and _28663_ (_03343_, _03342_, _01530_);
  and _28664_ (_03344_, _03343_, _02162_);
  nand _28665_ (_03345_, _03344_, _02280_);
  not _28666_ (_03346_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _28667_ (_03347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _03346_);
  not _28668_ (_03348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _28669_ (_03349_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor _28670_ (_03350_, _03349_, _03347_);
  nor _28671_ (_03351_, _00835_, _00921_);
  and _28672_ (_03352_, _03351_, _02163_);
  and _28673_ (_03353_, _03352_, _01190_);
  or _28674_ (_03354_, _03353_, _03350_);
  and _28675_ (_03355_, _03354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _28676_ (_03356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _28677_ (_03357_, t1_i);
  and _28678_ (_03358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _03357_);
  nor _28679_ (_03359_, _03358_, _03356_);
  not _28680_ (_03360_, _03359_);
  not _28681_ (_03361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _28682_ (_03362_, _03361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nor _28683_ (_03363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _28684_ (_03364_, _03363_);
  and _28685_ (_03365_, _03364_, _03362_);
  and _28686_ (_03366_, _03365_, _03360_);
  and _28687_ (_03367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _28688_ (_03368_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _28689_ (_03369_, _03368_, _03367_);
  and _28690_ (_03370_, _03369_, _03366_);
  and _28691_ (_03371_, _03370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _28692_ (_03372_, _03371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _28693_ (_03373_, _03372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _28694_ (_03374_, _03373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _28695_ (_03375_, _03369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _28696_ (_03376_, _03375_, _03366_);
  and _28697_ (_03377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _28698_ (_03378_, _03377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _28699_ (_03379_, _03378_, _03376_);
  nor _28700_ (_03380_, _03379_, _03350_);
  and _28701_ (_03381_, _03380_, _03374_);
  and _28702_ (_03382_, _03379_, _03347_);
  and _28703_ (_03383_, _03382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _28704_ (_03384_, _03383_, _03381_);
  nor _28705_ (_03385_, _03384_, _03353_);
  or _28706_ (_03386_, _03385_, _03355_);
  or _28707_ (_03387_, _03386_, _03344_);
  and _28708_ (_03388_, _03387_, _25365_);
  and _28709_ (_25308_, _03388_, _03345_);
  and _28710_ (_03389_, _03344_, _25365_);
  and _28711_ (_03390_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _28712_ (_03391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _28713_ (_03392_, _03391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _28714_ (_03393_, _03392_, _03376_);
  and _28715_ (_03394_, _03393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _28716_ (_03395_, _03394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _28717_ (_03396_, _03395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _28718_ (_03397_, _03396_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _28719_ (_03398_, _03397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _28720_ (_03399_, _03397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _28721_ (_03400_, _03399_, _03378_);
  not _28722_ (_03401_, _03349_);
  nor _28723_ (_03402_, _03378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _28724_ (_03403_, _03402_, _03401_);
  nor _28725_ (_03404_, _03403_, _03400_);
  and _28726_ (_03405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _28727_ (_03406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not _28728_ (_03407_, _03406_);
  nor _28729_ (_03408_, _03399_, _03407_);
  or _28730_ (_03409_, _03408_, _03405_);
  or _28731_ (_03410_, _03409_, _03404_);
  nand _28732_ (_03411_, _03410_, _03398_);
  nor _28733_ (_03412_, _03411_, _03353_);
  not _28734_ (_03413_, _03353_);
  nor _28735_ (_03414_, _03413_, _02280_);
  or _28736_ (_03415_, _03414_, _03412_);
  nor _28737_ (_03416_, _03344_, rst);
  and _28738_ (_03417_, _03416_, _03415_);
  or _28739_ (_25309_, _03417_, _03390_);
  not _28740_ (_03418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _28741_ (_03419_, _03366_, _03418_);
  or _28742_ (_03420_, _03419_, _03400_);
  and _28743_ (_03421_, _03420_, _03349_);
  or _28744_ (_03422_, _03419_, _03399_);
  and _28745_ (_03423_, _03422_, _03406_);
  nand _28746_ (_03424_, _03366_, _03346_);
  and _28747_ (_03425_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _28748_ (_03426_, _03425_, _03424_);
  or _28749_ (_03427_, _03426_, _03382_);
  or _28750_ (_03428_, _03427_, _03423_);
  nor _28751_ (_03429_, _03428_, _03421_);
  nor _28752_ (_03430_, _03429_, _03353_);
  and _28753_ (_25310_, _03430_, _03416_);
  and _28754_ (_03431_, _03342_, _01597_);
  and _28755_ (_03432_, _03431_, _02162_);
  nor _28756_ (_03433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not _28757_ (_03434_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _28758_ (_03435_, t0_i);
  and _28759_ (_03436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _03435_);
  nor _28760_ (_03437_, _03436_, _03434_);
  not _28761_ (_03438_, _03437_);
  not _28762_ (_03439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _28763_ (_03440_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _28764_ (_03441_, _03440_, _03439_);
  and _28765_ (_03442_, _03441_, _03438_);
  and _28766_ (_03443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _28767_ (_03444_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _28768_ (_03445_, _03444_, _03443_);
  and _28769_ (_03446_, _03445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _28770_ (_03447_, _03446_, _03442_);
  and _28771_ (_03448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _28772_ (_03449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _28773_ (_03450_, _03449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _28774_ (_03451_, _03450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _28775_ (_03452_, _03451_, _03448_);
  and _28776_ (_03453_, _03452_, _03447_);
  and _28777_ (_03454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _28778_ (_03455_, _03454_, _03453_);
  and _28779_ (_03456_, _03455_, _03433_);
  not _28780_ (_03457_, _03442_);
  and _28781_ (_03458_, _03457_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _28782_ (_03459_, _03454_, _03452_);
  or _28783_ (_03460_, _03459_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _28784_ (_03461_, _03433_);
  and _28785_ (_03462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _28786_ (_03463_, _03462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _28787_ (_03464_, _03463_, _03447_);
  and _28788_ (_03465_, _03464_, _03461_);
  and _28789_ (_03466_, _03465_, _03460_);
  or _28790_ (_03467_, _03466_, _03458_);
  or _28791_ (_03468_, _03467_, _03456_);
  nand _28792_ (_03469_, _03468_, _25365_);
  nor _28793_ (_03470_, _03469_, _03432_);
  and _28794_ (_03471_, _03342_, _01468_);
  and _28795_ (_03472_, _03471_, _02162_);
  not _28796_ (_03473_, _03472_);
  and _28797_ (_25311_, _03473_, _03470_);
  nand _28798_ (_03474_, _03472_, _02280_);
  not _28799_ (_03475_, _03432_);
  or _28800_ (_03476_, _03475_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _28801_ (_03477_, _03433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _28802_ (_03478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _28803_ (_03479_, _03478_, _03447_);
  or _28804_ (_03480_, _03479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _28805_ (_03481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _28806_ (_03482_, _03481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _28807_ (_03483_, _03482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _28808_ (_03484_, _03483_, _03464_);
  and _28809_ (_03485_, _03484_, _03461_);
  or _28810_ (_03486_, _03485_, _03432_);
  and _28811_ (_03487_, _03486_, _03480_);
  or _28812_ (_03488_, _03487_, _03477_);
  and _28813_ (_03489_, _03488_, _03476_);
  or _28814_ (_03490_, _03489_, _03472_);
  and _28815_ (_03491_, _03490_, _25365_);
  and _28816_ (_25312_, _03491_, _03474_);
  nand _28817_ (_03492_, _03432_, _02280_);
  and _28818_ (_03493_, _03481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _28819_ (_03494_, _03482_, _03493_);
  not _28820_ (_03495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _28821_ (_03496_, _03463_, _03446_);
  and _28822_ (_03497_, _03442_, _03481_);
  and _28823_ (_03498_, _03497_, _03496_);
  and _28824_ (_03500_, _03498_, _03452_);
  and _28825_ (_03501_, _03500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _28826_ (_03502_, _03501_, _03495_);
  and _28827_ (_03503_, _03501_, _03495_);
  or _28828_ (_03504_, _03503_, _03502_);
  and _28829_ (_03505_, _03504_, _03494_);
  and _28830_ (_03506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _28831_ (_03507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _28832_ (_03508_, _03507_, _03451_);
  and _28833_ (_03509_, _03508_, _03448_);
  and _28834_ (_03510_, _03509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _28835_ (_03511_, _03510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _28836_ (_03512_, _03510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _28837_ (_03513_, _03512_, _03511_);
  and _28838_ (_03514_, _03513_, _03506_);
  and _28839_ (_03515_, _03453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _28840_ (_03516_, _03515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _28841_ (_03517_, _03455_, _03461_);
  and _28842_ (_03518_, _03517_, _03516_);
  or _28843_ (_03519_, _03518_, _03514_);
  or _28844_ (_03520_, _03519_, _03505_);
  or _28845_ (_03521_, _03520_, _03432_);
  and _28846_ (_03522_, _03521_, _03473_);
  and _28847_ (_03523_, _03522_, _03492_);
  and _28848_ (_03524_, _03472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _28849_ (_03525_, _03524_, _03523_);
  and _28850_ (_25313_, _03525_, _25365_);
  not _28851_ (_03526_, _03507_);
  or _28852_ (_03527_, _03526_, _03459_);
  or _28853_ (_03528_, _03507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _28854_ (_03529_, _03506_, _25365_);
  and _28855_ (_03530_, _03529_, _03528_);
  nand _28856_ (_03531_, _03530_, _03527_);
  nor _28857_ (_03532_, _03531_, _03432_);
  and _28858_ (_25314_, _03532_, _03473_);
  nor _28859_ (_03533_, _01291_, _00921_);
  and _28860_ (_03534_, _03533_, _02163_);
  and _28861_ (_03535_, _03534_, _01190_);
  or _28862_ (_03536_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _28863_ (_03537_, _03536_, _25365_);
  nand _28864_ (_03538_, _03535_, _02280_);
  and _28865_ (_25315_, _03538_, _03537_);
  and _28866_ (_03539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor _28867_ (_03540_, _03539_, _03353_);
  nor _28868_ (_03541_, _03366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _28869_ (_03542_, _03366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _28870_ (_03543_, _03542_, _03541_);
  and _28871_ (_03544_, _03543_, _03540_);
  not _28872_ (_03545_, _03540_);
  and _28873_ (_03546_, _03545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _28874_ (_03547_, _03546_, _03544_);
  and _28875_ (_03548_, _03378_, _03375_);
  and _28876_ (_03549_, _03548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _28877_ (_03550_, _03549_, _03347_);
  nor _28878_ (_03551_, _03550_, _03353_);
  or _28879_ (_03552_, _03551_, _03344_);
  or _28880_ (_03553_, _03552_, _03547_);
  nand _28881_ (_03554_, _03344_, _02259_);
  and _28882_ (_03555_, _03554_, _25365_);
  and _28883_ (_25316_, _03555_, _03553_);
  and _28884_ (_03556_, _03542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _28885_ (_03557_, _03542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _28886_ (_03558_, _03557_, _03556_);
  and _28887_ (_03559_, _03558_, _03540_);
  and _28888_ (_03560_, _03545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _28889_ (_03561_, _03560_, _03559_);
  and _28890_ (_03562_, _03373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _28891_ (_03563_, _03562_, _03347_);
  nand _28892_ (_03564_, _03563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _28893_ (_03565_, _03564_, _03353_);
  or _28894_ (_03566_, _03565_, _03344_);
  or _28895_ (_03567_, _03566_, _03561_);
  not _28896_ (_03568_, _03344_);
  or _28897_ (_03569_, _03568_, _02251_);
  and _28898_ (_03570_, _03569_, _25365_);
  and _28899_ (_25317_, _03570_, _03567_);
  nor _28900_ (_03571_, _03556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _28901_ (_03572_, _03542_, _03367_);
  nor _28902_ (_03573_, _03572_, _03571_);
  and _28903_ (_03574_, _03573_, _03540_);
  and _28904_ (_03575_, _03545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _28905_ (_03576_, _03575_, _03574_);
  nand _28906_ (_03577_, _03563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _28907_ (_03578_, _03577_, _03353_);
  or _28908_ (_03579_, _03578_, _03344_);
  or _28909_ (_03580_, _03579_, _03576_);
  or _28910_ (_03581_, _03568_, _02236_);
  and _28911_ (_03582_, _03581_, _25365_);
  and _28912_ (_25318_, _03582_, _03580_);
  and _28913_ (_03583_, _03545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _28914_ (_03584_, _03572_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _28915_ (_03585_, _03539_, _03370_);
  and _28916_ (_03586_, _03585_, _03584_);
  and _28917_ (_03587_, _03382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _28918_ (_03588_, _03587_, _03586_);
  nor _28919_ (_03589_, _03588_, _03353_);
  or _28920_ (_03590_, _03589_, _03583_);
  and _28921_ (_03591_, _03590_, _03416_);
  and _28922_ (_03592_, _03389_, _02220_);
  or _28923_ (_25319_, _03592_, _03591_);
  and _28924_ (_03593_, _03545_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _28925_ (_03594_, _03382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _28926_ (_03595_, _03594_, _03353_);
  or _28927_ (_03596_, _03595_, _03593_);
  nor _28928_ (_03597_, _03370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _28929_ (_03598_, _03597_, _03376_);
  and _28930_ (_03599_, _03598_, _03540_);
  or _28931_ (_03600_, _03599_, _03344_);
  or _28932_ (_03601_, _03600_, _03596_);
  nand _28933_ (_03602_, _03344_, _02204_);
  and _28934_ (_03603_, _03602_, _25365_);
  and _28935_ (_25320_, _03603_, _03601_);
  not _28936_ (_03604_, _02190_);
  and _28937_ (_03605_, _03389_, _03604_);
  and _28938_ (_03606_, _03354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _28939_ (_03607_, _03563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _28940_ (_03608_, _03350_);
  and _28941_ (_03609_, _03376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _28942_ (_03610_, _03376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _28943_ (_03611_, _03610_, _03609_);
  and _28944_ (_03612_, _03611_, _03608_);
  nor _28945_ (_03613_, _03612_, _03607_);
  nor _28946_ (_03614_, _03613_, _03353_);
  or _28947_ (_03615_, _03614_, _03606_);
  and _28948_ (_03616_, _03615_, _03416_);
  or _28949_ (_25321_, _03616_, _03605_);
  and _28950_ (_03617_, _03354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _28951_ (_03618_, _03347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _28952_ (_03619_, _03618_, _03366_);
  and _28953_ (_03620_, _03619_, _03548_);
  or _28954_ (_03621_, _03609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _28955_ (_03622_, _03621_, _03608_);
  nor _28956_ (_03623_, _03622_, _03373_);
  nor _28957_ (_03624_, _03623_, _03620_);
  nor _28958_ (_03625_, _03624_, _03353_);
  or _28959_ (_03626_, _03625_, _03617_);
  and _28960_ (_03627_, _03626_, _03416_);
  not _28961_ (_03628_, _02177_);
  and _28962_ (_03629_, _03389_, _03628_);
  or _28963_ (_25322_, _03629_, _03627_);
  and _28964_ (_03630_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  not _28965_ (_03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _28966_ (_03632_, _03378_, _03346_);
  not _28967_ (_03633_, _03632_);
  and _28968_ (_03634_, _03376_, _03348_);
  and _28969_ (_03635_, _03634_, _03633_);
  nor _28970_ (_03636_, _03635_, _03631_);
  and _28971_ (_03637_, _03635_, _03631_);
  or _28972_ (_03638_, _03637_, _03636_);
  or _28973_ (_03639_, _03638_, _03353_);
  nand _28974_ (_03640_, _03353_, _02259_);
  and _28975_ (_03641_, _03640_, _03416_);
  and _28976_ (_03642_, _03641_, _03639_);
  or _28977_ (_25323_, _03642_, _03630_);
  and _28978_ (_03643_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _28979_ (_03644_, _03413_, _02251_);
  not _28980_ (_03645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _28981_ (_03646_, _03634_, _03401_);
  and _28982_ (_03647_, _03379_, _03349_);
  nor _28983_ (_03648_, _03647_, _03646_);
  nor _28984_ (_03649_, _03648_, _03631_);
  nor _28985_ (_03650_, _03649_, _03645_);
  and _28986_ (_03651_, _03649_, _03645_);
  or _28987_ (_03652_, _03651_, _03650_);
  or _28988_ (_03653_, _03652_, _03353_);
  and _28989_ (_03654_, _03653_, _03416_);
  and _28990_ (_03655_, _03654_, _03644_);
  or _28991_ (_25324_, _03655_, _03643_);
  and _28992_ (_03656_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _28993_ (_03657_, _03413_, _02236_);
  nand _28994_ (_03658_, _03393_, _03348_);
  or _28995_ (_03659_, _03658_, _03632_);
  and _28996_ (_03660_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _28997_ (_03661_, _03632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _28998_ (_03662_, _03661_);
  not _28999_ (_03663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _29000_ (_03664_, _03391_, _03663_);
  and _29001_ (_03665_, _03664_, _03376_);
  and _29002_ (_03666_, _03665_, _03662_);
  or _29003_ (_03667_, _03666_, _03660_);
  or _29004_ (_03668_, _03667_, _03353_);
  and _29005_ (_03669_, _03668_, _03416_);
  and _29006_ (_03670_, _03669_, _03657_);
  or _29007_ (_25325_, _03670_, _03656_);
  and _29008_ (_03671_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _29009_ (_03672_, _03413_, _02220_);
  and _29010_ (_03673_, _03391_, _03548_);
  and _29011_ (_03674_, _03673_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _29012_ (_03675_, _03674_, _03366_);
  nor _29013_ (_03676_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _29014_ (_03677_, _03675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _29015_ (_03678_, _03677_, _03676_);
  nor _29016_ (_03679_, _03678_, _03401_);
  and _29017_ (_03680_, _03658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _29018_ (_03681_, _03658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _29019_ (_03682_, _03681_, _03680_);
  and _29020_ (_03683_, _03682_, _03401_);
  or _29021_ (_03684_, _03683_, _03679_);
  or _29022_ (_03685_, _03684_, _03353_);
  and _29023_ (_03686_, _03685_, _03416_);
  and _29024_ (_03688_, _03686_, _03672_);
  or _29025_ (_25326_, _03688_, _03671_);
  and _29026_ (_03689_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _29027_ (_03690_, _03353_, _02204_);
  or _29028_ (_03691_, _03677_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _29029_ (_03692_, _03691_, _03349_);
  and _29030_ (_03693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _29031_ (_03694_, _03675_, _03693_);
  nor _29032_ (_03695_, _03694_, _03692_);
  nor _29033_ (_03696_, _03394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _29034_ (_03697_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _29035_ (_03698_, _03395_, _03407_);
  nor _29036_ (_03699_, _03698_, _03697_);
  nor _29037_ (_03700_, _03699_, _03696_);
  or _29038_ (_03701_, _03700_, _03695_);
  or _29039_ (_03702_, _03701_, _03353_);
  and _29040_ (_03703_, _03702_, _03416_);
  and _29041_ (_03704_, _03703_, _03690_);
  or _29042_ (_25327_, _03704_, _03689_);
  and _29043_ (_03705_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand _29044_ (_03706_, _03353_, _02190_);
  and _29045_ (_03707_, _03694_, _03348_);
  nor _29046_ (_03708_, _03707_, _03406_);
  nor _29047_ (_03709_, _03708_, _03698_);
  or _29048_ (_03710_, _03709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand _29049_ (_03711_, _03709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _29050_ (_03712_, _03711_, _03710_);
  or _29051_ (_03713_, _03712_, _03353_);
  and _29052_ (_03714_, _03713_, _03416_);
  and _29053_ (_03715_, _03714_, _03706_);
  or _29054_ (_25328_, _03715_, _03705_);
  and _29055_ (_03716_, _03389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _29056_ (_03717_, _03353_, _02177_);
  and _29057_ (_03718_, _03662_, _03396_);
  or _29058_ (_03719_, _03718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _29059_ (_03720_, _03718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _29060_ (_03721_, _03720_, _03719_);
  or _29061_ (_03722_, _03721_, _03353_);
  and _29062_ (_03723_, _03722_, _03416_);
  and _29063_ (_03724_, _03723_, _03717_);
  or _29064_ (_25329_, _03724_, _03716_);
  nor _29065_ (_03725_, _03457_, _03432_);
  or _29066_ (_03726_, _03725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _29067_ (_03727_, _03442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _29068_ (_03728_, _03482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _29069_ (_03729_, _03728_, _03496_);
  nand _29070_ (_03730_, _03729_, _03727_);
  or _29071_ (_03731_, _03730_, _03432_);
  and _29072_ (_03732_, _03731_, _03726_);
  or _29073_ (_03733_, _03732_, _03472_);
  nand _29074_ (_03734_, _03472_, _02259_);
  and _29075_ (_03735_, _03734_, _25365_);
  and _29076_ (_25330_, _03735_, _03733_);
  nor _29077_ (_03736_, _03727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _29078_ (_03737_, _03727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _29079_ (_03738_, _03737_, _03736_);
  and _29080_ (_03739_, _03482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _29081_ (_03740_, _03739_, _03464_);
  nor _29082_ (_03741_, _03740_, _03738_);
  nor _29083_ (_03742_, _03741_, _03432_);
  and _29084_ (_03743_, _03432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _29085_ (_03744_, _03743_, _03742_);
  and _29086_ (_03745_, _03744_, _03473_);
  and _29087_ (_03746_, _03472_, _02251_);
  or _29088_ (_03747_, _03746_, _03745_);
  and _29089_ (_25331_, _03747_, _25365_);
  and _29090_ (_03748_, _03342_, _02424_);
  not _29091_ (_03749_, _03748_);
  or _29092_ (_03750_, _03749_, _02236_);
  nor _29093_ (_03751_, _03737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _29094_ (_03752_, _03727_, _03443_);
  nor _29095_ (_03753_, _03752_, _03751_);
  and _29096_ (_03754_, _03482_, _03464_);
  and _29097_ (_03755_, _03754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _29098_ (_03756_, _03755_, _03753_);
  nor _29099_ (_03757_, _03756_, _03432_);
  and _29100_ (_03758_, _03432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _29101_ (_03759_, _03758_, _03757_);
  or _29102_ (_03760_, _03759_, _03748_);
  and _29103_ (_03761_, _03760_, _25365_);
  and _29104_ (_25332_, _03761_, _03750_);
  or _29105_ (_03762_, _03749_, _02220_);
  and _29106_ (_03763_, _03445_, _03442_);
  nor _29107_ (_03764_, _03752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _29108_ (_03765_, _03764_, _03763_);
  and _29109_ (_03766_, _03754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _29110_ (_03767_, _03766_, _03765_);
  nor _29111_ (_03768_, _03767_, _03432_);
  and _29112_ (_03769_, _03432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _29113_ (_03770_, _03769_, _03768_);
  or _29114_ (_03771_, _03770_, _03748_);
  and _29115_ (_03772_, _03771_, _25365_);
  and _29116_ (_25333_, _03772_, _03762_);
  nand _29117_ (_03773_, _03748_, _02204_);
  nor _29118_ (_03774_, _03763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _29119_ (_03775_, _03774_, _03447_);
  and _29120_ (_03776_, _03754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _29121_ (_03777_, _03776_, _03775_);
  nor _29122_ (_03778_, _03777_, _03432_);
  and _29123_ (_03779_, _03432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _29124_ (_03780_, _03779_, _03778_);
  or _29125_ (_03781_, _03780_, _03748_);
  and _29126_ (_03782_, _03781_, _25365_);
  and _29127_ (_25334_, _03782_, _03773_);
  and _29128_ (_03783_, _03754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _29129_ (_03784_, _03447_, _03461_);
  or _29130_ (_03785_, _03784_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _29131_ (_03786_, _03784_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand _29132_ (_03787_, _03786_, _03475_);
  and _29133_ (_03788_, _03787_, _03785_);
  or _29134_ (_03789_, _03788_, _03783_);
  or _29135_ (_03790_, _03475_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _29136_ (_03791_, _03790_, _03473_);
  and _29137_ (_03792_, _03791_, _03789_);
  nor _29138_ (_03793_, _03473_, _02190_);
  or _29139_ (_03794_, _03793_, _03792_);
  and _29140_ (_25335_, _03794_, _25365_);
  not _29141_ (_03795_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _29142_ (_03796_, _03786_, _03795_);
  and _29143_ (_03797_, _03482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _29144_ (_03798_, _03797_, _03442_);
  and _29145_ (_03799_, _03798_, _03496_);
  nor _29146_ (_03800_, _03799_, _03796_);
  nor _29147_ (_03801_, _03800_, _03432_);
  and _29148_ (_03802_, _03787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _29149_ (_03803_, _03802_, _03801_);
  and _29150_ (_03804_, _03803_, _03473_);
  nor _29151_ (_03805_, _03473_, _02177_);
  or _29152_ (_03806_, _03805_, _03804_);
  and _29153_ (_25336_, _03806_, _25365_);
  or _29154_ (_03807_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _29155_ (_03808_, _03807_, _03494_);
  and _29156_ (_03809_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _29157_ (_03810_, _03809_, _03808_);
  and _29158_ (_03811_, _03507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _29159_ (_03812_, _03507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _29160_ (_03813_, _03812_, _03506_);
  nor _29161_ (_03814_, _03813_, _03811_);
  and _29162_ (_03815_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _29163_ (_03816_, _03447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _29164_ (_03817_, _03816_, _03433_);
  nor _29165_ (_03818_, _03817_, _03815_);
  or _29166_ (_03819_, _03818_, _03814_);
  or _29167_ (_03820_, _03819_, _03810_);
  or _29168_ (_03821_, _03820_, _03432_);
  nand _29169_ (_03822_, _03432_, _02259_);
  and _29170_ (_03823_, _03822_, _03821_);
  or _29171_ (_03824_, _03823_, _03472_);
  or _29172_ (_03825_, _03473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _29173_ (_03826_, _03825_, _25365_);
  and _29174_ (_25337_, _03826_, _03824_);
  or _29175_ (_03827_, _03475_, _02251_);
  or _29176_ (_03828_, _03809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _29177_ (_03829_, _03496_, _03442_);
  and _29178_ (_03830_, _03829_, _03449_);
  not _29179_ (_03831_, _03830_);
  or _29180_ (_03832_, _03831_, _03482_);
  and _29181_ (_03833_, _03832_, _03494_);
  and _29182_ (_03834_, _03833_, _03828_);
  and _29183_ (_03835_, _03507_, _03449_);
  or _29184_ (_03836_, _03811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _29185_ (_03837_, _03836_, _03506_);
  nor _29186_ (_03838_, _03837_, _03835_);
  and _29187_ (_03839_, _03815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _29188_ (_03840_, _03815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _29189_ (_03841_, _03840_, _03433_);
  nor _29190_ (_03842_, _03841_, _03839_);
  or _29191_ (_03843_, _03842_, _03838_);
  or _29192_ (_03844_, _03843_, _03834_);
  nor _29193_ (_03845_, _03844_, _03432_);
  nor _29194_ (_03846_, _03845_, _03748_);
  and _29195_ (_03847_, _03846_, _03827_);
  and _29196_ (_03848_, _03748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _29197_ (_03849_, _03848_, _03847_);
  and _29198_ (_25338_, _03849_, _25365_);
  or _29199_ (_03850_, _03475_, _02236_);
  or _29200_ (_03851_, _03830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _29201_ (_03852_, _03829_, _03450_);
  not _29202_ (_03853_, _03852_);
  and _29203_ (_03854_, _03853_, _03493_);
  and _29204_ (_03855_, _03854_, _03851_);
  and _29205_ (_03856_, _03449_, _03442_);
  and _29206_ (_03857_, _03856_, _03446_);
  or _29207_ (_03858_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _29208_ (_03859_, _03450_, _03447_);
  nor _29209_ (_03860_, _03859_, _03461_);
  and _29210_ (_03861_, _03860_, _03858_);
  and _29211_ (_03862_, _03835_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _29212_ (_03863_, _03862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _29213_ (_03864_, _03507_, _03450_);
  nand _29214_ (_03865_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _29215_ (_03866_, _03865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _29216_ (_03867_, _03866_, _03863_);
  or _29217_ (_03868_, _03867_, _03861_);
  or _29218_ (_03869_, _03868_, _03855_);
  nor _29219_ (_03870_, _03869_, _03432_);
  nor _29220_ (_03871_, _03870_, _03748_);
  and _29221_ (_03872_, _03871_, _03850_);
  and _29222_ (_03873_, _03472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _29223_ (_03874_, _03873_, _03872_);
  and _29224_ (_25339_, _03874_, _25365_);
  or _29225_ (_03876_, _03475_, _02220_);
  not _29226_ (_03877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _29227_ (_03878_, _03852_, _03481_);
  nor _29228_ (_03879_, _03878_, _03877_);
  and _29229_ (_03880_, _03878_, _03877_);
  or _29230_ (_03881_, _03880_, _03879_);
  and _29231_ (_03882_, _03881_, _03494_);
  or _29232_ (_03883_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _29233_ (_03884_, _03508_);
  and _29234_ (_03885_, _03884_, _03506_);
  and _29235_ (_03886_, _03885_, _03883_);
  or _29236_ (_03887_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _29237_ (_03888_, _03451_, _03447_);
  nor _29238_ (_03889_, _03888_, _03461_);
  and _29239_ (_03890_, _03889_, _03887_);
  or _29240_ (_03891_, _03890_, _03886_);
  or _29241_ (_03892_, _03891_, _03882_);
  nor _29242_ (_03893_, _03892_, _03432_);
  nor _29243_ (_03894_, _03893_, _03748_);
  and _29244_ (_03895_, _03894_, _03876_);
  and _29245_ (_03896_, _03472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _29246_ (_03897_, _03896_, _03895_);
  and _29247_ (_25340_, _03897_, _25365_);
  nand _29248_ (_03898_, _03432_, _02204_);
  or _29249_ (_03899_, _03888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _29250_ (_03900_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _29251_ (_03901_, _03900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _29252_ (_03902_, _03901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _29253_ (_03903_, _03902_, _03461_);
  and _29254_ (_03904_, _03903_, _03899_);
  and _29255_ (_03905_, _03829_, _03451_);
  or _29256_ (_03906_, _03905_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _29257_ (_03907_, _03906_, _03493_);
  nand _29258_ (_03908_, _03905_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _29259_ (_03909_, _03908_, _03907_);
  and _29260_ (_03910_, _03508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _29261_ (_03911_, _03910_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _29262_ (_03912_, _03508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _29263_ (_03913_, _03912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _29264_ (_03914_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _29265_ (_03915_, _03914_, _03911_);
  or _29266_ (_03916_, _03915_, _03909_);
  or _29267_ (_03917_, _03916_, _03904_);
  nor _29268_ (_03918_, _03917_, _03432_);
  nor _29269_ (_03919_, _03918_, _03748_);
  and _29270_ (_03920_, _03919_, _03898_);
  and _29271_ (_03921_, _03748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _29272_ (_03922_, _03921_, _03920_);
  and _29273_ (_25341_, _03922_, _25365_);
  nand _29274_ (_03923_, _03432_, _02190_);
  not _29275_ (_03924_, _03902_);
  nor _29276_ (_03925_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _29277_ (_03926_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _29278_ (_03927_, _03926_, _03925_);
  and _29279_ (_03928_, _03927_, _03433_);
  nor _29280_ (_03929_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _29281_ (_03930_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _29282_ (_03931_, _03929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _29283_ (_03932_, _03931_, _03494_);
  and _29284_ (_03933_, _03932_, _03930_);
  not _29285_ (_03934_, _03509_);
  and _29286_ (_03935_, _03934_, _03506_);
  or _29287_ (_03936_, _03910_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _29288_ (_03937_, _03936_, _03935_);
  or _29289_ (_03938_, _03937_, _03933_);
  or _29290_ (_03939_, _03938_, _03928_);
  or _29291_ (_03940_, _03939_, _03432_);
  and _29292_ (_03941_, _03940_, _03749_);
  and _29293_ (_03942_, _03941_, _03923_);
  and _29294_ (_03943_, _03472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _29295_ (_03944_, _03943_, _03942_);
  and _29296_ (_25342_, _03944_, _25365_);
  nand _29297_ (_03945_, _03432_, _02177_);
  or _29298_ (_03946_, _03500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _29299_ (_03947_, _03946_, _03494_);
  nor _29300_ (_03948_, _03947_, _03501_);
  or _29301_ (_03949_, _03509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _29302_ (_03950_, _03510_);
  and _29303_ (_03951_, _03950_, _03506_);
  and _29304_ (_03952_, _03951_, _03949_);
  or _29305_ (_03953_, _03453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _29306_ (_03954_, _03515_, _03461_);
  and _29307_ (_03955_, _03954_, _03953_);
  or _29308_ (_03956_, _03955_, _03952_);
  or _29309_ (_03957_, _03956_, _03948_);
  nor _29310_ (_03958_, _03957_, _03432_);
  nor _29311_ (_03959_, _03958_, _03748_);
  and _29312_ (_03960_, _03959_, _03945_);
  and _29313_ (_03961_, _03472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _29314_ (_03962_, _03961_, _03960_);
  and _29315_ (_25343_, _03962_, _25365_);
  nand _29316_ (_03963_, _03535_, _02259_);
  or _29317_ (_03964_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _29318_ (_03965_, _03964_, _25365_);
  and _29319_ (_25344_, _03965_, _03963_);
  or _29320_ (_03966_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _29321_ (_03967_, _03966_, _25365_);
  not _29322_ (_03968_, _03535_);
  or _29323_ (_03969_, _03968_, _02251_);
  and _29324_ (_25345_, _03969_, _03967_);
  or _29325_ (_03970_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _29326_ (_03971_, _03970_, _25365_);
  or _29327_ (_03972_, _03968_, _02236_);
  and _29328_ (_25346_, _03972_, _03971_);
  or _29329_ (_03973_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _29330_ (_03974_, _03973_, _25365_);
  or _29331_ (_03975_, _03968_, _02220_);
  and _29332_ (_25347_, _03975_, _03974_);
  or _29333_ (_03976_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _29334_ (_03977_, _03976_, _25365_);
  nand _29335_ (_03978_, _03535_, _02204_);
  and _29336_ (_25348_, _03978_, _03977_);
  or _29337_ (_03979_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _29338_ (_03980_, _03979_, _25365_);
  nand _29339_ (_03981_, _03535_, _02190_);
  and _29340_ (_25349_, _03981_, _03980_);
  or _29341_ (_03982_, _03535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _29342_ (_03983_, _03982_, _25365_);
  nand _29343_ (_03984_, _03535_, _02177_);
  and _29344_ (_25350_, _03984_, _03983_);
  not _29345_ (_03985_, _00938_);
  nor _29346_ (_03986_, _02795_, _00921_);
  nand _29347_ (_03987_, _03986_, _03985_);
  nor _29348_ (_03988_, _03987_, _00906_);
  and _29349_ (_03989_, _03988_, _02936_);
  and _29350_ (_03990_, _03989_, _01294_);
  nand _29351_ (_03991_, _03990_, _01289_);
  and _29352_ (_03992_, _02157_, _01294_);
  and _29353_ (_03993_, _03992_, _02960_);
  not _29354_ (_03994_, _03993_);
  or _29355_ (_03995_, _03990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _29356_ (_03996_, _03995_, _03994_);
  and _29357_ (_03997_, _03996_, _03991_);
  nor _29358_ (_03998_, _03994_, _02280_);
  or _29359_ (_03999_, _03998_, _03997_);
  and _29360_ (_25351_, _03999_, _25365_);
  and _29361_ (_04000_, _03342_, _00860_);
  and _29362_ (_04001_, _04000_, _02943_);
  not _29363_ (_04002_, _04001_);
  and _29364_ (_04003_, _00938_, _00922_);
  and _29365_ (_04004_, _04003_, _02796_);
  and _29366_ (_04005_, _04004_, _02936_);
  and _29367_ (_04006_, _04005_, _01294_);
  or _29368_ (_04007_, _04006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _29369_ (_04008_, _04007_, _04002_);
  nand _29370_ (_04009_, _04006_, _01289_);
  and _29371_ (_04010_, _04009_, _04008_);
  nor _29372_ (_04011_, _04002_, _02280_);
  or _29373_ (_04012_, _04011_, _04010_);
  and _29374_ (_25352_, _04012_, _25365_);
  and _29375_ (_04013_, _04000_, _02162_);
  and _29376_ (_04014_, _03986_, _00938_);
  and _29377_ (_04015_, _04014_, _00907_);
  and _29378_ (_04016_, _04015_, _02903_);
  nand _29379_ (_04017_, _04016_, _00858_);
  and _29380_ (_04018_, _04017_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _29381_ (_04019_, _04018_, _04013_);
  or _29382_ (_04020_, _00859_, _01467_);
  and _29383_ (_04021_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _29384_ (_04022_, _04021_, _02773_);
  and _29385_ (_04023_, _04022_, _04016_);
  or _29386_ (_04024_, _04023_, _04019_);
  nand _29387_ (_04025_, _04013_, _02177_);
  and _29388_ (_04026_, _04025_, _25365_);
  and _29389_ (_25353_, _04026_, _04024_);
  not _29390_ (_04027_, _04013_);
  nor _29391_ (_04028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _29392_ (_04029_, _04028_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _29393_ (_04030_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _29394_ (_04031_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _29395_ (_04032_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _29396_ (_04033_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _04032_);
  and _29397_ (_04034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29398_ (_04035_, _04034_, _04033_);
  nor _29399_ (_04036_, _04035_, _04031_);
  or _29400_ (_04037_, _04036_, _04030_);
  and _29401_ (_04038_, _04032_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _29402_ (_04039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _29403_ (_04040_, _04039_, _04038_);
  nor _29404_ (_04041_, _04040_, _04031_);
  and _29405_ (_04042_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _04032_);
  and _29406_ (_04043_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29407_ (_04044_, _04043_, _04042_);
  nand _29408_ (_04045_, _04044_, _04041_);
  or _29409_ (_04046_, _04045_, _04037_);
  and _29410_ (_04047_, _04046_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _29411_ (_04048_, _04047_, _04029_);
  and _29412_ (_04049_, _02162_, _01294_);
  and _29413_ (_04050_, _04049_, _03986_);
  or _29414_ (_04051_, _04050_, _04048_);
  and _29415_ (_04052_, _04051_, _04027_);
  nand _29416_ (_04053_, _04050_, _01289_);
  and _29417_ (_04054_, _04053_, _04052_);
  nor _29418_ (_04055_, _04027_, _02280_);
  or _29419_ (_04056_, _04055_, _04054_);
  and _29420_ (_25354_, _04056_, _25365_);
  and _29421_ (_04057_, _03352_, _01298_);
  nand _29422_ (_04058_, _04057_, _01289_);
  not _29423_ (_04059_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _29424_ (_04061_, _04059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _29425_ (_04062_, _04044_, _04031_);
  not _29426_ (_04063_, _04062_);
  or _29427_ (_04064_, _04063_, _04041_);
  or _29428_ (_04065_, _04064_, _04037_);
  and _29429_ (_04066_, _04065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _29430_ (_04067_, _04066_, _04061_);
  or _29431_ (_04068_, _04067_, _04057_);
  and _29432_ (_04069_, _04068_, _04027_);
  and _29433_ (_04070_, _04069_, _04058_);
  nor _29434_ (_04071_, _04027_, _02190_);
  or _29435_ (_04072_, _04071_, _04070_);
  and _29436_ (_25355_, _04072_, _25365_);
  not _29437_ (_04073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _29438_ (_04074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _04073_);
  nand _29439_ (_04075_, _04036_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _29440_ (_04076_, _04062_, _04041_);
  or _29441_ (_04077_, _04076_, _04075_);
  and _29442_ (_04078_, _04077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _29443_ (_04079_, _04078_, _04074_);
  and _29444_ (_04080_, _03534_, _01298_);
  or _29445_ (_04081_, _04080_, _04079_);
  and _29446_ (_04082_, _04081_, _04027_);
  nand _29447_ (_04083_, _04080_, _01289_);
  and _29448_ (_04084_, _04083_, _04082_);
  and _29449_ (_04085_, _04013_, _02251_);
  or _29450_ (_04086_, _04085_, _04084_);
  and _29451_ (_25356_, _04086_, _25365_);
  and _29452_ (_04087_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _29453_ (_04088_, _04075_, _04064_);
  and _29454_ (_04089_, _04088_, _04087_);
  and _29455_ (_04090_, _03986_, _02416_);
  or _29456_ (_04091_, _04090_, _04089_);
  and _29457_ (_04092_, _04091_, _04027_);
  nand _29458_ (_04093_, _04090_, _01289_);
  and _29459_ (_04094_, _04093_, _04092_);
  and _29460_ (_04095_, _04013_, _02220_);
  or _29461_ (_04096_, _04095_, _04094_);
  and _29462_ (_25357_, _04096_, _25365_);
  nand _29463_ (_04097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _29464_ (_04098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _04032_);
  and _29465_ (_04099_, _04098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _29466_ (_04100_, _04099_, _04097_);
  or _29467_ (_04101_, _04100_, _04031_);
  and _29468_ (_04102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _29469_ (_04103_, _04102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _29470_ (_04104_, _04103_);
  and _29471_ (_04105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _29472_ (_04106_, _04105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _29473_ (_04107_, _04106_);
  and _29474_ (_04108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _29475_ (_04109_, _04108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29476_ (_04110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _29477_ (_04111_, _04110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _29478_ (_04112_, _04111_, _04109_);
  and _29479_ (_04113_, _04112_, _04107_);
  and _29480_ (_04114_, _04113_, _04104_);
  not _29481_ (_04115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _29482_ (_04116_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _29483_ (_04117_, _04116_, _04115_);
  nand _29484_ (_04118_, _04117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _29485_ (_04119_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _29486_ (_04120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _29487_ (_04121_, _04120_, _04119_);
  and _29488_ (_04122_, _04121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _29489_ (_04123_, _04122_);
  and _29490_ (_04124_, _04123_, _04118_);
  nand _29491_ (_04125_, _04124_, _04114_);
  and _29492_ (_04126_, _04125_, _04101_);
  and _29493_ (_04127_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _29494_ (_04128_, _04127_, _04032_);
  and _29495_ (_04129_, _04128_, _04126_);
  not _29496_ (_04130_, _04129_);
  not _29497_ (_04131_, _04128_);
  and _29498_ (_04132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _04031_);
  not _29499_ (_04133_, _04132_);
  not _29500_ (_04134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _29501_ (_04135_, _04105_, _04134_);
  not _29502_ (_04136_, _04135_);
  not _29503_ (_04137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29504_ (_04138_, _04108_, _04137_);
  not _29505_ (_04139_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _29506_ (_04140_, _04110_, _04139_);
  nor _29507_ (_04141_, _04140_, _04138_);
  and _29508_ (_04142_, _04141_, _04136_);
  nor _29509_ (_04143_, _04142_, _04133_);
  not _29510_ (_04144_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _29511_ (_04145_, _04117_, _04144_);
  not _29512_ (_04146_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _29513_ (_04147_, _04121_, _04146_);
  nor _29514_ (_04148_, _04147_, _04145_);
  not _29515_ (_04149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _29516_ (_04150_, _04102_, _04149_);
  not _29517_ (_04151_, _04150_);
  and _29518_ (_04152_, _04151_, _04148_);
  nor _29519_ (_04153_, _04152_, _04133_);
  nor _29520_ (_04154_, _04153_, _04143_);
  or _29521_ (_04155_, _04154_, _04131_);
  and _29522_ (_04156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _25365_);
  and _29523_ (_04157_, _04156_, _04155_);
  and _29524_ (_25358_, _04157_, _04130_);
  nor _29525_ (_04158_, _04127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _29526_ (_04159_, _04158_);
  not _29527_ (_04160_, _04126_);
  and _29528_ (_04161_, _04154_, _04160_);
  nor _29529_ (_04162_, _04161_, _04159_);
  nand _29530_ (_04163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _25365_);
  nor _29531_ (_25359_, _04163_, _04162_);
  and _29532_ (_04164_, _04124_, _04104_);
  nand _29533_ (_04165_, _04164_, _04126_);
  or _29534_ (_04166_, _04153_, _04126_);
  and _29535_ (_04167_, _04166_, _04128_);
  and _29536_ (_04168_, _04167_, _04165_);
  or _29537_ (_04169_, _04168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _29538_ (_04170_, _04130_, _04113_);
  nor _29539_ (_04171_, _04131_, _04126_);
  nand _29540_ (_04172_, _04171_, _04143_);
  and _29541_ (_04173_, _04172_, _25365_);
  and _29542_ (_04174_, _04173_, _04170_);
  and _29543_ (_25360_, _04174_, _04169_);
  and _29544_ (_04175_, _04165_, _04158_);
  or _29545_ (_04176_, _04175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _29546_ (_04177_, _04158_, _04126_);
  not _29547_ (_04178_, _04177_);
  or _29548_ (_04179_, _04178_, _04113_);
  or _29549_ (_04180_, _04153_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand _29550_ (_04181_, _04158_, _04143_);
  and _29551_ (_04182_, _04181_, _04180_);
  or _29552_ (_04183_, _04182_, _04126_);
  and _29553_ (_04184_, _04183_, _25365_);
  and _29554_ (_04185_, _04184_, _04179_);
  and _29555_ (_25361_, _04185_, _04176_);
  nand _29556_ (_04186_, _04161_, _04031_);
  nor _29557_ (_04187_, _04032_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _29558_ (_04188_, _04187_, _04127_);
  and _29559_ (_04189_, _04188_, _25365_);
  and _29560_ (_25362_, _04189_, _04186_);
  and _29561_ (_04190_, _04161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _29562_ (_04191_, _04032_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _29563_ (_04192_, _04191_, _04187_);
  nor _29564_ (_04193_, _04192_, _04160_);
  or _29565_ (_04194_, _04193_, _04127_);
  or _29566_ (_04195_, _04194_, _04190_);
  not _29567_ (_04196_, _04127_);
  or _29568_ (_04197_, _04192_, _04196_);
  and _29569_ (_04198_, _04197_, _25365_);
  and _29570_ (_25363_, _04198_, _04195_);
  and _29571_ (_04199_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _25365_);
  and _29572_ (_25364_, _04199_, _04127_);
  nor _29573_ (_25366_, _04028_, rst);
  and _29574_ (_25367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _25365_);
  nor _29575_ (_04200_, _04161_, _04127_);
  and _29576_ (_04201_, _04127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _29577_ (_04202_, _04201_, _04200_);
  and _29578_ (_00010_, _04202_, _25365_);
  and _29579_ (_04203_, _04127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _29580_ (_04204_, _04203_, _04200_);
  and _29581_ (_00012_, _04204_, _25365_);
  and _29582_ (_04205_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _25365_);
  and _29583_ (_00014_, _04205_, _04127_);
  not _29584_ (_04206_, _04140_);
  nor _29585_ (_04207_, _04147_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _29586_ (_04208_, _04207_, _04145_);
  or _29587_ (_04209_, _04208_, _04150_);
  and _29588_ (_04210_, _04209_, _04206_);
  or _29589_ (_04211_, _04210_, _04138_);
  nor _29590_ (_04212_, _04154_, _04126_);
  and _29591_ (_04213_, _04212_, _04136_);
  and _29592_ (_04214_, _04213_, _04211_);
  not _29593_ (_04215_, _04111_);
  or _29594_ (_04216_, _04122_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _29595_ (_04217_, _04216_, _04118_);
  or _29596_ (_04218_, _04217_, _04103_);
  and _29597_ (_04219_, _04218_, _04215_);
  or _29598_ (_04220_, _04219_, _04109_);
  and _29599_ (_04221_, _04126_, _04107_);
  and _29600_ (_04222_, _04221_, _04220_);
  or _29601_ (_04223_, _04222_, _04127_);
  or _29602_ (_04224_, _04223_, _04214_);
  or _29603_ (_04225_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _29604_ (_04226_, _04225_, _25365_);
  and _29605_ (_00016_, _04226_, _04224_);
  not _29606_ (_04227_, _04109_);
  or _29607_ (_04228_, _04111_, _04103_);
  and _29608_ (_04229_, _04124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _29609_ (_04230_, _04229_, _04228_);
  and _29610_ (_04231_, _04230_, _04227_);
  and _29611_ (_04232_, _04231_, _04221_);
  nor _29612_ (_04233_, _04138_, _04135_);
  or _29613_ (_04234_, _04150_, _04140_);
  and _29614_ (_04235_, _04148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _29615_ (_04236_, _04235_, _04234_);
  and _29616_ (_04237_, _04236_, _04233_);
  and _29617_ (_04238_, _04237_, _04212_);
  or _29618_ (_04239_, _04238_, _04127_);
  or _29619_ (_04240_, _04239_, _04232_);
  or _29620_ (_04241_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _29621_ (_04242_, _04241_, _25365_);
  and _29622_ (_00017_, _04242_, _04240_);
  and _29623_ (_04244_, _04151_, _04132_);
  nand _29624_ (_04245_, _04244_, _04142_);
  or _29625_ (_04246_, _04245_, _04148_);
  nor _29626_ (_04247_, _04246_, _04126_);
  nand _29627_ (_04248_, _04114_, _04101_);
  nor _29628_ (_04249_, _04248_, _04124_);
  or _29629_ (_04250_, _04249_, _04127_);
  or _29630_ (_04251_, _04250_, _04247_);
  or _29631_ (_04252_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _29632_ (_04253_, _04252_, _25365_);
  and _29633_ (_00019_, _04253_, _04251_);
  and _29634_ (_04254_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _25365_);
  and _29635_ (_00021_, _04254_, _04127_);
  and _29636_ (_04255_, _04127_, _04032_);
  or _29637_ (_04256_, _04255_, _04162_);
  or _29638_ (_04257_, _04256_, _04171_);
  and _29639_ (_00022_, _04257_, _25365_);
  not _29640_ (_04258_, _04200_);
  and _29641_ (_04259_, _04258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _29642_ (_04260_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _29643_ (_04261_, _04122_, _04032_);
  or _29644_ (_04262_, _04261_, _04260_);
  nor _29645_ (_04263_, _04118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29646_ (_04264_, _04263_, _04103_);
  nand _29647_ (_04265_, _04264_, _04262_);
  or _29648_ (_04266_, _04104_, _04034_);
  and _29649_ (_04267_, _04266_, _04265_);
  or _29650_ (_04268_, _04267_, _04111_);
  or _29651_ (_04269_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _04032_);
  or _29652_ (_04270_, _04269_, _04215_);
  and _29653_ (_04271_, _04270_, _04227_);
  and _29654_ (_04272_, _04271_, _04268_);
  and _29655_ (_04273_, _04109_, _04034_);
  or _29656_ (_04274_, _04273_, _04106_);
  or _29657_ (_04275_, _04274_, _04272_);
  or _29658_ (_04276_, _04269_, _04107_);
  and _29659_ (_04277_, _04276_, _04126_);
  and _29660_ (_04278_, _04277_, _04275_);
  and _29661_ (_04279_, _04147_, _04032_);
  or _29662_ (_04280_, _04279_, _04260_);
  and _29663_ (_04281_, _04145_, _04032_);
  nor _29664_ (_04282_, _04281_, _04150_);
  nand _29665_ (_04283_, _04282_, _04280_);
  or _29666_ (_04284_, _04151_, _04034_);
  and _29667_ (_04285_, _04284_, _04283_);
  or _29668_ (_04286_, _04285_, _04140_);
  not _29669_ (_04287_, _04138_);
  or _29670_ (_04288_, _04269_, _04206_);
  and _29671_ (_04289_, _04288_, _04287_);
  and _29672_ (_04290_, _04289_, _04286_);
  and _29673_ (_04291_, _04138_, _04034_);
  or _29674_ (_04292_, _04291_, _04135_);
  or _29675_ (_04293_, _04292_, _04290_);
  and _29676_ (_04294_, _04269_, _04212_);
  or _29677_ (_04295_, _04294_, _04213_);
  and _29678_ (_04296_, _04295_, _04293_);
  or _29679_ (_04297_, _04296_, _04278_);
  and _29680_ (_04298_, _04297_, _04196_);
  or _29681_ (_04299_, _04298_, _04259_);
  and _29682_ (_00024_, _04299_, _25365_);
  and _29683_ (_04300_, _04135_, _04043_);
  or _29684_ (_04301_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _04032_);
  and _29685_ (_04302_, _04301_, _04136_);
  or _29686_ (_04303_, _04302_, _04142_);
  and _29687_ (_04304_, _04150_, _04043_);
  not _29688_ (_04305_, _04141_);
  or _29689_ (_04306_, _04279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _29690_ (_04307_, _04306_, _04282_);
  or _29691_ (_04308_, _04307_, _04305_);
  or _29692_ (_04309_, _04308_, _04304_);
  and _29693_ (_04310_, _04309_, _04303_);
  or _29694_ (_04311_, _04310_, _04300_);
  and _29695_ (_04312_, _04311_, _04212_);
  or _29696_ (_04313_, _04261_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _29697_ (_04314_, _04313_, _04264_);
  and _29698_ (_04315_, _04103_, _04043_);
  or _29699_ (_04316_, _04315_, _04314_);
  and _29700_ (_04317_, _04316_, _04112_);
  not _29701_ (_04318_, _04112_);
  and _29702_ (_04319_, _04301_, _04318_);
  or _29703_ (_04320_, _04319_, _04106_);
  or _29704_ (_04321_, _04320_, _04317_);
  or _29705_ (_04322_, _04107_, _04043_);
  and _29706_ (_04323_, _04322_, _04126_);
  and _29707_ (_04324_, _04323_, _04321_);
  and _29708_ (_04325_, _04161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _29709_ (_04326_, _04325_, _04127_);
  or _29710_ (_04327_, _04326_, _04324_);
  or _29711_ (_04328_, _04327_, _04312_);
  or _29712_ (_04329_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _29713_ (_04330_, _04329_, _25365_);
  and _29714_ (_00026_, _04330_, _04328_);
  and _29715_ (_04331_, _04258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _29716_ (_04332_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29717_ (_04333_, _04332_, _04107_);
  and _29718_ (_04334_, _04333_, _04126_);
  not _29719_ (_04335_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _29720_ (_04336_, _04122_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29721_ (_04337_, _04336_, _04335_);
  nor _29722_ (_04338_, _04118_, _04032_);
  nor _29723_ (_04340_, _04338_, _04103_);
  nand _29724_ (_04341_, _04340_, _04337_);
  or _29725_ (_04342_, _04104_, _04033_);
  and _29726_ (_04343_, _04342_, _04341_);
  or _29727_ (_04344_, _04343_, _04111_);
  or _29728_ (_04345_, _04332_, _04215_);
  and _29729_ (_04346_, _04345_, _04227_);
  and _29730_ (_04347_, _04346_, _04344_);
  and _29731_ (_04348_, _04109_, _04033_);
  or _29732_ (_04349_, _04348_, _04106_);
  or _29733_ (_04350_, _04349_, _04347_);
  and _29734_ (_04351_, _04350_, _04334_);
  or _29735_ (_04352_, _04332_, _04136_);
  and _29736_ (_04353_, _04147_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29737_ (_04354_, _04353_, _04335_);
  and _29738_ (_04355_, _04145_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29739_ (_04356_, _04355_, _04150_);
  nand _29740_ (_04357_, _04356_, _04354_);
  or _29741_ (_04358_, _04151_, _04033_);
  and _29742_ (_04359_, _04358_, _04357_);
  or _29743_ (_04360_, _04359_, _04140_);
  or _29744_ (_04361_, _04332_, _04206_);
  and _29745_ (_04362_, _04361_, _04287_);
  and _29746_ (_04363_, _04362_, _04360_);
  and _29747_ (_04364_, _04138_, _04033_);
  or _29748_ (_04365_, _04364_, _04135_);
  or _29749_ (_04366_, _04365_, _04363_);
  and _29750_ (_04367_, _04366_, _04212_);
  and _29751_ (_04368_, _04367_, _04352_);
  or _29752_ (_04369_, _04368_, _04351_);
  and _29753_ (_04370_, _04369_, _04196_);
  or _29754_ (_04371_, _04370_, _04331_);
  and _29755_ (_00028_, _04371_, _25365_);
  and _29756_ (_04372_, _04258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _29757_ (_04373_, _04336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _29758_ (_04374_, _04373_, _04340_);
  and _29759_ (_04375_, _04103_, _04042_);
  or _29760_ (_04376_, _04375_, _04374_);
  and _29761_ (_04377_, _04376_, _04112_);
  or _29762_ (_04378_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _29763_ (_04379_, _04378_, _04318_);
  or _29764_ (_04380_, _04379_, _04106_);
  or _29765_ (_04381_, _04380_, _04377_);
  or _29766_ (_04382_, _04107_, _04042_);
  and _29767_ (_04383_, _04382_, _04126_);
  and _29768_ (_04384_, _04383_, _04381_);
  and _29769_ (_04385_, _04135_, _04042_);
  and _29770_ (_04386_, _04378_, _04136_);
  or _29771_ (_04387_, _04386_, _04142_);
  and _29772_ (_04388_, _04150_, _04042_);
  or _29773_ (_04389_, _04353_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _29774_ (_04390_, _04389_, _04356_);
  or _29775_ (_04391_, _04390_, _04305_);
  or _29776_ (_04392_, _04391_, _04388_);
  and _29777_ (_04393_, _04392_, _04387_);
  or _29778_ (_04394_, _04393_, _04385_);
  and _29779_ (_04395_, _04394_, _04212_);
  or _29780_ (_04396_, _04395_, _04384_);
  and _29781_ (_04397_, _04396_, _04196_);
  or _29782_ (_04398_, _04397_, _04372_);
  and _29783_ (_00030_, _04398_, _25365_);
  or _29784_ (_04399_, _04159_, _04154_);
  and _29785_ (_04400_, _04399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _29786_ (_04401_, _04400_, _04177_);
  and _29787_ (_00032_, _04401_, _25365_);
  and _29788_ (_04402_, _04155_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _29789_ (_04403_, _04402_, _04129_);
  and _29790_ (_00034_, _04403_, _25365_);
  and _29791_ (_04404_, _04016_, _00860_);
  or _29792_ (_04405_, _04404_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _29793_ (_04406_, _04405_, _04027_);
  nand _29794_ (_04407_, _04404_, _01289_);
  and _29795_ (_04408_, _04407_, _04406_);
  and _29796_ (_04409_, _04013_, _02260_);
  or _29797_ (_04410_, _04409_, _04408_);
  and _29798_ (_00036_, _04410_, _25365_);
  not _29799_ (_04411_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _29800_ (_04412_, _04016_, _01468_);
  nand _29801_ (_04413_, _04412_, _04411_);
  and _29802_ (_04414_, _04413_, _04027_);
  or _29803_ (_04415_, _04412_, _01344_);
  and _29804_ (_04416_, _04415_, _04414_);
  and _29805_ (_04417_, _04013_, _02236_);
  or _29806_ (_04418_, _04417_, _04416_);
  and _29807_ (_00038_, _04418_, _25365_);
  nand _29808_ (_04419_, _04016_, _01597_);
  nand _29809_ (_04420_, _04419_, _03439_);
  and _29810_ (_04421_, _04420_, _04027_);
  or _29811_ (_04422_, _04419_, _01344_);
  and _29812_ (_04423_, _04422_, _04421_);
  nor _29813_ (_04424_, _04027_, _02204_);
  or _29814_ (_04425_, _04424_, _04423_);
  and _29815_ (_00040_, _04425_, _25365_);
  and _29816_ (_04426_, _04005_, _00860_);
  or _29817_ (_04427_, _04426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _29818_ (_04428_, _04427_, _04002_);
  nand _29819_ (_04429_, _04426_, _01289_);
  and _29820_ (_04430_, _04429_, _04428_);
  and _29821_ (_04431_, _04001_, _02260_);
  or _29822_ (_04432_, _04431_, _04430_);
  and _29823_ (_00042_, _04432_, _25365_);
  and _29824_ (_04434_, _04005_, _02689_);
  or _29825_ (_04435_, _04434_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _29826_ (_04436_, _04435_, _04002_);
  nand _29827_ (_04437_, _04434_, _01289_);
  and _29828_ (_04438_, _04437_, _04436_);
  and _29829_ (_04439_, _04001_, _02251_);
  or _29830_ (_04440_, _04439_, _04438_);
  and _29831_ (_00044_, _04440_, _25365_);
  nand _29832_ (_04441_, _04005_, _02998_);
  and _29833_ (_04442_, _04441_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _29834_ (_04443_, _04442_, _04001_);
  and _29835_ (_04444_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _29836_ (_04445_, _04444_, _01470_);
  and _29837_ (_04446_, _04445_, _04005_);
  or _29838_ (_04447_, _04446_, _04443_);
  or _29839_ (_04448_, _04002_, _02236_);
  and _29840_ (_04449_, _04448_, _25365_);
  and _29841_ (_00046_, _04449_, _04447_);
  and _29842_ (_04450_, _04005_, _01530_);
  or _29843_ (_04451_, _04450_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _29844_ (_04452_, _04451_, _04002_);
  nand _29845_ (_04453_, _04450_, _01289_);
  and _29846_ (_04454_, _04453_, _04452_);
  and _29847_ (_04455_, _04001_, _02220_);
  or _29848_ (_04456_, _04455_, _04454_);
  and _29849_ (_00048_, _04456_, _25365_);
  and _29850_ (_04457_, _04005_, _01597_);
  or _29851_ (_04458_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _29852_ (_04459_, _04458_, _04002_);
  nand _29853_ (_04460_, _04457_, _01289_);
  and _29854_ (_04461_, _04460_, _04459_);
  nor _29855_ (_04462_, _04002_, _02204_);
  or _29856_ (_04463_, _04462_, _04461_);
  and _29857_ (_00050_, _04463_, _25365_);
  and _29858_ (_04464_, _04005_, _01680_);
  or _29859_ (_04465_, _04464_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _29860_ (_04466_, _04465_, _04002_);
  nand _29861_ (_04467_, _04464_, _01289_);
  and _29862_ (_04468_, _04467_, _04466_);
  nor _29863_ (_04469_, _04002_, _02190_);
  or _29864_ (_04470_, _04469_, _04468_);
  and _29865_ (_00052_, _04470_, _25365_);
  and _29866_ (_04471_, _04005_, _01745_);
  or _29867_ (_04472_, _04471_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _29868_ (_04473_, _04472_, _04002_);
  nand _29869_ (_04474_, _04471_, _01289_);
  and _29870_ (_04475_, _04474_, _04473_);
  nor _29871_ (_04476_, _04002_, _02177_);
  or _29872_ (_04477_, _04476_, _04475_);
  and _29873_ (_00054_, _04477_, _25365_);
  and _29874_ (_04478_, _03989_, _00860_);
  nand _29875_ (_04479_, _04478_, _01289_);
  or _29876_ (_04480_, _04478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _29877_ (_04481_, _04480_, _03994_);
  and _29878_ (_04482_, _04481_, _04479_);
  and _29879_ (_04483_, _03993_, _02260_);
  or _29880_ (_04484_, _04483_, _04482_);
  and _29881_ (_00056_, _04484_, _25365_);
  and _29882_ (_04485_, _03989_, _02689_);
  nand _29883_ (_04486_, _04485_, _01289_);
  or _29884_ (_04487_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29885_ (_04488_, _04487_, _03994_);
  and _29886_ (_04489_, _04488_, _04486_);
  and _29887_ (_04490_, _03993_, _02251_);
  or _29888_ (_04491_, _04490_, _04489_);
  and _29889_ (_00058_, _04491_, _25365_);
  and _29890_ (_04492_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _29891_ (_04493_, _04492_, _01470_);
  and _29892_ (_04494_, _04493_, _03989_);
  nand _29893_ (_04495_, _03989_, _02998_);
  and _29894_ (_04496_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _29895_ (_04497_, _04496_, _03993_);
  or _29896_ (_04498_, _04497_, _04494_);
  or _29897_ (_04499_, _03994_, _02236_);
  and _29898_ (_04500_, _04499_, _25365_);
  and _29899_ (_00060_, _04500_, _04498_);
  and _29900_ (_04501_, _03989_, _01530_);
  nand _29901_ (_04502_, _04501_, _01289_);
  or _29902_ (_04503_, _04501_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _29903_ (_04504_, _04503_, _03994_);
  and _29904_ (_04505_, _04504_, _04502_);
  and _29905_ (_04506_, _03993_, _02220_);
  or _29906_ (_04507_, _04506_, _04505_);
  and _29907_ (_00062_, _04507_, _25365_);
  and _29908_ (_04508_, _03989_, _01597_);
  nand _29909_ (_04509_, _04508_, _01289_);
  or _29910_ (_04510_, _04508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _29911_ (_04511_, _04510_, _03994_);
  and _29912_ (_04512_, _04511_, _04509_);
  nor _29913_ (_04513_, _03994_, _02204_);
  or _29914_ (_04514_, _04513_, _04512_);
  and _29915_ (_00064_, _04514_, _25365_);
  and _29916_ (_04515_, _03989_, _01680_);
  nand _29917_ (_04516_, _04515_, _01289_);
  or _29918_ (_04517_, _04515_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _29919_ (_04518_, _04517_, _03994_);
  and _29920_ (_04519_, _04518_, _04516_);
  nor _29921_ (_04520_, _03994_, _02190_);
  or _29922_ (_04521_, _04520_, _04519_);
  and _29923_ (_00066_, _04521_, _25365_);
  and _29924_ (_04523_, _03989_, _01745_);
  nand _29925_ (_04524_, _04523_, _01289_);
  or _29926_ (_04525_, _04523_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _29927_ (_04526_, _04525_, _03994_);
  and _29928_ (_04527_, _04526_, _04524_);
  nor _29929_ (_04528_, _03994_, _02177_);
  or _29930_ (_04529_, _04528_, _04527_);
  and _29931_ (_00068_, _04529_, _25365_);
  and _29932_ (_04530_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _29933_ (_04531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _29934_ (_04532_, _04028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _29935_ (_04533_, _04532_, _04531_);
  not _29936_ (_04534_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _29937_ (_04535_, _04534_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _29938_ (_04536_, _04535_, _04533_);
  nor _29939_ (_04537_, _04536_, _04530_);
  or _29940_ (_04538_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _29941_ (_04539_, _04538_, _25365_);
  nor _29942_ (_00491_, _04539_, _04537_);
  nor _29943_ (_04540_, _04537_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _29944_ (_04541_, _04540_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _29945_ (_04542_, _04540_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _29946_ (_04543_, _04542_, _25365_);
  and _29947_ (_00493_, _04543_, _04541_);
  not _29948_ (_04544_, rxd_i);
  and _29949_ (_04545_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _04544_);
  nor _29950_ (_04546_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _29951_ (_04547_, _04546_);
  and _29952_ (_04548_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _29953_ (_04549_, _04548_, _04547_);
  and _29954_ (_04550_, _04549_, _04545_);
  not _29955_ (_04551_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _29956_ (_04552_, _04551_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _29957_ (_04553_, _04552_, _04546_);
  or _29958_ (_04554_, _04553_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or _29959_ (_04555_, _04554_, _04550_);
  and _29960_ (_04556_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _25365_);
  and _29961_ (_00496_, _04556_, _04555_);
  and _29962_ (_04557_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _29963_ (_04558_, _04557_, _04547_);
  nor _29964_ (_04559_, _04546_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _29965_ (_04560_, _04559_, _04551_);
  nor _29966_ (_04561_, _04560_, _04558_);
  not _29967_ (_04562_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _29968_ (_04563_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _04562_);
  not _29969_ (_04564_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _29970_ (_04565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _04564_);
  and _29971_ (_04566_, _04565_, _04563_);
  not _29972_ (_04567_, _04566_);
  or _29973_ (_04568_, _04567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and _29974_ (_04569_, _04566_, _04558_);
  and _29975_ (_04570_, _04558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _29976_ (_04571_, _04570_, _04569_);
  and _29977_ (_04572_, _04571_, _04568_);
  or _29978_ (_04573_, _04572_, _04561_);
  and _29979_ (_04574_, _04546_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _29980_ (_04575_, _04574_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not _29981_ (_04576_, _04575_);
  or _29982_ (_04577_, _04576_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _29983_ (_04578_, _04577_, _04573_);
  nand _29984_ (_00498_, _04578_, _04556_);
  not _29985_ (_04579_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _29986_ (_04580_, _04558_);
  nor _29987_ (_04581_, _04551_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _29988_ (_04582_, _04581_);
  not _29989_ (_04583_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _29990_ (_04584_, _04546_, _04583_);
  and _29991_ (_04585_, _04584_, _04582_);
  and _29992_ (_04586_, _04585_, _04580_);
  nor _29993_ (_04587_, _04586_, _04579_);
  and _29994_ (_04588_, _04586_, rxd_i);
  or _29995_ (_04589_, _04588_, rst);
  or _29996_ (_00501_, _04589_, _04587_);
  nor _29997_ (_04590_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _29998_ (_04591_, _04590_, _04563_);
  and _29999_ (_04592_, _04591_, _04570_);
  nand _30000_ (_04593_, _04592_, _04544_);
  or _30001_ (_04594_, _04592_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _30002_ (_04595_, _04594_, _25365_);
  and _30003_ (_00503_, _04595_, _04593_);
  and _30004_ (_04596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _30005_ (_04597_, _04596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _30006_ (_04598_, _04597_, _04562_);
  and _30007_ (_04599_, _04598_, _04570_);
  and _30008_ (_04600_, _04549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _30009_ (_04601_, _04600_, _04570_);
  nor _30010_ (_04602_, _04597_, _04580_);
  or _30011_ (_04603_, _04602_, _04601_);
  and _30012_ (_04604_, _04603_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _30013_ (_04605_, _04604_, _04599_);
  and _30014_ (_00506_, _04605_, _25365_);
  and _30015_ (_04606_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _25365_);
  nand _30016_ (_04607_, _04606_, _04583_);
  nand _30017_ (_04608_, _04556_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _30018_ (_00509_, _04608_, _04607_);
  and _30019_ (_04609_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _04583_);
  not _30020_ (_04610_, _04549_);
  not _30021_ (_04611_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _30022_ (_04612_, _04553_, _04611_);
  and _30023_ (_04614_, _04612_, _04610_);
  nand _30024_ (_04615_, _04614_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _30025_ (_04616_, _04615_, _04580_);
  or _30026_ (_04617_, _04566_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _30027_ (_04618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _30028_ (_04619_, _04618_, _04569_);
  and _30029_ (_04620_, _04619_, _04617_);
  and _30030_ (_04621_, _04620_, _04616_);
  or _30031_ (_04622_, _04621_, _04575_);
  nand _30032_ (_04623_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _30033_ (_04624_, _04623_, _04558_);
  or _30034_ (_04625_, _04624_, _04567_);
  and _30035_ (_04626_, _04625_, _04576_);
  or _30036_ (_04627_, _04626_, rxd_i);
  and _30037_ (_04628_, _04627_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _30038_ (_04629_, _04628_, _04622_);
  or _30039_ (_04630_, _04629_, _04609_);
  and _30040_ (_00511_, _04630_, _25365_);
  and _30041_ (_04631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _30042_ (_04632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _30043_ (_04633_, _04532_, _04632_);
  or _30044_ (_04634_, _04633_, _04535_);
  nor _30045_ (_04635_, _04634_, _04631_);
  or _30046_ (_04636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _30047_ (_04637_, _04636_, _25365_);
  nor _30048_ (_00514_, _04637_, _04635_);
  nor _30049_ (_04638_, _04635_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _30050_ (_04639_, _04638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _30051_ (_04640_, _04638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _30052_ (_04641_, _04640_, _25365_);
  and _30053_ (_00517_, _04641_, _04639_);
  and _30054_ (_04642_, _04574_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _30055_ (_04643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _30056_ (_04644_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _30057_ (_04645_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _30058_ (_04646_, _04645_, _04644_);
  and _30059_ (_04647_, _04646_, _04643_);
  not _30060_ (_04648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _30061_ (_04649_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _30062_ (_04650_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _30063_ (_04651_, _04650_, _04649_);
  and _30064_ (_04652_, _04651_, _04648_);
  and _30065_ (_04653_, _04652_, _04647_);
  or _30066_ (_04654_, _04653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _30067_ (_04655_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _30068_ (_04656_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _30069_ (_04657_, _04656_, _04655_);
  and _30070_ (_04658_, _04547_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _30071_ (_04659_, _04658_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _30072_ (_04660_, _04659_, _04657_);
  not _30073_ (_04661_, _04660_);
  or _30074_ (_04662_, _04661_, _04654_);
  and _30075_ (_04663_, _04657_, _04658_);
  not _30076_ (_04664_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or _30077_ (_04665_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _04664_);
  or _30078_ (_04666_, _04665_, _04663_);
  and _30079_ (_04667_, _04666_, _04662_);
  or _30080_ (_04668_, _04667_, _04642_);
  not _30081_ (_04669_, _04642_);
  not _30082_ (_04670_, _04653_);
  or _30083_ (_04671_, _04670_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _30084_ (_04672_, _04671_, _04654_);
  or _30085_ (_04673_, _04672_, _04669_);
  nand _30086_ (_04674_, _04673_, _04668_);
  and _30087_ (_04675_, _03533_, _01406_);
  and _30088_ (_04676_, _04675_, _01190_);
  and _30089_ (_04677_, _04676_, _02927_);
  nor _30090_ (_04678_, _04677_, rst);
  nand _30091_ (_04679_, _04678_, _04674_);
  not _30092_ (_04680_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _30093_ (_04681_, _04677_, _25365_);
  nand _30094_ (_04682_, _04681_, _04680_);
  and _30095_ (_00519_, _04682_, _04679_);
  nor _30096_ (_04683_, _04670_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _30097_ (_04684_, _04663_, _04683_);
  and _30098_ (_04685_, _04653_, _04642_);
  or _30099_ (_04686_, _04664_, rst);
  nor _30100_ (_04687_, _04686_, _04685_);
  and _30101_ (_04688_, _04687_, _04684_);
  or _30102_ (_00522_, _04688_, _04681_);
  or _30103_ (_04689_, _04661_, _04683_);
  or _30104_ (_04690_, _04663_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _30105_ (_04691_, _04574_, _04664_);
  and _30106_ (_04692_, _04691_, _04690_);
  and _30107_ (_04693_, _04692_, _04689_);
  or _30108_ (_04694_, _04693_, _04685_);
  and _30109_ (_00525_, _04694_, _04678_);
  and _30110_ (_04695_, _04659_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _30111_ (_04696_, _04695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _30112_ (_04697_, _04696_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _30113_ (_04698_, _04697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _30114_ (_04699_, _04697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _30115_ (_04700_, _04699_, _04698_);
  and _30116_ (_00527_, _04700_, _04678_);
  nor _30117_ (_04701_, _04660_, _04642_);
  and _30118_ (_04702_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _30119_ (_04703_, _04702_, _04678_);
  and _30120_ (_04704_, _04681_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _30121_ (_00530_, _04704_, _04703_);
  and _30122_ (_04705_, _03992_, _02162_);
  or _30123_ (_04707_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _30124_ (_04708_, _04707_, _25365_);
  nand _30125_ (_04709_, _04705_, _02280_);
  and _30126_ (_00532_, _04709_, _04708_);
  and _30127_ (_04710_, _03988_, _02903_);
  and _30128_ (_04711_, _04710_, _01294_);
  nand _30129_ (_04712_, _04711_, _01289_);
  and _30130_ (_04713_, _04000_, _02927_);
  not _30131_ (_04714_, _04713_);
  or _30132_ (_04715_, _04711_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _30133_ (_04716_, _04715_, _04714_);
  and _30134_ (_04717_, _04716_, _04712_);
  nor _30135_ (_04718_, _04714_, _02280_);
  or _30136_ (_04719_, _04718_, _04717_);
  and _30137_ (_00535_, _04719_, _25365_);
  nor _30138_ (_04720_, _04575_, _04569_);
  not _30139_ (_04721_, _04720_);
  nor _30140_ (_04722_, _04614_, _04558_);
  nor _30141_ (_04723_, _04722_, _04721_);
  nor _30142_ (_04724_, _04723_, _04583_);
  or _30143_ (_04725_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _30144_ (_04726_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _04583_);
  or _30145_ (_04727_, _04726_, _04720_);
  and _30146_ (_04728_, _04727_, _25365_);
  and _30147_ (_01196_, _04728_, _04725_);
  or _30148_ (_04729_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _30149_ (_04730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _04583_);
  or _30150_ (_04731_, _04730_, _04720_);
  and _30151_ (_04732_, _04731_, _25365_);
  and _30152_ (_01198_, _04732_, _04729_);
  or _30153_ (_04733_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _30154_ (_04734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _04583_);
  or _30155_ (_04735_, _04734_, _04720_);
  and _30156_ (_04736_, _04735_, _25365_);
  and _30157_ (_01200_, _04736_, _04733_);
  or _30158_ (_04737_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _30159_ (_04738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _04583_);
  or _30160_ (_04739_, _04738_, _04720_);
  and _30161_ (_04740_, _04739_, _25365_);
  and _30162_ (_01202_, _04740_, _04737_);
  or _30163_ (_04741_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _30164_ (_04742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _04583_);
  or _30165_ (_04743_, _04742_, _04720_);
  and _30166_ (_04744_, _04743_, _25365_);
  and _30167_ (_01204_, _04744_, _04741_);
  or _30168_ (_04745_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _30169_ (_04746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _04583_);
  or _30170_ (_04747_, _04746_, _04720_);
  and _30171_ (_04748_, _04747_, _25365_);
  and _30172_ (_01206_, _04748_, _04745_);
  or _30173_ (_04749_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _30174_ (_04750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _04583_);
  or _30175_ (_04751_, _04750_, _04720_);
  and _30176_ (_04752_, _04751_, _25365_);
  and _30177_ (_01208_, _04752_, _04749_);
  or _30178_ (_04753_, _04724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _30179_ (_04754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _04583_);
  or _30180_ (_04755_, _04754_, _04720_);
  and _30181_ (_04756_, _04755_, _25365_);
  and _30182_ (_01210_, _04756_, _04753_);
  nor _30183_ (_04757_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _30184_ (_04758_, _04757_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _30185_ (_04759_, _04567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _30186_ (_04760_, _04566_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _30187_ (_04761_, _04760_, _04558_);
  and _30188_ (_04762_, _04761_, _04759_);
  or _30189_ (_04763_, _04549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _30190_ (_04764_, _04763_, _04612_);
  and _30191_ (_04765_, _04764_, _04580_);
  or _30192_ (_04766_, _04765_, _04762_);
  or _30193_ (_04767_, _04766_, _04575_);
  or _30194_ (_04768_, _04576_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _30195_ (_04769_, _04768_, _04556_);
  and _30196_ (_04770_, _04769_, _04767_);
  or _30197_ (_01212_, _04770_, _04758_);
  and _30198_ (_04771_, _04566_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _30199_ (_04772_, _04771_, _04614_);
  or _30200_ (_04773_, _04772_, _04723_);
  and _30201_ (_04774_, _04773_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _30202_ (_04775_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _04583_);
  nand _30203_ (_04776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _30204_ (_04777_, _04776_, _04720_);
  or _30205_ (_04778_, _04777_, _04775_);
  or _30206_ (_04779_, _04778_, _04774_);
  and _30207_ (_01214_, _04779_, _25365_);
  not _30208_ (_04780_, _04724_);
  and _30209_ (_04781_, _04780_, _04606_);
  or _30210_ (_04782_, _04772_, _04721_);
  and _30211_ (_04783_, _04556_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _30212_ (_04784_, _04783_, _04782_);
  or _30213_ (_01216_, _04784_, _04781_);
  or _30214_ (_04785_, _04599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _30215_ (_04786_, _04599_, _04544_);
  and _30216_ (_04787_, _04786_, _25365_);
  and _30217_ (_01218_, _04787_, _04785_);
  or _30218_ (_04788_, _04601_, _04564_);
  or _30219_ (_04789_, _04570_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _30220_ (_04790_, _04789_, _25365_);
  and _30221_ (_01220_, _04790_, _04788_);
  and _30222_ (_04791_, _04601_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _30223_ (_04793_, _04590_, _04596_);
  and _30224_ (_04794_, _04793_, _04570_);
  or _30225_ (_04795_, _04794_, _04791_);
  and _30226_ (_01222_, _04795_, _25365_);
  and _30227_ (_04796_, _04603_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _30228_ (_04797_, _04596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _30229_ (_04798_, _04797_, _04602_);
  or _30230_ (_04799_, _04798_, _04796_);
  and _30231_ (_01224_, _04799_, _25365_);
  and _30232_ (_04800_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _04583_);
  and _30233_ (_04801_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _30234_ (_04802_, _04801_, _04800_);
  and _30235_ (_01226_, _04802_, _25365_);
  and _30236_ (_04803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _04583_);
  and _30237_ (_04804_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _30238_ (_04805_, _04804_, _04803_);
  and _30239_ (_01228_, _04805_, _25365_);
  and _30240_ (_04806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _04583_);
  and _30241_ (_04807_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _30242_ (_04808_, _04807_, _04806_);
  and _30243_ (_01230_, _04808_, _25365_);
  and _30244_ (_04809_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _04583_);
  and _30245_ (_04810_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _30246_ (_04811_, _04810_, _04809_);
  and _30247_ (_01232_, _04811_, _25365_);
  and _30248_ (_04812_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _04583_);
  and _30249_ (_04813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _30250_ (_04814_, _04813_, _04812_);
  and _30251_ (_01234_, _04814_, _25365_);
  and _30252_ (_04815_, _04556_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _30253_ (_01236_, _04815_, _04758_);
  and _30254_ (_04816_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _30255_ (_04817_, _04816_, _04775_);
  and _30256_ (_01238_, _04817_, _25365_);
  nor _30257_ (_04818_, _04659_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _30258_ (_04819_, _04818_, _04695_);
  and _30259_ (_01240_, _04819_, _04678_);
  nor _30260_ (_04820_, _04695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _30261_ (_04821_, _04820_, _04696_);
  and _30262_ (_01242_, _04821_, _04678_);
  nor _30263_ (_04822_, _04696_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _30264_ (_04823_, _04822_, _04697_);
  and _30265_ (_01244_, _04823_, _04678_);
  or _30266_ (_04824_, _04660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _30267_ (_04825_, _04661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _30268_ (_04826_, _04825_, _04824_);
  and _30269_ (_04827_, _04826_, _04669_);
  and _30270_ (_04828_, _04653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _30271_ (_04829_, _04828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _30272_ (_04830_, _04829_, _04642_);
  nor _30273_ (_04831_, _04830_, _04827_);
  nor _30274_ (_04832_, _04831_, _04677_);
  nor _30275_ (_04833_, _04547_, _02259_);
  and _30276_ (_04834_, _04833_, _04677_);
  or _30277_ (_04835_, _04834_, _04832_);
  and _30278_ (_01246_, _04835_, _25365_);
  not _30279_ (_04836_, _04701_);
  and _30280_ (_04837_, _04836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _30281_ (_04838_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _30282_ (_04839_, _04838_, _04837_);
  and _30283_ (_04840_, _04839_, _04678_);
  or _30284_ (_04841_, _04547_, _02251_);
  nand _30285_ (_04842_, _04547_, _02259_);
  and _30286_ (_04843_, _04842_, _04681_);
  and _30287_ (_04844_, _04843_, _04841_);
  or _30288_ (_01248_, _04844_, _04840_);
  nor _30289_ (_04845_, _04701_, _04648_);
  and _30290_ (_04846_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _30291_ (_04847_, _04846_, _04845_);
  and _30292_ (_04848_, _04847_, _04678_);
  or _30293_ (_04849_, _04547_, _02236_);
  or _30294_ (_04850_, _04546_, _02251_);
  and _30295_ (_04851_, _04850_, _04681_);
  and _30296_ (_04852_, _04851_, _04849_);
  or _30297_ (_01250_, _04852_, _04848_);
  nor _30298_ (_04853_, _04701_, _04644_);
  and _30299_ (_04854_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _30300_ (_04855_, _04854_, _04853_);
  and _30301_ (_04856_, _04855_, _04678_);
  or _30302_ (_04857_, _04546_, _02236_);
  or _30303_ (_04858_, _04547_, _02220_);
  and _30304_ (_04859_, _04858_, _04681_);
  and _30305_ (_04860_, _04859_, _04857_);
  or _30306_ (_01252_, _04860_, _04856_);
  and _30307_ (_04861_, _04836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _30308_ (_04862_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or _30309_ (_04863_, _04862_, _04861_);
  and _30310_ (_04864_, _04863_, _04678_);
  or _30311_ (_04865_, _04546_, _02220_);
  nand _30312_ (_04866_, _04546_, _02204_);
  and _30313_ (_04867_, _04866_, _04681_);
  and _30314_ (_04868_, _04867_, _04865_);
  or _30315_ (_01254_, _04868_, _04864_);
  and _30316_ (_04869_, _04836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _30317_ (_04870_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _30318_ (_04871_, _04870_, _04869_);
  and _30319_ (_04872_, _04871_, _04678_);
  nand _30320_ (_04873_, _04546_, _02190_);
  nand _30321_ (_04874_, _04547_, _02204_);
  and _30322_ (_04875_, _04874_, _04681_);
  and _30323_ (_04877_, _04875_, _04873_);
  or _30324_ (_01256_, _04877_, _04872_);
  and _30325_ (_04878_, _04836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _30326_ (_04879_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or _30327_ (_04880_, _04879_, _04878_);
  and _30328_ (_04881_, _04880_, _04678_);
  nand _30329_ (_04882_, _04546_, _02177_);
  nand _30330_ (_04883_, _04547_, _02190_);
  and _30331_ (_04884_, _04883_, _04681_);
  and _30332_ (_04885_, _04884_, _04882_);
  or _30333_ (_01258_, _04885_, _04881_);
  and _30334_ (_04886_, _04836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _30335_ (_04887_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _30336_ (_04888_, _04887_, _04886_);
  and _30337_ (_04889_, _04888_, _04678_);
  nand _30338_ (_04890_, _04546_, _02280_);
  nand _30339_ (_04891_, _04547_, _02177_);
  and _30340_ (_04892_, _04891_, _04681_);
  and _30341_ (_04893_, _04892_, _04890_);
  or _30342_ (_01260_, _04893_, _04889_);
  and _30343_ (_04894_, _04677_, _04547_);
  nand _30344_ (_04895_, _04894_, _02280_);
  and _30345_ (_04896_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _30346_ (_04897_, _04836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _30347_ (_04898_, _04897_, _04896_);
  or _30348_ (_04899_, _04898_, _04677_);
  and _30349_ (_04900_, _04899_, _25365_);
  and _30350_ (_01262_, _04900_, _04895_);
  and _30351_ (_04901_, _04836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _30352_ (_04902_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _30353_ (_04903_, _04902_, _04901_);
  and _30354_ (_04904_, _04903_, _04678_);
  or _30355_ (_04905_, _04534_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _30356_ (_04906_, _04905_, _04547_);
  and _30357_ (_04907_, _04906_, _04681_);
  or _30358_ (_01264_, _04907_, _04904_);
  nand _30359_ (_04908_, _04705_, _02259_);
  or _30360_ (_04909_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _30361_ (_04910_, _04909_, _25365_);
  and _30362_ (_01266_, _04910_, _04908_);
  or _30363_ (_04911_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _30364_ (_04912_, _04911_, _25365_);
  not _30365_ (_04913_, _04705_);
  or _30366_ (_04914_, _04913_, _02251_);
  and _30367_ (_01268_, _04914_, _04912_);
  or _30368_ (_04915_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _30369_ (_04916_, _04915_, _25365_);
  or _30370_ (_04917_, _04913_, _02236_);
  and _30371_ (_01270_, _04917_, _04916_);
  or _30372_ (_04918_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _30373_ (_04919_, _04918_, _25365_);
  or _30374_ (_04920_, _04913_, _02220_);
  and _30375_ (_01272_, _04920_, _04919_);
  or _30376_ (_04921_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _30377_ (_04922_, _04921_, _25365_);
  nand _30378_ (_04923_, _04705_, _02204_);
  and _30379_ (_01274_, _04923_, _04922_);
  or _30380_ (_04924_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _30381_ (_04925_, _04924_, _25365_);
  nand _30382_ (_04926_, _04705_, _02190_);
  and _30383_ (_01276_, _04926_, _04925_);
  or _30384_ (_04927_, _04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _30385_ (_04928_, _04927_, _25365_);
  nand _30386_ (_04929_, _04705_, _02177_);
  and _30387_ (_01278_, _04929_, _04928_);
  nand _30388_ (_04930_, _01289_, _00860_);
  or _30389_ (_04931_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _30390_ (_04932_, _04931_, _04710_);
  and _30391_ (_04933_, _04932_, _04930_);
  not _30392_ (_04934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _30393_ (_04935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _04934_);
  or _30394_ (_04936_, _04935_, _04546_);
  nor _30395_ (_04937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _30396_ (_04938_, _04937_, _04936_);
  nor _30397_ (_04939_, _04938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _30398_ (_04940_, _04939_, _04710_);
  or _30399_ (_04941_, _04940_, _04713_);
  or _30400_ (_04942_, _04941_, _04933_);
  nand _30401_ (_04943_, _04713_, _02259_);
  and _30402_ (_04944_, _04943_, _25365_);
  and _30403_ (_01280_, _04944_, _04942_);
  and _30404_ (_04945_, _02689_, _01344_);
  not _30405_ (_04946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _30406_ (_04947_, _02689_, _04946_);
  nand _30407_ (_04948_, _04947_, _04710_);
  or _30408_ (_04949_, _04948_, _04945_);
  or _30409_ (_04950_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _30410_ (_04951_, _04950_, _04710_);
  and _30411_ (_04952_, _04951_, _04949_);
  or _30412_ (_04953_, _04952_, _04713_);
  or _30413_ (_04954_, _04714_, _02251_);
  and _30414_ (_04955_, _04954_, _25365_);
  and _30415_ (_01282_, _04955_, _04953_);
  not _30416_ (_04956_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not _30417_ (_04957_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _30418_ (_04958_, _04559_, _04957_);
  nor _30419_ (_04959_, _04958_, _04956_);
  and _30420_ (_04960_, _04958_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _30421_ (_04961_, _04960_, _04959_);
  or _30422_ (_04962_, _04961_, _04710_);
  or _30423_ (_04963_, _01468_, _04956_);
  nand _30424_ (_04964_, _04963_, _04710_);
  or _30425_ (_04965_, _04964_, _01470_);
  and _30426_ (_04966_, _04965_, _04962_);
  or _30427_ (_04967_, _04966_, _04713_);
  or _30428_ (_04968_, _04714_, _02236_);
  and _30429_ (_04969_, _04968_, _25365_);
  and _30430_ (_01284_, _04969_, _04967_);
  and _30431_ (_04970_, _04710_, _01530_);
  nand _30432_ (_04971_, _04970_, _01289_);
  or _30433_ (_04972_, _04970_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _30434_ (_04973_, _04972_, _04714_);
  and _30435_ (_04974_, _04973_, _04971_);
  and _30436_ (_04975_, _04713_, _02220_);
  or _30437_ (_04976_, _04975_, _04974_);
  and _30438_ (_01286_, _04976_, _25365_);
  and _30439_ (_04977_, _04710_, _01597_);
  nand _30440_ (_04978_, _04977_, _01289_);
  or _30441_ (_04979_, _04977_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _30442_ (_04980_, _04979_, _04714_);
  and _30443_ (_04981_, _04980_, _04978_);
  nor _30444_ (_04982_, _04714_, _02204_);
  or _30445_ (_04983_, _04982_, _04981_);
  and _30446_ (_01288_, _04983_, _25365_);
  and _30447_ (_04984_, _04710_, _01680_);
  nand _30448_ (_04985_, _04984_, _01289_);
  or _30449_ (_04986_, _04984_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _30450_ (_04987_, _04986_, _04714_);
  and _30451_ (_04988_, _04987_, _04985_);
  nor _30452_ (_04989_, _04714_, _02190_);
  or _30453_ (_04990_, _04989_, _04988_);
  and _30454_ (_01290_, _04990_, _25365_);
  and _30455_ (_04991_, _04710_, _01745_);
  nand _30456_ (_04992_, _04991_, _01289_);
  or _30457_ (_04993_, _04991_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _30458_ (_04994_, _04993_, _04714_);
  and _30459_ (_04995_, _04994_, _04992_);
  nor _30460_ (_04996_, _04714_, _02177_);
  or _30461_ (_04997_, _04996_, _04995_);
  and _30462_ (_01292_, _04997_, _25365_);
  and _30463_ (_01625_, t2_i, _25365_);
  nor _30464_ (_04998_, t2_i, rst);
  and _30465_ (_01628_, _04998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand _30466_ (_04999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _25365_);
  nor _30467_ (_01631_, _04999_, t2ex_i);
  and _30468_ (_01634_, t2ex_i, _25365_);
  and _30469_ (_05000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _30470_ (_05001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _30471_ (_05002_, _05001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _30472_ (_05003_, _05002_, _05000_);
  not _30473_ (_05004_, _05003_);
  and _30474_ (_05005_, _05004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _30475_ (_05006_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor _30476_ (_05007_, _05006_, _05005_);
  and _30477_ (_05008_, _02159_, _02681_);
  and _30478_ (_05009_, _05008_, _03471_);
  nor _30479_ (_05010_, _05009_, _05007_);
  and _30480_ (_05011_, _00858_, _01466_);
  and _30481_ (_05012_, _03533_, _05011_);
  and _30482_ (_05013_, _05008_, _05012_);
  and _30483_ (_05014_, _05013_, _01190_);
  not _30484_ (_05015_, _05014_);
  nor _30485_ (_05016_, _05015_, _02280_);
  or _30486_ (_05017_, _05016_, _05010_);
  and _30487_ (_05018_, _05008_, _03343_);
  not _30488_ (_05019_, _05018_);
  and _30489_ (_05020_, _05019_, _05017_);
  and _30490_ (_05021_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _30491_ (_05022_, _05021_, _05020_);
  and _30492_ (_01637_, _05022_, _25365_);
  nand _30493_ (_05023_, _05018_, _02280_);
  nor _30494_ (_05024_, _05009_, _05004_);
  or _30495_ (_05025_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _30496_ (_05026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _30497_ (_05027_, _05024_, _05026_);
  and _30498_ (_05028_, _05027_, _05025_);
  or _30499_ (_05029_, _05028_, _05018_);
  and _30500_ (_05030_, _05029_, _25365_);
  and _30501_ (_01640_, _05030_, _05023_);
  and _30502_ (_05031_, _05008_, _01680_);
  and _30503_ (_05032_, _05031_, _03342_);
  and _30504_ (_05033_, _05008_, _03431_);
  nor _30505_ (_05034_, _05033_, _05032_);
  not _30506_ (_05035_, _05001_);
  or _30507_ (_05036_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _30508_ (_05037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _30509_ (_05038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _05037_);
  and _30510_ (_05039_, _05038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _30511_ (_05040_, _05039_, _05036_);
  and _30512_ (_05041_, _05040_, _05035_);
  and _30513_ (_05042_, _05041_, _05034_);
  and _30514_ (_05043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _30515_ (_05044_, _05043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _30516_ (_05045_, _05044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _30517_ (_05046_, _05045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _30518_ (_05047_, _05046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _30519_ (_05048_, _05047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _30520_ (_05049_, _05048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _30521_ (_05050_, _05049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _30522_ (_05051_, _05050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _30523_ (_05052_, _05051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _30524_ (_05053_, _05052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _30525_ (_05054_, _05053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _30526_ (_05055_, _05054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _30527_ (_05056_, _05055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _30528_ (_05057_, _05056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _30529_ (_05058_, _05057_);
  nand _30530_ (_05059_, _05058_, _05042_);
  or _30531_ (_05060_, _05042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _30532_ (_05061_, _05060_, _25365_);
  and _30533_ (_01643_, _05061_, _05059_);
  nand _30534_ (_05062_, _05033_, _02280_);
  not _30535_ (_05063_, _05032_);
  not _30536_ (_05064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _30537_ (_05065_, _05000_, _05064_);
  and _30538_ (_05066_, _05065_, _05001_);
  and _30539_ (_05067_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not _30540_ (_05068_, _05066_);
  not _30541_ (_05069_, _05002_);
  and _30542_ (_05070_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _30543_ (_05071_, _05057_, _05040_);
  and _30544_ (_05072_, _05071_, _05070_);
  and _30545_ (_05073_, _05048_, _05040_);
  or _30546_ (_05074_, _05073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _30547_ (_05075_, _05073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _30548_ (_05076_, _05075_, _05074_);
  or _30549_ (_05077_, _05076_, _05072_);
  and _30550_ (_05078_, _05077_, _05068_);
  or _30551_ (_05079_, _05078_, _05067_);
  or _30552_ (_05080_, _05079_, _05033_);
  and _30553_ (_05081_, _05080_, _05063_);
  and _30554_ (_05082_, _05081_, _05062_);
  and _30555_ (_05083_, _05032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _30556_ (_05084_, _05083_, _05082_);
  and _30557_ (_01646_, _05084_, _25365_);
  nand _30558_ (_05085_, _05032_, _02280_);
  nor _30559_ (_05086_, _05066_, _05026_);
  and _30560_ (_05087_, _05068_, _05040_);
  and _30561_ (_05088_, _05087_, _05056_);
  or _30562_ (_05089_, _05088_, _05086_);
  nand _30563_ (_05090_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _30564_ (_05091_, _05090_, _05071_);
  and _30565_ (_05092_, _05091_, _05089_);
  nand _30566_ (_05093_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _30567_ (_05094_, _05093_, _05034_);
  or _30568_ (_05095_, _05094_, _05092_);
  nand _30569_ (_05096_, _05033_, _05026_);
  and _30570_ (_05097_, _05096_, _25365_);
  and _30571_ (_05098_, _05097_, _05095_);
  and _30572_ (_01649_, _05098_, _05085_);
  and _30573_ (_05099_, _05001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _30574_ (_05100_, _05099_, _05088_);
  nand _30575_ (_05101_, _05100_, _05034_);
  or _30576_ (_05102_, _05034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _30577_ (_05103_, _05102_, _25365_);
  and _30578_ (_01652_, _05103_, _05101_);
  or _30579_ (_05104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _30580_ (_05105_, _04004_, _02664_);
  or _30581_ (_05106_, _05105_, _05104_);
  nand _30582_ (_05107_, _02667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _30583_ (_05108_, _05107_, _05105_);
  or _30584_ (_05109_, _05108_, _02669_);
  and _30585_ (_05110_, _05109_, _05106_);
  and _30586_ (_05111_, _05008_, _04000_);
  or _30587_ (_05112_, _05111_, _05110_);
  nand _30588_ (_05113_, _05111_, _02280_);
  and _30589_ (_05114_, _05113_, _25365_);
  and _30590_ (_01655_, _05114_, _05112_);
  or _30591_ (_05115_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not _30592_ (_05116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _30593_ (_05117_, _05003_, _05116_);
  and _30594_ (_05118_, _05117_, _05115_);
  or _30595_ (_05119_, _05118_, _05009_);
  nand _30596_ (_05120_, _05009_, _02259_);
  and _30597_ (_05121_, _05120_, _05119_);
  or _30598_ (_05122_, _05121_, _05018_);
  not _30599_ (_05123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _30600_ (_05124_, _05018_, _05123_);
  and _30601_ (_05125_, _05124_, _25365_);
  and _30602_ (_02181_, _05125_, _05122_);
  not _30603_ (_05126_, _05009_);
  or _30604_ (_05127_, _05126_, _02251_);
  not _30605_ (_05128_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nor _30606_ (_05129_, _05003_, _05128_);
  and _30607_ (_05130_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _30608_ (_05131_, _05130_, _05129_);
  or _30609_ (_05132_, _05131_, _05009_);
  and _30610_ (_05133_, _05132_, _05127_);
  or _30611_ (_05134_, _05133_, _05018_);
  nand _30612_ (_05135_, _05018_, _05128_);
  and _30613_ (_05136_, _05135_, _25365_);
  and _30614_ (_02183_, _05136_, _05134_);
  and _30615_ (_05137_, _05004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _30616_ (_05138_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _30617_ (_05139_, _05138_, _05137_);
  nor _30618_ (_05140_, _05139_, _05009_);
  and _30619_ (_05141_, _05014_, _02236_);
  or _30620_ (_05142_, _05141_, _05140_);
  and _30621_ (_05143_, _05142_, _05019_);
  and _30622_ (_05144_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _30623_ (_05145_, _05144_, _05143_);
  and _30624_ (_02185_, _05145_, _25365_);
  and _30625_ (_05146_, _05004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _30626_ (_05147_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _30627_ (_05148_, _05147_, _05146_);
  nor _30628_ (_05149_, _05148_, _05009_);
  and _30629_ (_05150_, _05014_, _02220_);
  or _30630_ (_05151_, _05150_, _05149_);
  and _30631_ (_05152_, _05151_, _05019_);
  and _30632_ (_05153_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _30633_ (_05154_, _05153_, _05152_);
  and _30634_ (_02187_, _05154_, _25365_);
  and _30635_ (_05155_, _05004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _30636_ (_05156_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _30637_ (_05157_, _05156_, _05155_);
  nor _30638_ (_05158_, _05157_, _05009_);
  nor _30639_ (_05159_, _05015_, _02204_);
  or _30640_ (_05160_, _05159_, _05158_);
  and _30641_ (_05161_, _05160_, _05019_);
  and _30642_ (_05162_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _30643_ (_05163_, _05162_, _05161_);
  and _30644_ (_02189_, _05163_, _25365_);
  and _30645_ (_05164_, _05004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _30646_ (_05165_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _30647_ (_05166_, _05165_, _05164_);
  nor _30648_ (_05167_, _05166_, _05009_);
  nor _30649_ (_05168_, _05015_, _02190_);
  or _30650_ (_05169_, _05168_, _05167_);
  and _30651_ (_05170_, _05169_, _05019_);
  and _30652_ (_05171_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _30653_ (_05172_, _05171_, _05170_);
  and _30654_ (_02191_, _05172_, _25365_);
  not _30655_ (_05173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _30656_ (_05174_, _05003_, _05173_);
  and _30657_ (_05175_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _30658_ (_05176_, _05175_, _05174_);
  nor _30659_ (_05177_, _05176_, _05009_);
  nor _30660_ (_05178_, _05015_, _02177_);
  or _30661_ (_05179_, _05178_, _05177_);
  and _30662_ (_05180_, _05179_, _05019_);
  and _30663_ (_05181_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _30664_ (_05182_, _05181_, _05180_);
  and _30665_ (_02193_, _05182_, _25365_);
  or _30666_ (_05183_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _30667_ (_05184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _30668_ (_05185_, _05024_, _05184_);
  and _30669_ (_05186_, _05185_, _05183_);
  or _30670_ (_05187_, _05186_, _05018_);
  nand _30671_ (_05188_, _05018_, _02259_);
  and _30672_ (_05189_, _05188_, _25365_);
  and _30673_ (_02195_, _05189_, _05187_);
  not _30674_ (_05190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _30675_ (_05191_, _05024_, _05190_);
  and _30676_ (_05192_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _30677_ (_05193_, _05192_, _05191_);
  and _30678_ (_05194_, _05193_, _05019_);
  and _30679_ (_05195_, _05018_, _02251_);
  or _30680_ (_05196_, _05195_, _05194_);
  and _30681_ (_02197_, _05196_, _25365_);
  or _30682_ (_05197_, _05019_, _02236_);
  not _30683_ (_05198_, _05024_);
  and _30684_ (_05199_, _05198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _30685_ (_05200_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _30686_ (_05201_, _05200_, _05199_);
  or _30687_ (_05202_, _05201_, _05018_);
  and _30688_ (_05203_, _05202_, _25365_);
  and _30689_ (_02199_, _05203_, _05197_);
  or _30690_ (_05204_, _05019_, _02220_);
  and _30691_ (_05205_, _05198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _30692_ (_05206_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _30693_ (_05207_, _05206_, _05205_);
  or _30694_ (_05208_, _05207_, _05018_);
  and _30695_ (_05209_, _05208_, _25365_);
  and _30696_ (_02201_, _05209_, _05204_);
  nand _30697_ (_05210_, _05018_, _02204_);
  and _30698_ (_05211_, _05198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _30699_ (_05212_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _30700_ (_05213_, _05212_, _05211_);
  or _30701_ (_05214_, _05213_, _05018_);
  and _30702_ (_05215_, _05214_, _25365_);
  and _30703_ (_02203_, _05215_, _05210_);
  nand _30704_ (_05216_, _05018_, _02190_);
  not _30705_ (_05217_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor _30706_ (_05218_, _05024_, _05217_);
  and _30707_ (_05219_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _30708_ (_05220_, _05219_, _05218_);
  or _30709_ (_05221_, _05220_, _05018_);
  and _30710_ (_05222_, _05221_, _25365_);
  and _30711_ (_02205_, _05222_, _05216_);
  nand _30712_ (_05223_, _05018_, _02177_);
  not _30713_ (_05224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _30714_ (_05225_, _05024_, _05224_);
  and _30715_ (_05226_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _30716_ (_05227_, _05226_, _05225_);
  or _30717_ (_05228_, _05227_, _05018_);
  and _30718_ (_05229_, _05228_, _25365_);
  and _30719_ (_02207_, _05229_, _05223_);
  and _30720_ (_05230_, _05040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _30721_ (_05231_, _05002_, _05123_);
  nand _30722_ (_05232_, _05231_, _05057_);
  nand _30723_ (_05233_, _05232_, _05230_);
  or _30724_ (_05234_, _05040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _30725_ (_05235_, _05234_, _05068_);
  and _30726_ (_05236_, _05235_, _05233_);
  nand _30727_ (_05237_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _30728_ (_05238_, _05237_, _05034_);
  or _30729_ (_05239_, _05238_, _05236_);
  nand _30730_ (_05240_, _05032_, _05116_);
  nand _30731_ (_05241_, _05033_, _02259_);
  and _30732_ (_05242_, _05241_, _25365_);
  and _30733_ (_05243_, _05242_, _05240_);
  and _30734_ (_02209_, _05243_, _05239_);
  nor _30735_ (_05244_, _05002_, _05128_);
  and _30736_ (_05245_, _05244_, _05087_);
  and _30737_ (_05246_, _05245_, _05057_);
  and _30738_ (_05247_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  not _30739_ (_05248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor _30740_ (_05249_, _05230_, _05248_);
  and _30741_ (_05250_, _05230_, _05248_);
  or _30742_ (_05251_, _05250_, _05249_);
  and _30743_ (_05252_, _05251_, _05068_);
  nor _30744_ (_05253_, _05252_, _05247_);
  nand _30745_ (_05254_, _05253_, _05034_);
  or _30746_ (_05255_, _05254_, _05246_);
  not _30747_ (_05256_, _05033_);
  or _30748_ (_05257_, _05256_, _02251_);
  nand _30749_ (_05258_, _05032_, _05248_);
  and _30750_ (_05259_, _05258_, _25365_);
  and _30751_ (_05260_, _05259_, _05257_);
  and _30752_ (_02211_, _05260_, _05255_);
  and _30753_ (_05261_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _30754_ (_05262_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _30755_ (_05263_, _05262_, _05071_);
  nand _30756_ (_05264_, _05043_, _05040_);
  nor _30757_ (_05265_, _05264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _30758_ (_05266_, _05264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _30759_ (_05267_, _05266_, _05265_);
  or _30760_ (_05268_, _05267_, _05263_);
  and _30761_ (_05269_, _05268_, _05068_);
  or _30762_ (_05270_, _05269_, _05261_);
  or _30763_ (_05271_, _05270_, _05033_);
  or _30764_ (_05272_, _05256_, _02236_);
  and _30765_ (_05273_, _05272_, _05063_);
  and _30766_ (_05274_, _05273_, _05271_);
  and _30767_ (_05275_, _05032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _30768_ (_05276_, _05275_, _05274_);
  and _30769_ (_02213_, _05276_, _25365_);
  and _30770_ (_05277_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _30771_ (_05278_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _30772_ (_05279_, _05278_, _05071_);
  nand _30773_ (_05280_, _05044_, _05040_);
  nor _30774_ (_05281_, _05280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _30775_ (_05282_, _05280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _30776_ (_05283_, _05282_, _05281_);
  or _30777_ (_05284_, _05283_, _05279_);
  and _30778_ (_05285_, _05284_, _05068_);
  or _30779_ (_05286_, _05285_, _05277_);
  or _30780_ (_05287_, _05286_, _05033_);
  or _30781_ (_05288_, _05256_, _02220_);
  and _30782_ (_05289_, _05288_, _05063_);
  and _30783_ (_05290_, _05289_, _05287_);
  and _30784_ (_05291_, _05032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _30785_ (_05292_, _05291_, _05290_);
  and _30786_ (_02215_, _05292_, _25365_);
  and _30787_ (_05293_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _30788_ (_05294_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _30789_ (_05295_, _05294_, _05071_);
  nand _30790_ (_05296_, _05045_, _05040_);
  nor _30791_ (_05297_, _05296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _30792_ (_05298_, _05296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _30793_ (_05299_, _05298_, _05297_);
  or _30794_ (_05300_, _05299_, _05295_);
  and _30795_ (_05301_, _05300_, _05068_);
  or _30796_ (_05302_, _05301_, _05293_);
  or _30797_ (_05303_, _05302_, _05033_);
  nand _30798_ (_05304_, _05033_, _02204_);
  and _30799_ (_05305_, _05304_, _05063_);
  and _30800_ (_05306_, _05305_, _05303_);
  and _30801_ (_05307_, _05032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _30802_ (_05308_, _05307_, _05306_);
  and _30803_ (_02217_, _05308_, _25365_);
  and _30804_ (_05309_, _05066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _30805_ (_05310_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _30806_ (_05311_, _05310_, _05071_);
  nand _30807_ (_05312_, _05046_, _05040_);
  nor _30808_ (_05313_, _05312_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _30809_ (_05314_, _05312_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _30810_ (_05315_, _05314_, _05313_);
  or _30811_ (_05316_, _05315_, _05311_);
  and _30812_ (_05317_, _05316_, _05068_);
  or _30813_ (_05318_, _05317_, _05309_);
  and _30814_ (_05319_, _05318_, _05256_);
  nor _30815_ (_05320_, _05256_, _02190_);
  or _30816_ (_05321_, _05320_, _05032_);
  or _30817_ (_05322_, _05321_, _05319_);
  or _30818_ (_05323_, _05063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _30819_ (_05324_, _05323_, _25365_);
  and _30820_ (_02219_, _05324_, _05322_);
  nor _30821_ (_05325_, _05256_, _02177_);
  nor _30822_ (_05326_, _05002_, _05173_);
  and _30823_ (_05327_, _05326_, _05071_);
  and _30824_ (_05328_, _05047_, _05040_);
  nor _30825_ (_05329_, _05328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _30826_ (_05330_, _05329_, _05073_);
  or _30827_ (_05331_, _05330_, _05066_);
  or _30828_ (_05332_, _05331_, _05327_);
  nand _30829_ (_05333_, _05066_, _05173_);
  and _30830_ (_05334_, _05333_, _05034_);
  and _30831_ (_05335_, _05334_, _05332_);
  and _30832_ (_05336_, _05032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _30833_ (_05337_, _05336_, _05335_);
  or _30834_ (_05338_, _05337_, _05325_);
  and _30835_ (_02221_, _05338_, _25365_);
  not _30836_ (_05339_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _30837_ (_05340_, _05002_, _05339_);
  and _30838_ (_05341_, _05340_, _05071_);
  and _30839_ (_05342_, _05049_, _05040_);
  or _30840_ (_05343_, _05342_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _30841_ (_05344_, _05342_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _30842_ (_05345_, _05344_, _05343_);
  or _30843_ (_05346_, _05345_, _05066_);
  or _30844_ (_05347_, _05346_, _05341_);
  nand _30845_ (_05348_, _05066_, _05339_);
  and _30846_ (_05349_, _05348_, _05034_);
  and _30847_ (_05350_, _05349_, _05347_);
  and _30848_ (_05351_, _05033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _30849_ (_05352_, _05032_, _02260_);
  or _30850_ (_05353_, _05352_, _05351_);
  or _30851_ (_05354_, _05353_, _05350_);
  and _30852_ (_02223_, _05354_, _25365_);
  nor _30853_ (_05355_, _05002_, _05190_);
  and _30854_ (_05356_, _05355_, _05071_);
  and _30855_ (_05357_, _05050_, _05040_);
  or _30856_ (_05358_, _05357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _30857_ (_05359_, _05357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _30858_ (_05360_, _05359_, _05358_);
  or _30859_ (_05361_, _05360_, _05066_);
  or _30860_ (_05362_, _05361_, _05356_);
  not _30861_ (_05363_, _05034_);
  and _30862_ (_05364_, _05066_, _05190_);
  nor _30863_ (_05365_, _05364_, _05363_);
  and _30864_ (_05366_, _05365_, _05362_);
  and _30865_ (_05367_, _05032_, _02251_);
  and _30866_ (_05368_, _05033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _30867_ (_05369_, _05368_, _05367_);
  or _30868_ (_05370_, _05369_, _05366_);
  and _30869_ (_02225_, _05370_, _25365_);
  and _30870_ (_05371_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _30871_ (_05372_, _05371_, _05071_);
  and _30872_ (_05373_, _05051_, _05040_);
  or _30873_ (_05374_, _05373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _30874_ (_05375_, _05373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _30875_ (_05376_, _05375_, _05374_);
  or _30876_ (_05377_, _05376_, _05066_);
  or _30877_ (_05378_, _05377_, _05372_);
  nor _30878_ (_05379_, _05068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _30879_ (_05380_, _05379_, _05363_);
  and _30880_ (_05381_, _05380_, _05378_);
  and _30881_ (_05382_, _05032_, _02236_);
  and _30882_ (_05383_, _05033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _30883_ (_05384_, _05383_, _05382_);
  or _30884_ (_05385_, _05384_, _05381_);
  and _30885_ (_02227_, _05385_, _25365_);
  and _30886_ (_05386_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _30887_ (_05387_, _05386_, _05071_);
  nand _30888_ (_05388_, _05052_, _05040_);
  nor _30889_ (_05389_, _05388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _30890_ (_05390_, _05388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _30891_ (_05391_, _05390_, _05066_);
  or _30892_ (_05392_, _05391_, _05389_);
  or _30893_ (_05393_, _05392_, _05387_);
  or _30894_ (_05394_, _05068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _30895_ (_05395_, _05394_, _05034_);
  and _30896_ (_05396_, _05395_, _05393_);
  and _30897_ (_05397_, _05033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _30898_ (_05398_, _05397_, _05396_);
  and _30899_ (_05399_, _05032_, _02220_);
  or _30900_ (_05400_, _05399_, _05398_);
  and _30901_ (_02229_, _05400_, _25365_);
  and _30902_ (_05401_, _05069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _30903_ (_05402_, _05401_, _05071_);
  nand _30904_ (_05403_, _05053_, _05040_);
  and _30905_ (_05404_, _05403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _30906_ (_05405_, _05403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _30907_ (_05406_, _05405_, _05066_);
  or _30908_ (_05407_, _05406_, _05404_);
  or _30909_ (_05408_, _05407_, _05402_);
  or _30910_ (_05409_, _05068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _30911_ (_05410_, _05409_, _05034_);
  and _30912_ (_05411_, _05410_, _05408_);
  and _30913_ (_05412_, _05033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _30914_ (_05413_, _05412_, _05411_);
  nor _30915_ (_05414_, _05063_, _02204_);
  or _30916_ (_05415_, _05414_, _05413_);
  and _30917_ (_02231_, _05415_, _25365_);
  nor _30918_ (_05416_, _05002_, _05217_);
  nand _30919_ (_05417_, _05416_, _05071_);
  and _30920_ (_05418_, _05054_, _05040_);
  nor _30921_ (_05419_, _05418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _30922_ (_05420_, _05418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _30923_ (_05421_, _05420_, _05419_);
  and _30924_ (_05422_, _05421_, _05068_);
  nand _30925_ (_05423_, _05422_, _05417_);
  and _30926_ (_05424_, _05066_, _05217_);
  nor _30927_ (_05425_, _05424_, _05363_);
  and _30928_ (_05426_, _05425_, _05423_);
  and _30929_ (_05427_, _05033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _30930_ (_05428_, _05427_, _05426_);
  nor _30931_ (_05429_, _05063_, _02190_);
  or _30932_ (_05430_, _05429_, _05428_);
  and _30933_ (_02233_, _05430_, _25365_);
  and _30934_ (_05431_, _05033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _30935_ (_05432_, _05002_, _05224_);
  and _30936_ (_05433_, _05432_, _05071_);
  not _30937_ (_05434_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _30938_ (_05435_, _05055_, _05040_);
  nor _30939_ (_05436_, _05435_, _05434_);
  and _30940_ (_05437_, _05435_, _05434_);
  or _30941_ (_05438_, _05437_, _05066_);
  or _30942_ (_05439_, _05438_, _05436_);
  or _30943_ (_05440_, _05439_, _05433_);
  nand _30944_ (_05441_, _05066_, _05224_);
  and _30945_ (_05442_, _05441_, _05034_);
  and _30946_ (_05443_, _05442_, _05440_);
  or _30947_ (_05444_, _05443_, _05431_);
  nor _30948_ (_05445_, _05063_, _02177_);
  or _30949_ (_05446_, _05445_, _05444_);
  and _30950_ (_02235_, _05446_, _25365_);
  not _30951_ (_05447_, _05111_);
  and _30952_ (_05448_, _05105_, _00860_);
  or _30953_ (_05449_, _05448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _30954_ (_05450_, _05449_, _05447_);
  nand _30955_ (_05451_, _05448_, _01289_);
  and _30956_ (_05452_, _05451_, _05450_);
  and _30957_ (_05453_, _05111_, _02260_);
  or _30958_ (_05454_, _05453_, _05452_);
  and _30959_ (_02237_, _05454_, _25365_);
  and _30960_ (_05455_, _05105_, _02689_);
  or _30961_ (_05456_, _05455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _30962_ (_05457_, _05456_, _05447_);
  nand _30963_ (_05458_, _05455_, _01289_);
  and _30964_ (_05459_, _05458_, _05457_);
  and _30965_ (_05460_, _05111_, _02251_);
  or _30966_ (_05461_, _05460_, _05459_);
  and _30967_ (_02239_, _05461_, _25365_);
  nand _30968_ (_05462_, _05105_, _02998_);
  and _30969_ (_05463_, _05462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _30970_ (_05464_, _05463_, _05111_);
  and _30971_ (_05465_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _30972_ (_05466_, _05465_, _01470_);
  and _30973_ (_05467_, _05466_, _05105_);
  or _30974_ (_05468_, _05467_, _05464_);
  or _30975_ (_05469_, _05447_, _02236_);
  and _30976_ (_05470_, _05469_, _25365_);
  and _30977_ (_02241_, _05470_, _05468_);
  and _30978_ (_05471_, _05105_, _01530_);
  or _30979_ (_05472_, _05471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _30980_ (_05473_, _05472_, _05447_);
  nand _30981_ (_05474_, _05471_, _01289_);
  and _30982_ (_05475_, _05474_, _05473_);
  and _30983_ (_05476_, _05111_, _02220_);
  or _30984_ (_05477_, _05476_, _05475_);
  and _30985_ (_02243_, _05477_, _25365_);
  and _30986_ (_05478_, _05105_, _01597_);
  or _30987_ (_05479_, _05478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _30988_ (_05480_, _05479_, _05447_);
  nand _30989_ (_05481_, _05478_, _01289_);
  and _30990_ (_05482_, _05481_, _05480_);
  nor _30991_ (_05483_, _05447_, _02204_);
  or _30992_ (_05484_, _05483_, _05482_);
  and _30993_ (_02245_, _05484_, _25365_);
  and _30994_ (_05485_, _05105_, _01680_);
  or _30995_ (_05486_, _05485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _30996_ (_05487_, _05486_, _05447_);
  nand _30997_ (_05488_, _05485_, _01289_);
  and _30998_ (_05489_, _05488_, _05487_);
  nor _30999_ (_05490_, _05447_, _02190_);
  or _31000_ (_05491_, _05490_, _05489_);
  and _31001_ (_02247_, _05491_, _25365_);
  not _31002_ (_05492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _31003_ (_05493_, _05000_, _05492_);
  or _31004_ (_05494_, _05493_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _31005_ (_05495_, _05494_, _05105_);
  nand _31006_ (_05496_, _02772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _31007_ (_05497_, _05496_, _05105_);
  or _31008_ (_05498_, _05497_, _02773_);
  and _31009_ (_05499_, _05498_, _05495_);
  or _31010_ (_05500_, _05499_, _05111_);
  nand _31011_ (_05501_, _05111_, _02177_);
  and _31012_ (_05502_, _05501_, _25365_);
  and _31013_ (_02249_, _05502_, _05500_);
  nor _31014_ (_05503_, _02138_, _02088_);
  nand _31015_ (_05504_, _02282_, _05503_);
  not _31016_ (_05505_, _02138_);
  and _31017_ (_05506_, _05505_, _02088_);
  and _31018_ (_05507_, _02745_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _31019_ (_05508_, _05507_, _02740_);
  nor _31020_ (_05509_, _05508_, _00922_);
  and _31021_ (_05510_, _05508_, _00922_);
  or _31022_ (_05511_, _05510_, _05509_);
  not _31023_ (_05512_, _05511_);
  and _31024_ (_05513_, _01876_, _00858_);
  nor _31025_ (_05514_, _01876_, _00858_);
  nor _31026_ (_05515_, _05514_, _05513_);
  and _31027_ (_05516_, _00879_, _00906_);
  not _31028_ (_05517_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _31029_ (_05518_, _01187_, _05517_);
  and _31030_ (_05519_, _05518_, _01471_);
  and _31031_ (_05520_, _05519_, _05516_);
  and _31032_ (_05521_, _05520_, _05515_);
  and _31033_ (_05522_, _05521_, _00892_);
  and _31034_ (_05523_, _02748_, _03985_);
  nor _31035_ (_05524_, _02748_, _03985_);
  nor _31036_ (_05525_, _05524_, _05523_);
  and _31037_ (_05526_, _05525_, _05522_);
  and _31038_ (_05527_, _05526_, _05512_);
  not _31039_ (_05528_, _02748_);
  nor _31040_ (_05529_, _05508_, _01877_);
  and _31041_ (_05530_, _05529_, _05528_);
  nand _31042_ (_05531_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _31043_ (_05532_, _05508_, _01876_);
  and _31044_ (_05533_, _05532_, _05528_);
  nand _31045_ (_05534_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _31046_ (_05535_, _05534_, _05531_);
  and _31047_ (_05536_, _05508_, _01876_);
  and _31048_ (_05537_, _05536_, _05528_);
  nand _31049_ (_05538_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _31050_ (_05539_, _05536_, _02748_);
  nand _31051_ (_05540_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _31052_ (_05541_, _05540_, _05538_);
  and _31053_ (_05542_, _05541_, _05535_);
  and _31054_ (_05543_, _05508_, _01877_);
  and _31055_ (_05544_, _05543_, _02748_);
  nand _31056_ (_05545_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _31057_ (_05546_, _05529_, _02748_);
  nand _31058_ (_05547_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _31059_ (_05548_, _05547_, _05545_);
  and _31060_ (_05549_, _05532_, _02748_);
  nand _31061_ (_05550_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _31062_ (_05551_, _05543_, _05528_);
  nand _31063_ (_05552_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _31064_ (_05553_, _05552_, _05550_);
  and _31065_ (_05554_, _05553_, _05548_);
  and _31066_ (_05555_, _05554_, _05542_);
  nor _31067_ (_05556_, _05555_, _05527_);
  not _31068_ (_05557_, _02280_);
  and _31069_ (_05558_, _05527_, _05557_);
  or _31070_ (_05559_, _05558_, _05556_);
  nand _31071_ (_05560_, _05559_, _05506_);
  nor _31072_ (_05561_, _05505_, _02088_);
  not _31073_ (_05562_, _01760_);
  and _31074_ (_05563_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _31075_ (_05564_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  not _31076_ (_05565_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _31077_ (_05566_, _01789_, _05565_);
  nor _31078_ (_05567_, _05566_, _05564_);
  and _31079_ (_05568_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _31080_ (_05569_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _31081_ (_05570_, _05569_, _05568_);
  and _31082_ (_05571_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _31083_ (_05572_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _31084_ (_05573_, _05572_, _05571_);
  and _31085_ (_05574_, _05573_, _05570_);
  and _31086_ (_05575_, _05574_, _05567_);
  and _31087_ (_05576_, _01768_, _01760_);
  not _31088_ (_05577_, _05576_);
  nor _31089_ (_05578_, _05577_, _05575_);
  nor _31090_ (_05579_, _05578_, _05563_);
  not _31091_ (_05580_, _05579_);
  nand _31092_ (_05581_, _05580_, _05561_);
  and _31093_ (_05582_, _05581_, _02155_);
  and _31094_ (_05583_, _05582_, _05560_);
  and _31095_ (_05584_, _05583_, _05504_);
  not _31096_ (_05585_, _02055_);
  nor _31097_ (_05586_, _05585_, _02009_);
  and _31098_ (_05587_, _02049_, _01987_);
  not _31099_ (_05588_, _05587_);
  and _31100_ (_05589_, _05588_, _02059_);
  and _31101_ (_05590_, _01998_, _02052_);
  nor _31102_ (_05591_, _05590_, _02070_);
  and _31103_ (_05592_, _05591_, _02065_);
  and _31104_ (_05593_, _05592_, _05589_);
  and _31105_ (_05594_, _05593_, _05586_);
  nor _31106_ (_05595_, _05594_, _02140_);
  not _31107_ (_05596_, _05595_);
  not _31108_ (_05597_, _02079_);
  nor _31109_ (_05598_, _05597_, _02032_);
  nor _31110_ (_05599_, _02036_, _02140_);
  nor _31111_ (_05600_, _05599_, _05598_);
  and _31112_ (_05601_, _05600_, _05596_);
  not _31113_ (_05602_, _05601_);
  and _31114_ (_05603_, _05602_, _05584_);
  not _31115_ (_05604_, _05603_);
  and _31116_ (_05605_, _05561_, _02155_);
  and _31117_ (_05606_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _31118_ (_05607_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _31119_ (_05608_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _31120_ (_05609_, _05608_, _05607_);
  and _31121_ (_05610_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not _31122_ (_05611_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _31123_ (_05612_, _01789_, _05611_);
  nor _31124_ (_05613_, _05612_, _05610_);
  and _31125_ (_05614_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _31126_ (_05615_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _31127_ (_05616_, _05615_, _05614_);
  and _31128_ (_05617_, _05616_, _05613_);
  and _31129_ (_05618_, _05617_, _05609_);
  nor _31130_ (_05619_, _05618_, _05577_);
  nor _31131_ (_05620_, _05619_, _05606_);
  not _31132_ (_05621_, _05620_);
  nand _31133_ (_05622_, _05621_, _05605_);
  and _31134_ (_05623_, _05506_, _02155_);
  not _31135_ (_05624_, _05623_);
  and _31136_ (_05625_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _31137_ (_05626_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _31138_ (_05627_, _05626_, _05625_);
  and _31139_ (_05628_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _31140_ (_05629_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _31141_ (_05630_, _05629_, _05628_);
  and _31142_ (_05631_, _05630_, _05627_);
  and _31143_ (_05632_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _31144_ (_05633_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _31145_ (_05634_, _05633_, _05632_);
  and _31146_ (_05635_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _31147_ (_05636_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _31148_ (_05637_, _05636_, _05635_);
  and _31149_ (_05638_, _05637_, _05634_);
  and _31150_ (_05639_, _05638_, _05631_);
  nor _31151_ (_05640_, _05639_, _05527_);
  and _31152_ (_05641_, _05527_, _02220_);
  nor _31153_ (_05642_, _05641_, _05640_);
  or _31154_ (_05643_, _05642_, _05624_);
  and _31155_ (_05644_, _05643_, _05622_);
  and _31156_ (_05645_, _05503_, _02155_);
  not _31157_ (_05646_, _05645_);
  or _31158_ (_05647_, _02308_, _05646_);
  not _31159_ (_05648_, _05508_);
  and _31160_ (_05649_, _02138_, _02088_);
  and _31161_ (_05650_, _05649_, _02155_);
  nand _31162_ (_05651_, _05650_, _05648_);
  and _31163_ (_05652_, _05651_, _05647_);
  and _31164_ (_05653_, _05652_, _05644_);
  or _31165_ (_05654_, _05653_, _05604_);
  and _31166_ (_05655_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _31167_ (_05656_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _31168_ (_05657_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _31169_ (_05658_, _05657_, _05656_);
  and _31170_ (_05659_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not _31171_ (_05660_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _31172_ (_05661_, _01789_, _05660_);
  nor _31173_ (_05662_, _05661_, _05659_);
  and _31174_ (_05663_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _31175_ (_05664_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _31176_ (_05665_, _05664_, _05663_);
  and _31177_ (_05666_, _05665_, _05662_);
  and _31178_ (_05667_, _05666_, _05658_);
  nor _31179_ (_05668_, _05667_, _05577_);
  nor _31180_ (_05669_, _05668_, _05655_);
  not _31181_ (_05670_, _05669_);
  nand _31182_ (_05671_, _05670_, _05605_);
  and _31183_ (_05672_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _31184_ (_05673_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _31185_ (_05674_, _05673_, _05672_);
  and _31186_ (_05675_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _31187_ (_05676_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _31188_ (_05677_, _05676_, _05675_);
  and _31189_ (_05678_, _05677_, _05674_);
  and _31190_ (_05679_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _31191_ (_05680_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor _31192_ (_05681_, _05680_, _05679_);
  and _31193_ (_05682_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _31194_ (_05683_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _31195_ (_05684_, _05683_, _05682_);
  and _31196_ (_05685_, _05684_, _05681_);
  and _31197_ (_05686_, _05685_, _05678_);
  nor _31198_ (_05687_, _05686_, _05527_);
  and _31199_ (_05688_, _05527_, _02260_);
  nor _31200_ (_05689_, _05688_, _05687_);
  or _31201_ (_05690_, _05689_, _05624_);
  and _31202_ (_05691_, _05690_, _05671_);
  or _31203_ (_05704_, _02290_, _05646_);
  nand _31204_ (_05718_, _05650_, _01876_);
  and _31205_ (_05719_, _05718_, _05704_);
  and _31206_ (_05720_, _05719_, _05691_);
  or _31207_ (_05721_, _05720_, _05602_);
  nand _31208_ (_05722_, _05721_, _05654_);
  and _31209_ (_05723_, _00906_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _31210_ (_05724_, _05723_, _00922_);
  nor _31211_ (_05725_, _00858_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _31212_ (_05726_, _05725_, _05724_);
  nor _31213_ (_05727_, _05726_, _05722_);
  and _31214_ (_05728_, _05726_, _05722_);
  nor _31215_ (_05729_, _05728_, _05727_);
  and _31216_ (_05730_, _05650_, _05528_);
  and _31217_ (_05731_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _31218_ (_05732_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  not _31219_ (_05733_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _31220_ (_05734_, _01789_, _05733_);
  nor _31221_ (_05735_, _05734_, _05732_);
  and _31222_ (_05736_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _31223_ (_05737_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _31224_ (_05738_, _05737_, _05736_);
  and _31225_ (_05739_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _31226_ (_05740_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _31227_ (_05741_, _05740_, _05739_);
  and _31228_ (_05742_, _05741_, _05738_);
  and _31229_ (_05743_, _05742_, _05735_);
  nor _31230_ (_05744_, _05743_, _05577_);
  nor _31231_ (_05745_, _05744_, _05731_);
  not _31232_ (_05746_, _05745_);
  and _31233_ (_05747_, _05746_, _05605_);
  nor _31234_ (_05748_, _05747_, _05730_);
  and _31235_ (_05749_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _31236_ (_05750_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor _31237_ (_05751_, _05750_, _05749_);
  and _31238_ (_05752_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _31239_ (_05753_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _31240_ (_05754_, _05753_, _05752_);
  and _31241_ (_05755_, _05754_, _05751_);
  and _31242_ (_05756_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _31243_ (_05757_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _31244_ (_05758_, _05757_, _05756_);
  and _31245_ (_05759_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _31246_ (_05760_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _31247_ (_05761_, _05760_, _05759_);
  and _31248_ (_05762_, _05761_, _05758_);
  and _31249_ (_05763_, _05762_, _05755_);
  nor _31250_ (_05764_, _05763_, _05527_);
  not _31251_ (_05765_, _02204_);
  and _31252_ (_05766_, _05527_, _05765_);
  nor _31253_ (_05767_, _05766_, _05764_);
  nor _31254_ (_05768_, _05767_, _05624_);
  not _31255_ (_05769_, _05768_);
  nor _31256_ (_05770_, _02314_, _05646_);
  not _31257_ (_05771_, _02155_);
  and _31258_ (_05772_, _05771_, _02138_);
  nor _31259_ (_05773_, _05772_, _05770_);
  and _31260_ (_05774_, _05773_, _05769_);
  and _31261_ (_05775_, _05774_, _05748_);
  nor _31262_ (_05776_, _05775_, _05603_);
  nor _31263_ (_05777_, _05723_, _00938_);
  not _31264_ (_05778_, _05777_);
  and _31265_ (_05779_, _05778_, _05776_);
  and _31266_ (_05780_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _31267_ (_05781_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _31268_ (_05782_, _05781_, _05780_);
  and _31269_ (_05783_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _31270_ (_05784_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor _31271_ (_05785_, _05784_, _05783_);
  and _31272_ (_05786_, _05785_, _05782_);
  and _31273_ (_05787_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _31274_ (_05788_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _31275_ (_05789_, _05788_, _05787_);
  and _31276_ (_05790_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _31277_ (_05791_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _31278_ (_05792_, _05791_, _05790_);
  and _31279_ (_05793_, _05792_, _05789_);
  and _31280_ (_05794_, _05793_, _05786_);
  nor _31281_ (_05795_, _05794_, _05527_);
  and _31282_ (_05796_, _05527_, _03604_);
  nor _31283_ (_05797_, _05796_, _05795_);
  nor _31284_ (_05798_, _05797_, _05624_);
  and _31285_ (_05799_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _31286_ (_05800_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not _31287_ (_05801_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _31288_ (_05802_, _01789_, _05801_);
  nor _31289_ (_05803_, _05802_, _05800_);
  and _31290_ (_05804_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _31291_ (_05805_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _31292_ (_05806_, _05805_, _05804_);
  and _31293_ (_05807_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _31294_ (_05808_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _31295_ (_05809_, _05808_, _05807_);
  and _31296_ (_05810_, _05809_, _05806_);
  and _31297_ (_05811_, _05810_, _05803_);
  nor _31298_ (_05812_, _05811_, _05577_);
  nor _31299_ (_05813_, _05812_, _05799_);
  not _31300_ (_05814_, _05813_);
  and _31301_ (_05815_, _05814_, _05605_);
  nor _31302_ (_05816_, _02320_, _02138_);
  nor _31303_ (_05817_, _05816_, _05771_);
  or _31304_ (_05818_, _05561_, _05506_);
  nor _31305_ (_05819_, _05818_, _05817_);
  or _31306_ (_05820_, _05819_, _05815_);
  nor _31307_ (_05821_, _05820_, _05798_);
  and _31308_ (_05822_, _05821_, _05604_);
  nor _31309_ (_05823_, _05723_, _02663_);
  not _31310_ (_05824_, _05823_);
  and _31311_ (_05825_, _05824_, _05822_);
  nor _31312_ (_05826_, _05825_, _05779_);
  and _31313_ (_05827_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _31314_ (_05828_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _31315_ (_05829_, _05828_, _05827_);
  and _31316_ (_05830_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _31317_ (_05831_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor _31318_ (_05832_, _05831_, _05830_);
  and _31319_ (_05833_, _05832_, _05829_);
  and _31320_ (_05834_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _31321_ (_05835_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _31322_ (_05836_, _05835_, _05834_);
  and _31323_ (_05837_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _31324_ (_05838_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _31325_ (_05839_, _05838_, _05837_);
  and _31326_ (_05840_, _05839_, _05836_);
  and _31327_ (_05841_, _05840_, _05833_);
  nor _31328_ (_05842_, _05841_, _05527_);
  and _31329_ (_05843_, _05527_, _03628_);
  nor _31330_ (_05844_, _05843_, _05842_);
  nor _31331_ (_05845_, _05844_, _05624_);
  nor _31332_ (_05846_, _05506_, _02155_);
  nor _31333_ (_05847_, _05846_, _05845_);
  nor _31334_ (_05848_, _02326_, _05646_);
  and _31335_ (_05849_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _31336_ (_05850_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not _31337_ (_05851_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _31338_ (_05852_, _01789_, _05851_);
  nor _31339_ (_05853_, _05852_, _05850_);
  and _31340_ (_05854_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _31341_ (_05855_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _31342_ (_05856_, _05855_, _05854_);
  and _31343_ (_05857_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _31344_ (_05858_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _31345_ (_05859_, _05858_, _05857_);
  and _31346_ (_05860_, _05859_, _05856_);
  and _31347_ (_05861_, _05860_, _05853_);
  nor _31348_ (_05862_, _05861_, _05577_);
  nor _31349_ (_05863_, _05862_, _05849_);
  not _31350_ (_05864_, _05863_);
  and _31351_ (_05865_, _05864_, _05605_);
  nor _31352_ (_05866_, _05865_, _05848_);
  and _31353_ (_05867_, _05866_, _05847_);
  nor _31354_ (_05868_, _05867_, _05603_);
  nor _31355_ (_05869_, _05723_, _00879_);
  not _31356_ (_05870_, _05869_);
  and _31357_ (_05871_, _05870_, _05868_);
  nor _31358_ (_05872_, _05870_, _05868_);
  nor _31359_ (_05873_, _05872_, _05871_);
  and _31360_ (_05874_, _05873_, _05826_);
  and _31361_ (_05875_, _05874_, _05729_);
  nor _31362_ (_05876_, _05821_, _05604_);
  and _31363_ (_05877_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _31364_ (_05878_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _31365_ (_05879_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _31366_ (_05880_, _05879_, _05878_);
  and _31367_ (_05881_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  not _31368_ (_05882_, _01789_);
  and _31369_ (_05883_, _05882_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _31370_ (_05884_, _05883_, _05881_);
  and _31371_ (_05885_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _31372_ (_05886_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _31373_ (_05887_, _05886_, _05885_);
  and _31374_ (_05888_, _05887_, _05884_);
  and _31375_ (_05889_, _05888_, _05880_);
  nor _31376_ (_05890_, _05889_, _05577_);
  nor _31377_ (_05891_, _05890_, _05877_);
  not _31378_ (_05892_, _05891_);
  and _31379_ (_05893_, _05892_, _05605_);
  and _31380_ (_05894_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _31381_ (_05895_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _31382_ (_05896_, _05895_, _05894_);
  and _31383_ (_05897_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _31384_ (_05898_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _31385_ (_05899_, _05898_, _05897_);
  and _31386_ (_05900_, _05899_, _05896_);
  and _31387_ (_05901_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _31388_ (_05902_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _31389_ (_05903_, _05902_, _05901_);
  and _31390_ (_05904_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _31391_ (_05905_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _31392_ (_05906_, _05905_, _05904_);
  and _31393_ (_05907_, _05906_, _05903_);
  and _31394_ (_05908_, _05907_, _05900_);
  nor _31395_ (_05909_, _05908_, _05527_);
  and _31396_ (_05910_, _05527_, _02236_);
  nor _31397_ (_05911_, _05910_, _05909_);
  nor _31398_ (_05912_, _05911_, _05624_);
  nor _31399_ (_05913_, _05912_, _05893_);
  not _31400_ (_05914_, _02302_);
  and _31401_ (_05915_, _05914_, _05645_);
  and _31402_ (_05916_, _05650_, _01924_);
  nor _31403_ (_05917_, _05916_, _05915_);
  and _31404_ (_05918_, _05917_, _05913_);
  nor _31405_ (_05919_, _05918_, _05602_);
  nor _31406_ (_05920_, _05919_, _05876_);
  and _31407_ (_05921_, _05723_, _02663_);
  nor _31408_ (_05922_, _00835_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _31409_ (_05923_, _05922_, _05921_);
  not _31410_ (_05924_, _05923_);
  and _31411_ (_05925_, _05924_, _05920_);
  nor _31412_ (_05926_, _05924_, _05920_);
  nor _31413_ (_05927_, _05926_, _05925_);
  and _31414_ (_05928_, _05723_, _02160_);
  nor _31415_ (_05929_, _05723_, _00921_);
  nor _31416_ (_05930_, _05929_, _05928_);
  and _31417_ (_05931_, _05653_, _05604_);
  and _31418_ (_05932_, _05867_, _05603_);
  nor _31419_ (_05933_, _05932_, _05931_);
  and _31420_ (_05934_, _05933_, _05930_);
  nor _31421_ (_05935_, _05933_, _05930_);
  or _31422_ (_05936_, _05935_, _05934_);
  not _31423_ (_05937_, _05936_);
  and _31424_ (_05938_, _05937_, _05927_);
  or _31425_ (_05939_, _05775_, _05604_);
  and _31426_ (_05940_, _05650_, _01902_);
  and _31427_ (_05941_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _31428_ (_05942_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _31429_ (_05943_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _31430_ (_05944_, _05943_, _05942_);
  and _31431_ (_05945_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not _31432_ (_05946_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _31433_ (_05947_, _01789_, _05946_);
  nor _31434_ (_05948_, _05947_, _05945_);
  and _31435_ (_05949_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _31436_ (_05950_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _31437_ (_05962_, _05950_, _05949_);
  and _31438_ (_05963_, _05962_, _05948_);
  and _31439_ (_05964_, _05963_, _05944_);
  nor _31440_ (_05965_, _05964_, _05577_);
  nor _31441_ (_05966_, _05965_, _05941_);
  not _31442_ (_05967_, _05966_);
  and _31443_ (_05968_, _05967_, _05605_);
  nor _31444_ (_05969_, _05968_, _05940_);
  and _31445_ (_05970_, _05546_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _31446_ (_05971_, _05544_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _31447_ (_05972_, _05971_, _05970_);
  and _31448_ (_05973_, _05530_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _31449_ (_05974_, _05551_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _31450_ (_05975_, _05974_, _05973_);
  and _31451_ (_05976_, _05975_, _05972_);
  and _31452_ (_05977_, _05539_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _31453_ (_05978_, _05533_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _31454_ (_05979_, _05978_, _05977_);
  and _31455_ (_05980_, _05549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _31456_ (_05981_, _05537_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _31457_ (_05982_, _05981_, _05980_);
  and _31458_ (_05983_, _05982_, _05979_);
  and _31459_ (_05984_, _05983_, _05976_);
  nor _31460_ (_05985_, _05984_, _05527_);
  and _31461_ (_05986_, _05527_, _02251_);
  nor _31462_ (_05987_, _05986_, _05985_);
  nor _31463_ (_05988_, _05987_, _05624_);
  not _31464_ (_05989_, _05988_);
  and _31465_ (_05990_, _05506_, _05771_);
  nor _31466_ (_05991_, _02296_, _05646_);
  nor _31467_ (_05992_, _05991_, _05990_);
  and _31468_ (_05993_, _05992_, _05989_);
  and _31469_ (_05994_, _05993_, _05969_);
  or _31470_ (_05995_, _05994_, _05602_);
  and _31471_ (_05996_, _05995_, _05939_);
  not _31472_ (_05997_, _05996_);
  and _31473_ (_05998_, _05723_, _03985_);
  nor _31474_ (_05999_, _00847_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _31475_ (_06000_, _05999_, _05998_);
  nor _31476_ (_06001_, _06000_, _05997_);
  and _31477_ (_06002_, _06000_, _05997_);
  nor _31478_ (_06003_, _06002_, _06001_);
  nor _31479_ (_06004_, _05824_, _05822_);
  not _31480_ (_06005_, _06004_);
  nor _31481_ (_06006_, _05778_, _05776_);
  nor _31482_ (_06007_, _00906_, _00812_);
  nor _31483_ (_06008_, _06007_, _01188_);
  not _31484_ (_06009_, _06008_);
  nor _31485_ (_06010_, _05584_, _00906_);
  and _31486_ (_06011_, _05584_, _00906_);
  nor _31487_ (_06012_, _06011_, _06010_);
  nor _31488_ (_06013_, _06012_, _06009_);
  not _31489_ (_06014_, _06013_);
  nor _31490_ (_06015_, _06014_, _06006_);
  and _31491_ (_06016_, _06015_, _06005_);
  and _31492_ (_06017_, _06016_, _06003_);
  and _31493_ (_06018_, _06017_, _05938_);
  and _31494_ (_06019_, _06018_, _05875_);
  not _31495_ (_06020_, _05584_);
  not _31496_ (_06021_, _05920_);
  and _31497_ (_06022_, _05721_, _05654_);
  and _31498_ (_06023_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and _31499_ (_06024_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _31500_ (_06025_, _06024_, _06023_);
  and _31501_ (_06026_, _06025_, _05997_);
  and _31502_ (_06027_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and _31503_ (_06028_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _31504_ (_06029_, _06028_, _06027_);
  and _31505_ (_06030_, _06029_, _05996_);
  or _31506_ (_06031_, _06030_, _06026_);
  or _31507_ (_06032_, _06031_, _06021_);
  not _31508_ (_06033_, _05933_);
  and _31509_ (_06034_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and _31510_ (_06035_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _31511_ (_06036_, _06035_, _06034_);
  and _31512_ (_06037_, _06036_, _05997_);
  and _31513_ (_06038_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and _31514_ (_06039_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _31515_ (_06040_, _06039_, _06038_);
  and _31516_ (_06041_, _06040_, _05996_);
  or _31517_ (_06042_, _06041_, _06037_);
  or _31518_ (_06043_, _06042_, _05920_);
  and _31519_ (_06044_, _06043_, _06033_);
  and _31520_ (_06045_, _06044_, _06032_);
  or _31521_ (_06046_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _31522_ (_06047_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and _31523_ (_06048_, _06047_, _05996_);
  and _31524_ (_06049_, _06048_, _06046_);
  or _31525_ (_06050_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _31526_ (_06051_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and _31527_ (_06052_, _06051_, _05997_);
  and _31528_ (_06053_, _06052_, _06050_);
  or _31529_ (_06054_, _06053_, _06049_);
  or _31530_ (_06055_, _06054_, _06021_);
  or _31531_ (_06056_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _31532_ (_06057_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and _31533_ (_06058_, _06057_, _05996_);
  and _31534_ (_06059_, _06058_, _06056_);
  or _31535_ (_06060_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _31536_ (_06061_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and _31537_ (_06062_, _06061_, _05997_);
  and _31538_ (_06063_, _06062_, _06060_);
  or _31539_ (_06064_, _06063_, _06059_);
  or _31540_ (_06065_, _06064_, _05920_);
  and _31541_ (_06066_, _06065_, _05933_);
  and _31542_ (_06067_, _06066_, _06055_);
  or _31543_ (_06068_, _06067_, _06045_);
  or _31544_ (_06069_, _06068_, _05776_);
  not _31545_ (_06070_, _05822_);
  not _31546_ (_06071_, _05776_);
  and _31547_ (_06072_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and _31548_ (_06073_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _31549_ (_06074_, _06073_, _05996_);
  or _31550_ (_06075_, _06074_, _06072_);
  and _31551_ (_06076_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _31552_ (_06077_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _31553_ (_06078_, _06077_, _05997_);
  or _31554_ (_06082_, _06078_, _06076_);
  and _31555_ (_06095_, _06082_, _06075_);
  or _31556_ (_06105_, _06095_, _06021_);
  and _31557_ (_06106_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and _31558_ (_06109_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _31559_ (_06110_, _06109_, _05996_);
  or _31560_ (_06111_, _06110_, _06106_);
  and _31561_ (_06112_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and _31562_ (_06133_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _31563_ (_06147_, _06133_, _05997_);
  or _31564_ (_06148_, _06147_, _06112_);
  and _31565_ (_06149_, _06148_, _06111_);
  or _31566_ (_06153_, _06149_, _05920_);
  and _31567_ (_06181_, _06153_, _06033_);
  and _31568_ (_06182_, _06181_, _06105_);
  or _31569_ (_06183_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _31570_ (_06184_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and _31571_ (_06185_, _06184_, _06183_);
  or _31572_ (_06186_, _06185_, _05997_);
  or _31573_ (_06187_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _31574_ (_06188_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and _31575_ (_06189_, _06188_, _06187_);
  or _31576_ (_06190_, _06189_, _05996_);
  and _31577_ (_06191_, _06190_, _06186_);
  or _31578_ (_06192_, _06191_, _06021_);
  or _31579_ (_06193_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _31580_ (_06194_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and _31581_ (_06195_, _06194_, _06193_);
  or _31582_ (_06196_, _06195_, _05997_);
  or _31583_ (_06197_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _31584_ (_06198_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and _31585_ (_06199_, _06198_, _06197_);
  or _31586_ (_06257_, _06199_, _05996_);
  and _31587_ (_06358_, _06257_, _06196_);
  or _31588_ (_06396_, _06358_, _05920_);
  and _31589_ (_06397_, _06396_, _05933_);
  and _31590_ (_06398_, _06397_, _06192_);
  or _31591_ (_06399_, _06398_, _06182_);
  or _31592_ (_06400_, _06399_, _06071_);
  and _31593_ (_06401_, _06400_, _06070_);
  and _31594_ (_06402_, _06401_, _06069_);
  and _31595_ (_06403_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _31596_ (_06404_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _31597_ (_06405_, _06404_, _06403_);
  and _31598_ (_06406_, _06405_, _05996_);
  and _31599_ (_06407_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and _31600_ (_06408_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _31601_ (_06409_, _06408_, _06407_);
  and _31602_ (_06410_, _06409_, _05997_);
  or _31603_ (_06411_, _06410_, _06406_);
  and _31604_ (_06412_, _06411_, _05920_);
  and _31605_ (_06413_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and _31606_ (_06414_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _31607_ (_06415_, _06414_, _06413_);
  and _31608_ (_06416_, _06415_, _05996_);
  and _31609_ (_06417_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and _31610_ (_06418_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _31611_ (_06428_, _06418_, _06417_);
  and _31612_ (_06429_, _06428_, _05997_);
  or _31613_ (_06430_, _06429_, _06416_);
  and _31614_ (_06431_, _06430_, _06021_);
  or _31615_ (_06432_, _06431_, _06412_);
  and _31616_ (_06433_, _06432_, _06033_);
  or _31617_ (_06434_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _31618_ (_06435_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _31619_ (_06436_, _06435_, _06434_);
  and _31620_ (_06437_, _06436_, _05996_);
  or _31621_ (_06485_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _31622_ (_06495_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and _31623_ (_06496_, _06495_, _06485_);
  and _31624_ (_06497_, _06496_, _05997_);
  or _31625_ (_06498_, _06497_, _06437_);
  and _31626_ (_06499_, _06498_, _05920_);
  or _31627_ (_06500_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _31628_ (_06507_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _31629_ (_06508_, _06507_, _06500_);
  and _31630_ (_06509_, _06508_, _05996_);
  or _31631_ (_06510_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _31632_ (_06511_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _31633_ (_06512_, _06511_, _06510_);
  and _31634_ (_06513_, _06512_, _05997_);
  or _31635_ (_06514_, _06513_, _06509_);
  and _31636_ (_06525_, _06514_, _06021_);
  or _31637_ (_06526_, _06525_, _06499_);
  and _31638_ (_06527_, _06526_, _05933_);
  or _31639_ (_06528_, _06527_, _06433_);
  and _31640_ (_06529_, _06528_, _06071_);
  and _31641_ (_06530_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and _31642_ (_06531_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _31643_ (_06532_, _06531_, _06530_);
  and _31644_ (_06537_, _06532_, _05996_);
  and _31645_ (_06547_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and _31646_ (_06548_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _31647_ (_06549_, _06548_, _06547_);
  and _31648_ (_06550_, _06549_, _05997_);
  or _31649_ (_06551_, _06550_, _06537_);
  and _31650_ (_06552_, _06551_, _05920_);
  and _31651_ (_06553_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and _31652_ (_06554_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _31653_ (_06555_, _06554_, _06553_);
  and _31654_ (_06556_, _06555_, _05996_);
  and _31655_ (_06557_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and _31656_ (_06558_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _31657_ (_06559_, _06558_, _06557_);
  and _31658_ (_06560_, _06559_, _05997_);
  or _31659_ (_06561_, _06560_, _06556_);
  and _31660_ (_06562_, _06561_, _06021_);
  or _31661_ (_06563_, _06562_, _06552_);
  and _31662_ (_06564_, _06563_, _06033_);
  or _31663_ (_06565_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _31664_ (_06566_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and _31665_ (_06567_, _06566_, _06565_);
  and _31666_ (_06568_, _06567_, _05996_);
  or _31667_ (_06569_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _31668_ (_06570_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and _31669_ (_06571_, _06570_, _06569_);
  and _31670_ (_06572_, _06571_, _05997_);
  or _31671_ (_06573_, _06572_, _06568_);
  and _31672_ (_06574_, _06573_, _05920_);
  or _31673_ (_06575_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _31674_ (_06576_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and _31675_ (_06577_, _06576_, _06575_);
  and _31676_ (_06578_, _06577_, _05996_);
  or _31677_ (_06579_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _31678_ (_06580_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and _31679_ (_06581_, _06580_, _06579_);
  and _31680_ (_06582_, _06581_, _05997_);
  or _31681_ (_06589_, _06582_, _06578_);
  and _31682_ (_06607_, _06589_, _06021_);
  or _31683_ (_06608_, _06607_, _06574_);
  and _31684_ (_06609_, _06608_, _05933_);
  or _31685_ (_06610_, _06609_, _06564_);
  and _31686_ (_06611_, _06610_, _05776_);
  or _31687_ (_06612_, _06611_, _06529_);
  and _31688_ (_06613_, _06612_, _05822_);
  or _31689_ (_06614_, _06613_, _06402_);
  or _31690_ (_06615_, _06614_, _05868_);
  not _31691_ (_06616_, _05868_);
  and _31692_ (_06617_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and _31693_ (_06618_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _31694_ (_06619_, _06618_, _06617_);
  and _31695_ (_06620_, _06619_, _05996_);
  and _31696_ (_06621_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and _31697_ (_06622_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _31698_ (_06623_, _06622_, _06621_);
  and _31699_ (_06624_, _06623_, _05997_);
  or _31700_ (_06625_, _06624_, _06620_);
  or _31701_ (_06626_, _06625_, _06021_);
  and _31702_ (_06627_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and _31703_ (_06628_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _31704_ (_06629_, _06628_, _06627_);
  and _31705_ (_06630_, _06629_, _05996_);
  and _31706_ (_06631_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and _31707_ (_06632_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _31708_ (_06633_, _06632_, _06631_);
  and _31709_ (_06634_, _06633_, _05997_);
  or _31710_ (_06635_, _06634_, _06630_);
  or _31711_ (_06636_, _06635_, _05920_);
  and _31712_ (_06637_, _06636_, _06033_);
  and _31713_ (_06638_, _06637_, _06626_);
  or _31714_ (_06639_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _31715_ (_06640_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and _31716_ (_06641_, _06640_, _05997_);
  and _31717_ (_06642_, _06641_, _06639_);
  or _31718_ (_06643_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _31719_ (_06644_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and _31720_ (_06645_, _06644_, _05996_);
  and _31721_ (_06646_, _06645_, _06643_);
  or _31722_ (_06647_, _06646_, _06642_);
  or _31723_ (_06648_, _06647_, _06021_);
  or _31724_ (_06649_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _31725_ (_06650_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and _31726_ (_06651_, _06650_, _05997_);
  and _31727_ (_06652_, _06651_, _06649_);
  or _31728_ (_06653_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _31729_ (_06654_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and _31730_ (_06655_, _06654_, _05996_);
  and _31731_ (_06656_, _06655_, _06653_);
  or _31732_ (_06657_, _06656_, _06652_);
  or _31733_ (_06658_, _06657_, _05920_);
  and _31734_ (_06659_, _06658_, _05933_);
  and _31735_ (_06660_, _06659_, _06648_);
  or _31736_ (_06661_, _06660_, _06638_);
  and _31737_ (_06662_, _06661_, _06071_);
  and _31738_ (_06663_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and _31739_ (_06664_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _31740_ (_06665_, _06664_, _06663_);
  and _31741_ (_06666_, _06665_, _05996_);
  and _31742_ (_06667_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and _31743_ (_06668_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _31744_ (_06669_, _06668_, _06667_);
  and _31745_ (_06670_, _06669_, _05997_);
  or _31746_ (_06671_, _06670_, _06666_);
  or _31747_ (_06672_, _06671_, _06021_);
  and _31748_ (_06673_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and _31749_ (_06674_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _31750_ (_06675_, _06674_, _06673_);
  and _31751_ (_06676_, _06675_, _05996_);
  and _31752_ (_06677_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and _31753_ (_06678_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _31754_ (_06679_, _06678_, _06677_);
  and _31755_ (_06680_, _06679_, _05997_);
  or _31756_ (_06681_, _06680_, _06676_);
  or _31757_ (_06682_, _06681_, _05920_);
  and _31758_ (_06683_, _06682_, _06033_);
  and _31759_ (_06684_, _06683_, _06672_);
  or _31760_ (_06685_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _31761_ (_06686_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and _31762_ (_06687_, _06686_, _06685_);
  and _31763_ (_06688_, _06687_, _05996_);
  or _31764_ (_06689_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _31765_ (_06690_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _31766_ (_06691_, _06690_, _06689_);
  and _31767_ (_06692_, _06691_, _05997_);
  or _31768_ (_06693_, _06692_, _06688_);
  or _31769_ (_06694_, _06693_, _06021_);
  or _31770_ (_06695_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _31771_ (_06696_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and _31772_ (_06697_, _06696_, _06695_);
  and _31773_ (_06698_, _06697_, _05996_);
  or _31774_ (_06699_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _31775_ (_06700_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and _31776_ (_06701_, _06700_, _06699_);
  and _31777_ (_06702_, _06701_, _05997_);
  or _31778_ (_06703_, _06702_, _06698_);
  or _31779_ (_06704_, _06703_, _05920_);
  and _31780_ (_06705_, _06704_, _05933_);
  and _31781_ (_06706_, _06705_, _06694_);
  or _31782_ (_06707_, _06706_, _06684_);
  and _31783_ (_06708_, _06707_, _05776_);
  or _31784_ (_06709_, _06708_, _06662_);
  and _31785_ (_06716_, _06709_, _06070_);
  or _31786_ (_06718_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _31787_ (_06720_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and _31788_ (_06721_, _06720_, _06718_);
  and _31789_ (_06722_, _06721_, _05996_);
  or _31790_ (_06723_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _31791_ (_06724_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and _31792_ (_06725_, _06724_, _06723_);
  and _31793_ (_06745_, _06725_, _05997_);
  or _31794_ (_06777_, _06745_, _06722_);
  and _31795_ (_06809_, _06777_, _06021_);
  or _31796_ (_06842_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _31797_ (_06874_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and _31798_ (_06909_, _06874_, _06842_);
  and _31799_ (_06943_, _06909_, _05996_);
  or _31800_ (_06977_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _31801_ (_07010_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and _31802_ (_07045_, _07010_, _06977_);
  and _31803_ (_07079_, _07045_, _05997_);
  or _31804_ (_07113_, _07079_, _06943_);
  and _31805_ (_07147_, _07113_, _05920_);
  or _31806_ (_07181_, _07147_, _06809_);
  and _31807_ (_07216_, _07181_, _05933_);
  and _31808_ (_07250_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and _31809_ (_07283_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _31810_ (_07317_, _07283_, _07250_);
  and _31811_ (_07352_, _07317_, _05996_);
  and _31812_ (_07386_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and _31813_ (_07420_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _31814_ (_07454_, _07420_, _07386_);
  and _31815_ (_07489_, _07454_, _05997_);
  or _31816_ (_07523_, _07489_, _07352_);
  and _31817_ (_07557_, _07523_, _06021_);
  and _31818_ (_07591_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and _31819_ (_07626_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _31820_ (_07660_, _07626_, _07591_);
  and _31821_ (_07694_, _07660_, _05996_);
  and _31822_ (_07728_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and _31823_ (_07763_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _31824_ (_07796_, _07763_, _07728_);
  and _31825_ (_07830_, _07796_, _05997_);
  or _31826_ (_07864_, _07830_, _07694_);
  and _31827_ (_07899_, _07864_, _05920_);
  or _31828_ (_07933_, _07899_, _07557_);
  and _31829_ (_07967_, _07933_, _06033_);
  or _31830_ (_08001_, _07967_, _07216_);
  and _31831_ (_08036_, _08001_, _05776_);
  or _31832_ (_08070_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _31833_ (_08104_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and _31834_ (_08138_, _08104_, _05997_);
  and _31835_ (_08173_, _08138_, _08070_);
  or _31836_ (_08207_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or _31837_ (_08241_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and _31838_ (_08275_, _08241_, _05996_);
  and _31839_ (_08309_, _08275_, _08207_);
  or _31840_ (_08343_, _08309_, _08173_);
  and _31841_ (_08378_, _08343_, _06021_);
  or _31842_ (_08412_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _31843_ (_08446_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and _31844_ (_08481_, _08446_, _05997_);
  and _31845_ (_08515_, _08481_, _08412_);
  or _31846_ (_08549_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or _31847_ (_08583_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and _31848_ (_08617_, _08583_, _05996_);
  and _31849_ (_08652_, _08617_, _08549_);
  or _31850_ (_08686_, _08652_, _08515_);
  and _31851_ (_08720_, _08686_, _05920_);
  or _31852_ (_08754_, _08720_, _08378_);
  and _31853_ (_08789_, _08754_, _05933_);
  and _31854_ (_08823_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and _31855_ (_08835_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _31856_ (_08836_, _08835_, _08823_);
  and _31857_ (_08837_, _08836_, _05996_);
  and _31858_ (_08838_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and _31859_ (_08839_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _31860_ (_08840_, _08839_, _08838_);
  and _31861_ (_08841_, _08840_, _05997_);
  or _31862_ (_08842_, _08841_, _08837_);
  and _31863_ (_08843_, _08842_, _06021_);
  and _31864_ (_08844_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and _31865_ (_08845_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or _31866_ (_08846_, _08845_, _08844_);
  and _31867_ (_08847_, _08846_, _05996_);
  and _31868_ (_08848_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and _31869_ (_08849_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _31870_ (_08850_, _08849_, _08848_);
  and _31871_ (_08851_, _08850_, _05997_);
  or _31872_ (_08852_, _08851_, _08847_);
  and _31873_ (_08853_, _08852_, _05920_);
  or _31874_ (_08854_, _08853_, _08843_);
  and _31875_ (_08855_, _08854_, _06033_);
  or _31876_ (_08856_, _08855_, _08789_);
  and _31877_ (_08857_, _08856_, _06071_);
  or _31878_ (_08858_, _08857_, _08036_);
  and _31879_ (_08859_, _08858_, _05822_);
  or _31880_ (_08860_, _08859_, _06716_);
  or _31881_ (_08861_, _08860_, _06616_);
  and _31882_ (_08862_, _08861_, _06615_);
  or _31883_ (_08863_, _08862_, _06020_);
  and _31884_ (_08864_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and _31885_ (_08865_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _31886_ (_08866_, _08865_, _08864_);
  and _31887_ (_08867_, _08866_, _05996_);
  and _31888_ (_08868_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and _31889_ (_08869_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _31890_ (_08870_, _08869_, _08868_);
  and _31891_ (_08871_, _08870_, _05997_);
  or _31892_ (_08872_, _08871_, _08867_);
  or _31893_ (_08873_, _08872_, _06021_);
  and _31894_ (_08874_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and _31895_ (_08875_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _31896_ (_08876_, _08875_, _08874_);
  and _31897_ (_08877_, _08876_, _05996_);
  and _31898_ (_08878_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and _31899_ (_08879_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _31900_ (_08880_, _08879_, _08878_);
  and _31901_ (_08881_, _08880_, _05997_);
  or _31902_ (_08882_, _08881_, _08877_);
  or _31903_ (_08883_, _08882_, _05920_);
  and _31904_ (_08884_, _08883_, _06033_);
  and _31905_ (_08885_, _08884_, _08873_);
  or _31906_ (_08886_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _31907_ (_08887_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and _31908_ (_08888_, _08887_, _08886_);
  and _31909_ (_08889_, _08888_, _05996_);
  or _31910_ (_08890_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _31911_ (_08891_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and _31912_ (_08892_, _08891_, _08890_);
  and _31913_ (_08894_, _08892_, _05997_);
  or _31914_ (_08895_, _08894_, _08889_);
  or _31915_ (_08896_, _08895_, _06021_);
  or _31916_ (_08897_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _31917_ (_08898_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and _31918_ (_08899_, _08898_, _08897_);
  and _31919_ (_08900_, _08899_, _05996_);
  or _31920_ (_08901_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _31921_ (_08902_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and _31922_ (_08903_, _08902_, _08901_);
  and _31923_ (_08904_, _08903_, _05997_);
  or _31924_ (_08905_, _08904_, _08900_);
  or _31925_ (_08906_, _08905_, _05920_);
  and _31926_ (_08907_, _08906_, _05933_);
  and _31927_ (_08908_, _08907_, _08896_);
  or _31928_ (_08909_, _08908_, _08885_);
  and _31929_ (_08910_, _08909_, _05776_);
  and _31930_ (_08911_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _31931_ (_08912_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _31932_ (_08913_, _08912_, _08911_);
  and _31933_ (_08914_, _08913_, _05996_);
  and _31934_ (_08915_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _31935_ (_08916_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _31936_ (_08917_, _08916_, _08915_);
  and _31937_ (_08918_, _08917_, _05997_);
  or _31938_ (_08919_, _08918_, _08914_);
  or _31939_ (_08920_, _08919_, _06021_);
  and _31940_ (_08921_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _31941_ (_08922_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _31942_ (_08923_, _08922_, _08921_);
  and _31943_ (_08924_, _08923_, _05996_);
  and _31944_ (_08925_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _31945_ (_08926_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _31946_ (_08927_, _08926_, _08925_);
  and _31947_ (_08928_, _08927_, _05997_);
  or _31948_ (_08929_, _08928_, _08924_);
  or _31949_ (_08930_, _08929_, _05920_);
  and _31950_ (_08931_, _08930_, _06033_);
  and _31951_ (_08932_, _08931_, _08920_);
  or _31952_ (_08933_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _31953_ (_08934_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _31954_ (_08935_, _08934_, _05997_);
  and _31955_ (_08936_, _08935_, _08933_);
  or _31956_ (_08937_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or _31957_ (_08938_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _31958_ (_08939_, _08938_, _05996_);
  and _31959_ (_08940_, _08939_, _08937_);
  or _31960_ (_08941_, _08940_, _08936_);
  or _31961_ (_08942_, _08941_, _06021_);
  or _31962_ (_08943_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or _31963_ (_08944_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _31964_ (_08945_, _08944_, _05997_);
  and _31965_ (_08946_, _08945_, _08943_);
  or _31966_ (_08947_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _31967_ (_08948_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and _31968_ (_08949_, _08948_, _05996_);
  and _31969_ (_08950_, _08949_, _08947_);
  or _31970_ (_08951_, _08950_, _08946_);
  or _31971_ (_08952_, _08951_, _05920_);
  and _31972_ (_08953_, _08952_, _05933_);
  and _31973_ (_08954_, _08953_, _08942_);
  or _31974_ (_08955_, _08954_, _08932_);
  and _31975_ (_08956_, _08955_, _06071_);
  or _31976_ (_08957_, _08956_, _08910_);
  and _31977_ (_08958_, _08957_, _06070_);
  and _31978_ (_08959_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and _31979_ (_08960_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _31980_ (_08961_, _08960_, _08959_);
  and _31981_ (_08962_, _08961_, _05996_);
  and _31982_ (_08963_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and _31983_ (_08964_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _31984_ (_08965_, _08964_, _08963_);
  and _31985_ (_08966_, _08965_, _05997_);
  or _31986_ (_08967_, _08966_, _08962_);
  and _31987_ (_08968_, _08967_, _05920_);
  and _31988_ (_08969_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and _31989_ (_08970_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or _31990_ (_08971_, _08970_, _08969_);
  and _31991_ (_08972_, _08971_, _05996_);
  and _31992_ (_08973_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and _31993_ (_08974_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or _31994_ (_08975_, _08974_, _08973_);
  and _31995_ (_08976_, _08975_, _05997_);
  or _31996_ (_08977_, _08976_, _08972_);
  and _31997_ (_08978_, _08977_, _06021_);
  or _31998_ (_08979_, _08978_, _08968_);
  and _31999_ (_08980_, _08979_, _06033_);
  or _32000_ (_08981_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or _32001_ (_08982_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _32002_ (_08983_, _08982_, _05997_);
  and _32003_ (_08984_, _08983_, _08981_);
  or _32004_ (_08985_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or _32005_ (_08986_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and _32006_ (_08987_, _08986_, _05996_);
  and _32007_ (_08988_, _08987_, _08985_);
  or _32008_ (_08989_, _08988_, _08984_);
  and _32009_ (_08990_, _08989_, _05920_);
  or _32010_ (_08991_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or _32011_ (_08992_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and _32012_ (_08993_, _08992_, _05997_);
  and _32013_ (_08994_, _08993_, _08991_);
  or _32014_ (_08995_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or _32015_ (_08996_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and _32016_ (_08997_, _08996_, _05996_);
  and _32017_ (_08998_, _08997_, _08995_);
  or _32018_ (_08999_, _08998_, _08994_);
  and _32019_ (_09000_, _08999_, _06021_);
  or _32020_ (_09001_, _09000_, _08990_);
  and _32021_ (_09002_, _09001_, _05933_);
  or _32022_ (_09003_, _09002_, _08980_);
  and _32023_ (_09004_, _09003_, _06071_);
  and _32024_ (_09005_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and _32025_ (_09006_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _32026_ (_09007_, _09006_, _09005_);
  and _32027_ (_09008_, _09007_, _05996_);
  and _32028_ (_09009_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _32029_ (_09010_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _32030_ (_09011_, _09010_, _09009_);
  and _32031_ (_09012_, _09011_, _05997_);
  or _32032_ (_09013_, _09012_, _09008_);
  and _32033_ (_09014_, _09013_, _05920_);
  and _32034_ (_09015_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and _32035_ (_09016_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _32036_ (_09017_, _09016_, _09015_);
  and _32037_ (_09018_, _09017_, _05996_);
  and _32038_ (_09019_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and _32039_ (_09020_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _32040_ (_09021_, _09020_, _09019_);
  and _32041_ (_09022_, _09021_, _05997_);
  or _32042_ (_09023_, _09022_, _09018_);
  and _32043_ (_09024_, _09023_, _06021_);
  or _32044_ (_09025_, _09024_, _09014_);
  and _32045_ (_09026_, _09025_, _06033_);
  or _32046_ (_09027_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _32047_ (_09028_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and _32048_ (_09029_, _09028_, _09027_);
  and _32049_ (_09030_, _09029_, _05996_);
  or _32050_ (_09031_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _32051_ (_09032_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _32052_ (_09033_, _09032_, _09031_);
  and _32053_ (_09034_, _09033_, _05997_);
  or _32054_ (_09035_, _09034_, _09030_);
  and _32055_ (_09036_, _09035_, _05920_);
  or _32056_ (_09037_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _32057_ (_09038_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _32058_ (_09039_, _09038_, _09037_);
  and _32059_ (_09040_, _09039_, _05996_);
  or _32060_ (_09041_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _32061_ (_09042_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and _32062_ (_09043_, _09042_, _09041_);
  and _32063_ (_09044_, _09043_, _05997_);
  or _32064_ (_09045_, _09044_, _09040_);
  and _32065_ (_09046_, _09045_, _06021_);
  or _32066_ (_09047_, _09046_, _09036_);
  and _32067_ (_09048_, _09047_, _05933_);
  or _32068_ (_09049_, _09048_, _09026_);
  and _32069_ (_09050_, _09049_, _05776_);
  or _32070_ (_09051_, _09050_, _09004_);
  and _32071_ (_09052_, _09051_, _05822_);
  or _32072_ (_09053_, _09052_, _08958_);
  or _32073_ (_09054_, _09053_, _05868_);
  and _32074_ (_09055_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and _32075_ (_09056_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _32076_ (_09057_, _09056_, _09055_);
  and _32077_ (_09058_, _09057_, _05996_);
  and _32078_ (_09059_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and _32079_ (_09060_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _32080_ (_09061_, _09060_, _09059_);
  and _32081_ (_09062_, _09061_, _05997_);
  or _32082_ (_09063_, _09062_, _09058_);
  or _32083_ (_09064_, _09063_, _06021_);
  and _32084_ (_09065_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and _32085_ (_09066_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _32086_ (_09067_, _09066_, _09065_);
  and _32087_ (_09068_, _09067_, _05996_);
  and _32088_ (_09069_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and _32089_ (_09070_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _32090_ (_09071_, _09070_, _09069_);
  and _32091_ (_09072_, _09071_, _05997_);
  or _32092_ (_09073_, _09072_, _09068_);
  or _32093_ (_09074_, _09073_, _05920_);
  and _32094_ (_09075_, _09074_, _06033_);
  and _32095_ (_09076_, _09075_, _09064_);
  or _32096_ (_09077_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _32097_ (_09078_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and _32098_ (_09079_, _09078_, _05997_);
  and _32099_ (_09080_, _09079_, _09077_);
  or _32100_ (_09081_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _32101_ (_09082_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and _32102_ (_09083_, _09082_, _05996_);
  and _32103_ (_09084_, _09083_, _09081_);
  or _32104_ (_09085_, _09084_, _09080_);
  or _32105_ (_09086_, _09085_, _06021_);
  or _32106_ (_09087_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _32107_ (_09088_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and _32108_ (_09089_, _09088_, _05997_);
  and _32109_ (_09090_, _09089_, _09087_);
  or _32110_ (_09091_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _32111_ (_09092_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and _32112_ (_09093_, _09092_, _05996_);
  and _32113_ (_09094_, _09093_, _09091_);
  or _32114_ (_09095_, _09094_, _09090_);
  or _32115_ (_09096_, _09095_, _05920_);
  and _32116_ (_09097_, _09096_, _05933_);
  and _32117_ (_09098_, _09097_, _09086_);
  or _32118_ (_09099_, _09098_, _09076_);
  and _32119_ (_09100_, _09099_, _06071_);
  and _32120_ (_09101_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and _32121_ (_09102_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _32122_ (_09103_, _09102_, _09101_);
  and _32123_ (_09104_, _09103_, _05996_);
  and _32124_ (_09105_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _32125_ (_09106_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or _32126_ (_09107_, _09106_, _09105_);
  and _32127_ (_09108_, _09107_, _05997_);
  or _32128_ (_09109_, _09108_, _09104_);
  or _32129_ (_09110_, _09109_, _06021_);
  and _32130_ (_09111_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and _32131_ (_09112_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or _32132_ (_09113_, _09112_, _09111_);
  and _32133_ (_09114_, _09113_, _05996_);
  and _32134_ (_09115_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and _32135_ (_09116_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _32136_ (_09117_, _09116_, _09115_);
  and _32137_ (_09118_, _09117_, _05997_);
  or _32138_ (_09119_, _09118_, _09114_);
  or _32139_ (_09120_, _09119_, _05920_);
  and _32140_ (_09121_, _09120_, _06033_);
  and _32141_ (_09122_, _09121_, _09110_);
  or _32142_ (_09123_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _32143_ (_09124_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _32144_ (_09125_, _09124_, _09123_);
  and _32145_ (_09126_, _09125_, _05996_);
  or _32146_ (_09127_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _32147_ (_09128_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and _32148_ (_09129_, _09128_, _09127_);
  and _32149_ (_09130_, _09129_, _05997_);
  or _32150_ (_09131_, _09130_, _09126_);
  or _32151_ (_09132_, _09131_, _06021_);
  or _32152_ (_09133_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _32153_ (_09134_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _32154_ (_09135_, _09134_, _09133_);
  and _32155_ (_09136_, _09135_, _05996_);
  or _32156_ (_09137_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _32157_ (_09138_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _32158_ (_09139_, _09138_, _09137_);
  and _32159_ (_09140_, _09139_, _05997_);
  or _32160_ (_09141_, _09140_, _09136_);
  or _32161_ (_09142_, _09141_, _05920_);
  and _32162_ (_09143_, _09142_, _05933_);
  and _32163_ (_09144_, _09143_, _09132_);
  or _32164_ (_09145_, _09144_, _09122_);
  and _32165_ (_09146_, _09145_, _05776_);
  or _32166_ (_09147_, _09146_, _09100_);
  and _32167_ (_09148_, _09147_, _06070_);
  or _32168_ (_09149_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _32169_ (_09150_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _32170_ (_09151_, _09150_, _09149_);
  and _32171_ (_09152_, _09151_, _05996_);
  or _32172_ (_09153_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _32173_ (_09154_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and _32174_ (_09155_, _09154_, _09153_);
  and _32175_ (_09156_, _09155_, _05997_);
  or _32176_ (_09157_, _09156_, _09152_);
  and _32177_ (_09158_, _09157_, _06021_);
  or _32178_ (_09159_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _32179_ (_09160_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _32180_ (_09161_, _09160_, _09159_);
  and _32181_ (_09162_, _09161_, _05996_);
  or _32182_ (_09163_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or _32183_ (_09164_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _32184_ (_09165_, _09164_, _09163_);
  and _32185_ (_09166_, _09165_, _05997_);
  or _32186_ (_09167_, _09166_, _09162_);
  and _32187_ (_09168_, _09167_, _05920_);
  or _32188_ (_09169_, _09168_, _09158_);
  and _32189_ (_09170_, _09169_, _05933_);
  and _32190_ (_09171_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and _32191_ (_09172_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _32192_ (_09173_, _09172_, _09171_);
  and _32193_ (_09174_, _09173_, _05996_);
  and _32194_ (_09175_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _32195_ (_09176_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _32196_ (_09177_, _09176_, _09175_);
  and _32197_ (_09178_, _09177_, _05997_);
  or _32198_ (_09179_, _09178_, _09174_);
  and _32199_ (_09180_, _09179_, _06021_);
  and _32200_ (_09181_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _32201_ (_09182_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _32202_ (_09183_, _09182_, _09181_);
  and _32203_ (_09184_, _09183_, _05996_);
  and _32204_ (_09185_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _32205_ (_09186_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _32206_ (_09187_, _09186_, _09185_);
  and _32207_ (_09188_, _09187_, _05997_);
  or _32208_ (_09189_, _09188_, _09184_);
  and _32209_ (_09190_, _09189_, _05920_);
  or _32210_ (_09191_, _09190_, _09180_);
  and _32211_ (_09192_, _09191_, _06033_);
  or _32212_ (_09193_, _09192_, _09170_);
  and _32213_ (_09194_, _09193_, _05776_);
  or _32214_ (_09195_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or _32215_ (_09196_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and _32216_ (_09197_, _09196_, _05997_);
  and _32217_ (_09198_, _09197_, _09195_);
  or _32218_ (_09199_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _32219_ (_09200_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and _32220_ (_09201_, _09200_, _05996_);
  and _32221_ (_09202_, _09201_, _09199_);
  or _32222_ (_09203_, _09202_, _09198_);
  and _32223_ (_09204_, _09203_, _06021_);
  or _32224_ (_09205_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or _32225_ (_09206_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and _32226_ (_09207_, _09206_, _05997_);
  and _32227_ (_09208_, _09207_, _09205_);
  or _32228_ (_09209_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _32229_ (_09210_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and _32230_ (_09211_, _09210_, _05996_);
  and _32231_ (_09212_, _09211_, _09209_);
  or _32232_ (_09213_, _09212_, _09208_);
  and _32233_ (_09214_, _09213_, _05920_);
  or _32234_ (_09215_, _09214_, _09204_);
  and _32235_ (_09216_, _09215_, _05933_);
  and _32236_ (_09217_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and _32237_ (_09218_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _32238_ (_09219_, _09218_, _09217_);
  and _32239_ (_09220_, _09219_, _05996_);
  and _32240_ (_09221_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and _32241_ (_09222_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or _32242_ (_09223_, _09222_, _09221_);
  and _32243_ (_09224_, _09223_, _05997_);
  or _32244_ (_09225_, _09224_, _09220_);
  and _32245_ (_09226_, _09225_, _06021_);
  and _32246_ (_09227_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and _32247_ (_09228_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or _32248_ (_09229_, _09228_, _09227_);
  and _32249_ (_09230_, _09229_, _05996_);
  and _32250_ (_09231_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and _32251_ (_09232_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _32252_ (_09233_, _09232_, _09231_);
  and _32253_ (_09234_, _09233_, _05997_);
  or _32254_ (_09235_, _09234_, _09230_);
  and _32255_ (_09236_, _09235_, _05920_);
  or _32256_ (_09237_, _09236_, _09226_);
  and _32257_ (_09238_, _09237_, _06033_);
  or _32258_ (_09239_, _09238_, _09216_);
  and _32259_ (_09240_, _09239_, _06071_);
  or _32260_ (_09241_, _09240_, _09194_);
  and _32261_ (_09242_, _09241_, _05822_);
  or _32262_ (_09243_, _09242_, _09148_);
  or _32263_ (_09244_, _09243_, _06616_);
  and _32264_ (_09245_, _09244_, _09054_);
  or _32265_ (_09246_, _09245_, _05584_);
  and _32266_ (_09247_, _09246_, _08863_);
  or _32267_ (_09248_, _09247_, _06019_);
  not _32268_ (_09249_, _06019_);
  or _32269_ (_09250_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and _32270_ (_09251_, _09250_, _25365_);
  and _32271_ (_02659_, _09251_, _09248_);
  and _32272_ (_09252_, _06008_, _05777_);
  and _32273_ (_09253_, _06008_, _05824_);
  nor _32274_ (_09254_, _09253_, _09252_);
  nor _32275_ (_09255_, _05723_, _05516_);
  and _32276_ (_09256_, _09255_, _06008_);
  not _32277_ (_09257_, _09256_);
  and _32278_ (_09258_, _09257_, _09254_);
  nor _32279_ (_09259_, _06009_, _05726_);
  nor _32280_ (_09260_, _06009_, _06000_);
  nor _32281_ (_09261_, _09260_, _09259_);
  nor _32282_ (_09262_, _06009_, _05923_);
  nor _32283_ (_09263_, _06009_, _05930_);
  nor _32284_ (_09264_, _09263_, _09262_);
  and _32285_ (_09265_, _09264_, _09261_);
  and _32286_ (_09266_, _09265_, _06008_);
  and _32287_ (_09267_, _09266_, _09258_);
  not _32288_ (_09268_, _09267_);
  and _32289_ (_09269_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _32290_ (_09270_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _00986_);
  and _32291_ (_09271_, _09270_, _00973_);
  and _32292_ (_09272_, _09271_, _01344_);
  nor _32293_ (_09273_, _02259_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not _32294_ (_09274_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _32295_ (_09275_, _09271_, _09274_);
  and _32296_ (_09276_, _09275_, _00188_);
  or _32297_ (_09308_, _09276_, _09273_);
  or _32298_ (_09334_, _09308_, _09272_);
  and _32299_ (_09356_, _09334_, _09267_);
  or _32300_ (_12202_, _09356_, _09269_);
  and _32301_ (_09416_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nand _32302_ (_09443_, _09270_, _00979_);
  nor _32303_ (_09444_, _09443_, _01289_);
  and _32304_ (_09445_, _02251_, _09274_);
  and _32305_ (_09446_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _32306_ (_09447_, _09270_, _00981_);
  or _32307_ (_09448_, _09447_, _09446_);
  and _32308_ (_09449_, _09270_, _00976_);
  or _32309_ (_09450_, _09449_, _09448_);
  and _32310_ (_09451_, _09450_, _00137_);
  or _32311_ (_09452_, _09451_, _09445_);
  or _32312_ (_09453_, _09452_, _09444_);
  and _32313_ (_09454_, _09453_, _09267_);
  or _32314_ (_12204_, _09454_, _09416_);
  and _32315_ (_09455_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand _32316_ (_09456_, _09270_, _00977_);
  nor _32317_ (_09457_, _09456_, _01289_);
  and _32318_ (_09458_, _02236_, _09274_);
  nand _32319_ (_09459_, _00977_, _00986_);
  and _32320_ (_09460_, _00174_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _32321_ (_09461_, _09460_, _09459_);
  or _32322_ (_09462_, _09461_, _09458_);
  or _32323_ (_09463_, _09462_, _09457_);
  and _32324_ (_09464_, _09463_, _09267_);
  or _32325_ (_12205_, _09464_, _09455_);
  and _32326_ (_09465_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _32327_ (_09466_, _09447_, _01344_);
  and _32328_ (_09467_, _02220_, _09274_);
  nand _32329_ (_09468_, _00981_, _00986_);
  and _32330_ (_09469_, _00123_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _32331_ (_09470_, _09469_, _09468_);
  or _32332_ (_09471_, _09470_, _09467_);
  or _32333_ (_09472_, _09471_, _09466_);
  and _32334_ (_09473_, _09472_, _09267_);
  or _32335_ (_12207_, _09473_, _09465_);
  and _32336_ (_09474_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand _32337_ (_09475_, _09446_, _00973_);
  nor _32338_ (_09476_, _09475_, _01289_);
  nor _32339_ (_09477_, _02204_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _32340_ (_09478_, _00973_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _32341_ (_09479_, _00073_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _32342_ (_09480_, _09479_, _09478_);
  or _32343_ (_09481_, _09480_, _09477_);
  or _32344_ (_09482_, _09481_, _09476_);
  and _32345_ (_09483_, _09482_, _09267_);
  or _32346_ (_12208_, _09483_, _09474_);
  and _32347_ (_09484_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand _32348_ (_09485_, _09446_, _00979_);
  nor _32349_ (_09486_, _09485_, _01289_);
  nor _32350_ (_09487_, _02190_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _32351_ (_09488_, _00979_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _32352_ (_09489_, _00109_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _32353_ (_09490_, _09489_, _09488_);
  or _32354_ (_09491_, _09490_, _09487_);
  or _32355_ (_09492_, _09491_, _09486_);
  and _32356_ (_09493_, _09492_, _09267_);
  or _32357_ (_12210_, _09493_, _09484_);
  and _32358_ (_09494_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand _32359_ (_09495_, _09446_, _00977_);
  nor _32360_ (_09496_, _09495_, _01289_);
  nor _32361_ (_09497_, _02177_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _32362_ (_09498_, _00977_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _32363_ (_09499_, _00154_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _32364_ (_09500_, _09499_, _09498_);
  or _32365_ (_09501_, _09500_, _09497_);
  or _32366_ (_09502_, _09501_, _09496_);
  and _32367_ (_09503_, _09502_, _09267_);
  or _32368_ (_12211_, _09503_, _09494_);
  nand _32369_ (_09504_, _02280_, _09274_);
  and _32370_ (_09505_, _09446_, _00981_);
  nor _32371_ (_09506_, _00092_, _09274_);
  nor _32372_ (_09507_, _09506_, _09505_);
  and _32373_ (_09508_, _09507_, _09504_);
  and _32374_ (_09509_, _09505_, _01344_);
  or _32375_ (_09510_, _09509_, _09508_);
  and _32376_ (_09511_, _09510_, _09267_);
  and _32377_ (_09512_, _09268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _32378_ (_12213_, _09512_, _09511_);
  and _32379_ (_09513_, _09334_, _06008_);
  and _32380_ (_09514_, _09259_, _06000_);
  and _32381_ (_09515_, _09514_, _09264_);
  and _32382_ (_09516_, _09515_, _09258_);
  and _32383_ (_09517_, _09516_, _09513_);
  not _32384_ (_09518_, _09516_);
  and _32385_ (_09519_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _32386_ (_12214_, _09519_, _09517_);
  and _32387_ (_09520_, _09453_, _06008_);
  and _32388_ (_09521_, _09516_, _09520_);
  and _32389_ (_09522_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _32390_ (_12215_, _09522_, _09521_);
  and _32391_ (_09523_, _09463_, _06008_);
  and _32392_ (_09524_, _09516_, _09523_);
  and _32393_ (_09525_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _32394_ (_12216_, _09525_, _09524_);
  and _32395_ (_09526_, _09472_, _06008_);
  and _32396_ (_09527_, _09516_, _09526_);
  and _32397_ (_09528_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _32398_ (_12217_, _09528_, _09527_);
  and _32399_ (_09529_, _09482_, _06008_);
  and _32400_ (_09530_, _09516_, _09529_);
  and _32401_ (_09531_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or _32402_ (_12219_, _09531_, _09530_);
  and _32403_ (_09532_, _09492_, _06008_);
  and _32404_ (_09533_, _09516_, _09532_);
  and _32405_ (_09534_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _32406_ (_12220_, _09534_, _09533_);
  and _32407_ (_09535_, _09502_, _06008_);
  and _32408_ (_09536_, _09516_, _09535_);
  and _32409_ (_09537_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _32410_ (_12221_, _09537_, _09536_);
  and _32411_ (_09538_, _09510_, _06008_);
  and _32412_ (_09539_, _09516_, _09538_);
  and _32413_ (_09540_, _09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _32414_ (_12222_, _09540_, _09539_);
  and _32415_ (_09541_, _09260_, _05726_);
  and _32416_ (_09542_, _09541_, _09264_);
  and _32417_ (_09543_, _09542_, _09258_);
  and _32418_ (_09544_, _09543_, _09513_);
  not _32419_ (_09545_, _09543_);
  and _32420_ (_09546_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _32421_ (_12224_, _09546_, _09544_);
  and _32422_ (_09547_, _09543_, _09520_);
  and _32423_ (_09548_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _32424_ (_12225_, _09548_, _09547_);
  and _32425_ (_09549_, _09543_, _09523_);
  and _32426_ (_09550_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _32427_ (_12226_, _09550_, _09549_);
  and _32428_ (_09551_, _09543_, _09526_);
  and _32429_ (_09552_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _32430_ (_12227_, _09552_, _09551_);
  and _32431_ (_09553_, _09543_, _09529_);
  and _32432_ (_09554_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _32433_ (_12228_, _09554_, _09553_);
  and _32434_ (_09555_, _09543_, _09532_);
  and _32435_ (_09556_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _32436_ (_12230_, _09556_, _09555_);
  and _32437_ (_09557_, _09543_, _09535_);
  and _32438_ (_09558_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _32439_ (_12231_, _09558_, _09557_);
  and _32440_ (_09559_, _09543_, _09538_);
  and _32441_ (_09560_, _09545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _32442_ (_12232_, _09560_, _09559_);
  and _32443_ (_09561_, _09260_, _09259_);
  and _32444_ (_09562_, _09561_, _09264_);
  and _32445_ (_09563_, _09562_, _09258_);
  and _32446_ (_09564_, _09563_, _09513_);
  not _32447_ (_09565_, _09563_);
  and _32448_ (_09566_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _32449_ (_12234_, _09566_, _09564_);
  and _32450_ (_09567_, _09563_, _09520_);
  and _32451_ (_09568_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _32452_ (_12235_, _09568_, _09567_);
  and _32453_ (_09569_, _09563_, _09523_);
  and _32454_ (_09570_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _32455_ (_12236_, _09570_, _09569_);
  and _32456_ (_09571_, _09563_, _09526_);
  and _32457_ (_09572_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _32458_ (_12237_, _09572_, _09571_);
  and _32459_ (_09573_, _09563_, _09529_);
  and _32460_ (_09574_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _32461_ (_12238_, _09574_, _09573_);
  and _32462_ (_09575_, _09563_, _09532_);
  and _32463_ (_09576_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _32464_ (_12239_, _09576_, _09575_);
  and _32465_ (_09577_, _09563_, _09535_);
  and _32466_ (_09578_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _32467_ (_12241_, _09578_, _09577_);
  and _32468_ (_09579_, _09563_, _09538_);
  and _32469_ (_09580_, _09565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _32470_ (_12242_, _09580_, _09579_);
  and _32471_ (_09581_, _09262_, _05930_);
  and _32472_ (_09582_, _09581_, _09261_);
  and _32473_ (_09583_, _09582_, _09258_);
  and _32474_ (_09584_, _09583_, _09513_);
  not _32475_ (_09585_, _09583_);
  and _32476_ (_09586_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _32477_ (_12244_, _09586_, _09584_);
  and _32478_ (_09587_, _09583_, _09520_);
  and _32479_ (_09588_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _32480_ (_12245_, _09588_, _09587_);
  and _32481_ (_09589_, _09583_, _09523_);
  and _32482_ (_09590_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _32483_ (_12246_, _09590_, _09589_);
  and _32484_ (_09591_, _09583_, _09526_);
  and _32485_ (_09592_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _32486_ (_12247_, _09592_, _09591_);
  and _32487_ (_09593_, _09583_, _09529_);
  and _32488_ (_09594_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _32489_ (_12248_, _09594_, _09593_);
  and _32490_ (_09595_, _09583_, _09532_);
  and _32491_ (_09596_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _32492_ (_12249_, _09596_, _09595_);
  and _32493_ (_09597_, _09583_, _09535_);
  and _32494_ (_09598_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _32495_ (_12250_, _09598_, _09597_);
  and _32496_ (_09599_, _09583_, _09538_);
  and _32497_ (_09600_, _09585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _32498_ (_12252_, _09600_, _09599_);
  and _32499_ (_09601_, _09581_, _09514_);
  and _32500_ (_09602_, _09601_, _09258_);
  and _32501_ (_09603_, _09602_, _09513_);
  not _32502_ (_09604_, _09602_);
  and _32503_ (_09605_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _32504_ (_12253_, _09605_, _09603_);
  and _32505_ (_09606_, _09602_, _09520_);
  and _32506_ (_09607_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _32507_ (_12254_, _09607_, _09606_);
  and _32508_ (_09608_, _09602_, _09523_);
  and _32509_ (_09609_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _32510_ (_12256_, _09609_, _09608_);
  and _32511_ (_09610_, _09602_, _09526_);
  and _32512_ (_09611_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _32513_ (_12257_, _09611_, _09610_);
  and _32514_ (_09612_, _09602_, _09529_);
  and _32515_ (_09613_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or _32516_ (_12258_, _09613_, _09612_);
  and _32517_ (_09614_, _09602_, _09532_);
  and _32518_ (_09615_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or _32519_ (_12259_, _09615_, _09614_);
  and _32520_ (_09616_, _09602_, _09535_);
  and _32521_ (_09617_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or _32522_ (_12260_, _09617_, _09616_);
  and _32523_ (_09618_, _09602_, _09538_);
  and _32524_ (_09619_, _09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _32525_ (_12261_, _09619_, _09618_);
  and _32526_ (_09620_, _09581_, _09541_);
  and _32527_ (_09621_, _09620_, _09258_);
  and _32528_ (_09622_, _09621_, _09513_);
  not _32529_ (_09623_, _09621_);
  and _32530_ (_09624_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _32531_ (_12263_, _09624_, _09622_);
  and _32532_ (_09625_, _09621_, _09520_);
  and _32533_ (_09626_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _32534_ (_12264_, _09626_, _09625_);
  and _32535_ (_09627_, _09621_, _09523_);
  and _32536_ (_09628_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _32537_ (_12265_, _09628_, _09627_);
  and _32538_ (_09629_, _09621_, _09526_);
  and _32539_ (_09630_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _32540_ (_12266_, _09630_, _09629_);
  and _32541_ (_09631_, _09621_, _09529_);
  and _32542_ (_09632_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _32543_ (_12268_, _09632_, _09631_);
  and _32544_ (_09633_, _09621_, _09532_);
  and _32545_ (_09634_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _32546_ (_12269_, _09634_, _09633_);
  and _32547_ (_09635_, _09621_, _09535_);
  and _32548_ (_09636_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _32549_ (_12270_, _09636_, _09635_);
  and _32550_ (_09637_, _09621_, _09538_);
  and _32551_ (_09638_, _09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _32552_ (_12271_, _09638_, _09637_);
  and _32553_ (_09639_, _09581_, _09561_);
  and _32554_ (_09640_, _09639_, _09258_);
  and _32555_ (_09641_, _09640_, _09513_);
  not _32556_ (_09642_, _09640_);
  and _32557_ (_09643_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _32558_ (_12272_, _09643_, _09641_);
  and _32559_ (_09644_, _09640_, _09520_);
  and _32560_ (_09645_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _32561_ (_12273_, _09645_, _09644_);
  and _32562_ (_09646_, _09640_, _09523_);
  and _32563_ (_09647_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _32564_ (_12275_, _09647_, _09646_);
  and _32565_ (_09648_, _09640_, _09526_);
  and _32566_ (_09649_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _32567_ (_12276_, _09649_, _09648_);
  and _32568_ (_09650_, _09640_, _09529_);
  and _32569_ (_09651_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _32570_ (_12277_, _09651_, _09650_);
  and _32571_ (_09652_, _09640_, _09532_);
  and _32572_ (_09653_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _32573_ (_12279_, _09653_, _09652_);
  and _32574_ (_09654_, _09640_, _09535_);
  and _32575_ (_09655_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _32576_ (_12280_, _09655_, _09654_);
  and _32577_ (_09656_, _09640_, _09538_);
  and _32578_ (_09657_, _09642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _32579_ (_12281_, _09657_, _09656_);
  and _32580_ (_09658_, _09263_, _05923_);
  and _32581_ (_09659_, _09658_, _09261_);
  and _32582_ (_09660_, _09659_, _09258_);
  and _32583_ (_09661_, _09660_, _09513_);
  not _32584_ (_09662_, _09660_);
  and _32585_ (_09663_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _32586_ (_12282_, _09663_, _09661_);
  and _32587_ (_09664_, _09660_, _09520_);
  and _32588_ (_09665_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _32589_ (_12283_, _09665_, _09664_);
  and _32590_ (_09666_, _09660_, _09523_);
  and _32591_ (_09667_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _32592_ (_12284_, _09667_, _09666_);
  and _32593_ (_09668_, _09660_, _09526_);
  and _32594_ (_09669_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _32595_ (_12286_, _09669_, _09668_);
  and _32596_ (_09670_, _09660_, _09529_);
  and _32597_ (_09671_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _32598_ (_12287_, _09671_, _09670_);
  and _32599_ (_09672_, _09660_, _09532_);
  and _32600_ (_09673_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _32601_ (_12288_, _09673_, _09672_);
  and _32602_ (_09674_, _09660_, _09535_);
  and _32603_ (_09675_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or _32604_ (_12290_, _09675_, _09674_);
  and _32605_ (_09676_, _09660_, _09538_);
  and _32606_ (_09677_, _09662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _32607_ (_12291_, _09677_, _09676_);
  and _32608_ (_09678_, _09658_, _09514_);
  and _32609_ (_09679_, _09678_, _09258_);
  and _32610_ (_09680_, _09679_, _09513_);
  not _32611_ (_09681_, _09679_);
  and _32612_ (_09682_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _32613_ (_12292_, _09682_, _09680_);
  and _32614_ (_09683_, _09679_, _09520_);
  and _32615_ (_09684_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _32616_ (_12293_, _09684_, _09683_);
  and _32617_ (_09685_, _09679_, _09523_);
  and _32618_ (_09686_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _32619_ (_12294_, _09686_, _09685_);
  and _32620_ (_09687_, _09679_, _09526_);
  and _32621_ (_09688_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _32622_ (_12295_, _09688_, _09687_);
  and _32623_ (_09689_, _09679_, _09529_);
  and _32624_ (_09690_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _32625_ (_12297_, _09690_, _09689_);
  and _32626_ (_09691_, _09679_, _09532_);
  and _32627_ (_09692_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _32628_ (_12298_, _09692_, _09691_);
  and _32629_ (_09693_, _09679_, _09535_);
  and _32630_ (_09694_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _32631_ (_12299_, _09694_, _09693_);
  and _32632_ (_09695_, _09679_, _09538_);
  and _32633_ (_09696_, _09681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _32634_ (_12300_, _09696_, _09695_);
  and _32635_ (_09697_, _09658_, _09541_);
  and _32636_ (_09698_, _09697_, _09258_);
  and _32637_ (_09699_, _09698_, _09513_);
  not _32638_ (_09700_, _09698_);
  and _32639_ (_09701_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _32640_ (_12302_, _09701_, _09699_);
  and _32641_ (_09702_, _09698_, _09520_);
  and _32642_ (_09703_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _32643_ (_12303_, _09703_, _09702_);
  and _32644_ (_09704_, _09698_, _09523_);
  and _32645_ (_09705_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _32646_ (_12304_, _09705_, _09704_);
  and _32647_ (_09706_, _09698_, _09526_);
  and _32648_ (_09707_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _32649_ (_12306_, _09707_, _09706_);
  and _32650_ (_09708_, _09698_, _09529_);
  and _32651_ (_09709_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _32652_ (_12307_, _09709_, _09708_);
  and _32653_ (_09710_, _09698_, _09532_);
  and _32654_ (_09711_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _32655_ (_12308_, _09711_, _09710_);
  and _32656_ (_09712_, _09698_, _09535_);
  and _32657_ (_09713_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _32658_ (_12310_, _09713_, _09712_);
  and _32659_ (_09714_, _09698_, _09538_);
  and _32660_ (_09715_, _09700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _32661_ (_12311_, _09715_, _09714_);
  and _32662_ (_09716_, _09658_, _09561_);
  and _32663_ (_09717_, _09716_, _09258_);
  and _32664_ (_09718_, _09717_, _09513_);
  not _32665_ (_09719_, _09717_);
  and _32666_ (_09720_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or _32667_ (_12312_, _09720_, _09718_);
  and _32668_ (_09721_, _09717_, _09520_);
  and _32669_ (_09722_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _32670_ (_12313_, _09722_, _09721_);
  and _32671_ (_09723_, _09717_, _09523_);
  and _32672_ (_09724_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _32673_ (_12314_, _09724_, _09723_);
  and _32674_ (_09725_, _09717_, _09526_);
  and _32675_ (_09726_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _32676_ (_12315_, _09726_, _09725_);
  and _32677_ (_09727_, _09717_, _09529_);
  and _32678_ (_09728_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or _32679_ (_12317_, _09728_, _09727_);
  and _32680_ (_09729_, _09717_, _09532_);
  and _32681_ (_09730_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _32682_ (_12318_, _09730_, _09729_);
  and _32683_ (_09731_, _09717_, _09535_);
  and _32684_ (_09732_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _32685_ (_12319_, _09732_, _09731_);
  and _32686_ (_09733_, _09717_, _09538_);
  and _32687_ (_09734_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _32688_ (_12320_, _09734_, _09733_);
  and _32689_ (_09735_, _09263_, _09262_);
  and _32690_ (_09736_, _09735_, _09261_);
  and _32691_ (_09737_, _09736_, _09258_);
  and _32692_ (_09738_, _09737_, _09513_);
  not _32693_ (_09739_, _09737_);
  and _32694_ (_09740_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _32695_ (_12322_, _09740_, _09738_);
  and _32696_ (_09741_, _09737_, _09520_);
  and _32697_ (_09742_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _32698_ (_12323_, _09742_, _09741_);
  and _32699_ (_09743_, _09737_, _09523_);
  and _32700_ (_09744_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _32701_ (_12324_, _09744_, _09743_);
  and _32702_ (_09745_, _09737_, _09526_);
  and _32703_ (_09746_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or _32704_ (_12325_, _09746_, _09745_);
  and _32705_ (_09747_, _09737_, _09529_);
  and _32706_ (_09748_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _32707_ (_12326_, _09748_, _09747_);
  and _32708_ (_09749_, _09737_, _09532_);
  and _32709_ (_09750_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _32710_ (_12327_, _09750_, _09749_);
  and _32711_ (_09751_, _09737_, _09535_);
  and _32712_ (_09752_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _32713_ (_12329_, _09752_, _09751_);
  and _32714_ (_09753_, _09737_, _09538_);
  and _32715_ (_09754_, _09739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _32716_ (_12330_, _09754_, _09753_);
  and _32717_ (_09755_, _09735_, _09514_);
  and _32718_ (_09756_, _09755_, _09258_);
  and _32719_ (_09757_, _09756_, _09513_);
  not _32720_ (_09758_, _09756_);
  and _32721_ (_09759_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _32722_ (_12331_, _09759_, _09757_);
  and _32723_ (_09760_, _09756_, _09520_);
  and _32724_ (_09761_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _32725_ (_12333_, _09761_, _09760_);
  and _32726_ (_09762_, _09756_, _09523_);
  and _32727_ (_09763_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _32728_ (_12334_, _09763_, _09762_);
  and _32729_ (_09764_, _09756_, _09526_);
  and _32730_ (_09765_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _32731_ (_12335_, _09765_, _09764_);
  and _32732_ (_09766_, _09756_, _09529_);
  and _32733_ (_09767_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _32734_ (_12336_, _09767_, _09766_);
  and _32735_ (_09768_, _09756_, _09532_);
  and _32736_ (_09769_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _32737_ (_12337_, _09769_, _09768_);
  and _32738_ (_09770_, _09756_, _09535_);
  and _32739_ (_09771_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _32740_ (_12338_, _09771_, _09770_);
  and _32741_ (_09772_, _09756_, _09538_);
  and _32742_ (_09773_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _32743_ (_12339_, _09773_, _09772_);
  and _32744_ (_09774_, _09735_, _09541_);
  and _32745_ (_09775_, _09774_, _09258_);
  and _32746_ (_09776_, _09775_, _09513_);
  not _32747_ (_09777_, _09775_);
  and _32748_ (_09778_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _32749_ (_12341_, _09778_, _09776_);
  and _32750_ (_09779_, _09775_, _09520_);
  and _32751_ (_09780_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _32752_ (_12342_, _09780_, _09779_);
  and _32753_ (_09781_, _09775_, _09523_);
  and _32754_ (_09782_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _32755_ (_12344_, _09782_, _09781_);
  and _32756_ (_09783_, _09775_, _09526_);
  and _32757_ (_09784_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _32758_ (_12345_, _09784_, _09783_);
  and _32759_ (_09785_, _09775_, _09529_);
  and _32760_ (_09786_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _32761_ (_12346_, _09786_, _09785_);
  and _32762_ (_09787_, _09775_, _09532_);
  and _32763_ (_09788_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _32764_ (_12347_, _09788_, _09787_);
  and _32765_ (_09789_, _09775_, _09535_);
  and _32766_ (_09790_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _32767_ (_12348_, _09790_, _09789_);
  and _32768_ (_09791_, _09775_, _09538_);
  and _32769_ (_09792_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _32770_ (_12349_, _09792_, _09791_);
  and _32771_ (_09793_, _09735_, _09561_);
  and _32772_ (_09794_, _09793_, _09258_);
  and _32773_ (_09795_, _09794_, _09513_);
  not _32774_ (_09796_, _09794_);
  and _32775_ (_09797_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _32776_ (_12350_, _09797_, _09795_);
  and _32777_ (_09798_, _09794_, _09520_);
  and _32778_ (_09799_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _32779_ (_12352_, _09799_, _09798_);
  and _32780_ (_09800_, _09794_, _09523_);
  and _32781_ (_09801_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or _32782_ (_12353_, _09801_, _09800_);
  and _32783_ (_09802_, _09794_, _09526_);
  and _32784_ (_09803_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _32785_ (_12354_, _09803_, _09802_);
  and _32786_ (_09804_, _09794_, _09529_);
  and _32787_ (_09805_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or _32788_ (_12356_, _09805_, _09804_);
  and _32789_ (_09806_, _09794_, _09532_);
  and _32790_ (_09807_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _32791_ (_12357_, _09807_, _09806_);
  and _32792_ (_09808_, _09794_, _09535_);
  and _32793_ (_09809_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _32794_ (_12358_, _09809_, _09808_);
  and _32795_ (_09810_, _09794_, _09538_);
  and _32796_ (_09811_, _09796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _32797_ (_12359_, _09811_, _09810_);
  not _32798_ (_09812_, _09255_);
  and _32799_ (_09813_, _09252_, _00892_);
  and _32800_ (_09814_, _09813_, _09812_);
  and _32801_ (_09815_, _09814_, _09265_);
  and _32802_ (_09816_, _09815_, _09513_);
  not _32803_ (_09817_, _09815_);
  and _32804_ (_09818_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or _32805_ (_12360_, _09818_, _09816_);
  and _32806_ (_09819_, _09815_, _09520_);
  and _32807_ (_09820_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or _32808_ (_12362_, _09820_, _09819_);
  and _32809_ (_09821_, _09815_, _09523_);
  and _32810_ (_09822_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or _32811_ (_12363_, _09822_, _09821_);
  and _32812_ (_09823_, _09815_, _09526_);
  and _32813_ (_09824_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or _32814_ (_12364_, _09824_, _09823_);
  and _32815_ (_09825_, _09815_, _09529_);
  and _32816_ (_09826_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or _32817_ (_12365_, _09826_, _09825_);
  and _32818_ (_09827_, _09815_, _09532_);
  and _32819_ (_09828_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or _32820_ (_12367_, _09828_, _09827_);
  and _32821_ (_09829_, _09815_, _09535_);
  and _32822_ (_09830_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or _32823_ (_12368_, _09830_, _09829_);
  and _32824_ (_09831_, _09815_, _09538_);
  and _32825_ (_09832_, _09817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or _32826_ (_12369_, _09832_, _09831_);
  and _32827_ (_09833_, _09814_, _09515_);
  and _32828_ (_09834_, _09833_, _09513_);
  not _32829_ (_09835_, _09833_);
  and _32830_ (_09836_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _32831_ (_12370_, _09836_, _09834_);
  and _32832_ (_09837_, _09833_, _09520_);
  and _32833_ (_09838_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _32834_ (_12371_, _09838_, _09837_);
  and _32835_ (_09839_, _09833_, _09523_);
  and _32836_ (_09840_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _32837_ (_12372_, _09840_, _09839_);
  and _32838_ (_09841_, _09833_, _09526_);
  and _32839_ (_09842_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _32840_ (_12374_, _09842_, _09841_);
  and _32841_ (_09843_, _09833_, _09529_);
  and _32842_ (_09844_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _32843_ (_12375_, _09844_, _09843_);
  and _32844_ (_09845_, _09833_, _09532_);
  and _32845_ (_09846_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _32846_ (_12376_, _09846_, _09845_);
  and _32847_ (_09847_, _09833_, _09535_);
  and _32848_ (_09848_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _32849_ (_12377_, _09848_, _09847_);
  and _32850_ (_09849_, _09833_, _09538_);
  and _32851_ (_09850_, _09835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _32852_ (_12379_, _09850_, _09849_);
  and _32853_ (_09851_, _09814_, _09542_);
  and _32854_ (_09852_, _09851_, _09513_);
  not _32855_ (_09853_, _09851_);
  and _32856_ (_09854_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _32857_ (_12380_, _09854_, _09852_);
  and _32858_ (_09855_, _09851_, _09520_);
  and _32859_ (_09856_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _32860_ (_12381_, _09856_, _09855_);
  and _32861_ (_09857_, _09851_, _09523_);
  and _32862_ (_09858_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _32863_ (_12382_, _09858_, _09857_);
  and _32864_ (_09859_, _09851_, _09526_);
  and _32865_ (_09860_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _32866_ (_12383_, _09860_, _09859_);
  and _32867_ (_09861_, _09851_, _09529_);
  and _32868_ (_09862_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _32869_ (_12384_, _09862_, _09861_);
  and _32870_ (_09863_, _09851_, _09532_);
  and _32871_ (_09864_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _32872_ (_12386_, _09864_, _09863_);
  and _32873_ (_09865_, _09851_, _09535_);
  and _32874_ (_09866_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _32875_ (_12387_, _09866_, _09865_);
  and _32876_ (_09867_, _09851_, _09538_);
  and _32877_ (_09868_, _09853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _32878_ (_12388_, _09868_, _09867_);
  and _32879_ (_09869_, _09814_, _09562_);
  and _32880_ (_09870_, _09869_, _09513_);
  not _32881_ (_09871_, _09869_);
  and _32882_ (_09872_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or _32883_ (_12389_, _09872_, _09870_);
  and _32884_ (_09873_, _09869_, _09520_);
  and _32885_ (_09874_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or _32886_ (_12391_, _09874_, _09873_);
  and _32887_ (_09875_, _09869_, _09523_);
  and _32888_ (_09876_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or _32889_ (_12392_, _09876_, _09875_);
  and _32890_ (_09877_, _09869_, _09526_);
  and _32891_ (_09878_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or _32892_ (_12393_, _09878_, _09877_);
  and _32893_ (_09879_, _09869_, _09529_);
  and _32894_ (_09880_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or _32895_ (_12394_, _09880_, _09879_);
  and _32896_ (_09881_, _09869_, _09532_);
  and _32897_ (_09882_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or _32898_ (_12395_, _09882_, _09881_);
  and _32899_ (_09883_, _09869_, _09535_);
  and _32900_ (_09884_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or _32901_ (_12396_, _09884_, _09883_);
  and _32902_ (_09885_, _09869_, _09538_);
  and _32903_ (_09886_, _09871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or _32904_ (_12397_, _09886_, _09885_);
  and _32905_ (_09887_, _09814_, _09582_);
  and _32906_ (_09888_, _09887_, _09513_);
  not _32907_ (_09889_, _09887_);
  and _32908_ (_09890_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or _32909_ (_12399_, _09890_, _09888_);
  and _32910_ (_09891_, _09887_, _09520_);
  and _32911_ (_09892_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or _32912_ (_12400_, _09892_, _09891_);
  and _32913_ (_09893_, _09887_, _09523_);
  and _32914_ (_09894_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or _32915_ (_12401_, _09894_, _09893_);
  and _32916_ (_09895_, _09887_, _09526_);
  and _32917_ (_09896_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or _32918_ (_12403_, _09896_, _09895_);
  and _32919_ (_09897_, _09887_, _09529_);
  and _32920_ (_09898_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or _32921_ (_12404_, _09898_, _09897_);
  and _32922_ (_09899_, _09887_, _09532_);
  and _32923_ (_09900_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or _32924_ (_12405_, _09900_, _09899_);
  and _32925_ (_09901_, _09887_, _09535_);
  and _32926_ (_09902_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or _32927_ (_12407_, _09902_, _09901_);
  and _32928_ (_09903_, _09887_, _09538_);
  and _32929_ (_09904_, _09889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or _32930_ (_12408_, _09904_, _09903_);
  and _32931_ (_09905_, _09814_, _09601_);
  and _32932_ (_09906_, _09905_, _09513_);
  not _32933_ (_09907_, _09905_);
  and _32934_ (_09908_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _32935_ (_12409_, _09908_, _09906_);
  and _32936_ (_09909_, _09905_, _09520_);
  and _32937_ (_09910_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _32938_ (_12411_, _09910_, _09909_);
  and _32939_ (_09911_, _09905_, _09523_);
  and _32940_ (_09912_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _32941_ (_12412_, _09912_, _09911_);
  and _32942_ (_09913_, _09905_, _09526_);
  and _32943_ (_09914_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _32944_ (_12413_, _09914_, _09913_);
  and _32945_ (_09915_, _09905_, _09529_);
  and _32946_ (_09916_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _32947_ (_12414_, _09916_, _09915_);
  and _32948_ (_09917_, _09905_, _09532_);
  and _32949_ (_09918_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _32950_ (_12415_, _09918_, _09917_);
  and _32951_ (_09919_, _09905_, _09535_);
  and _32952_ (_09920_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _32953_ (_12416_, _09920_, _09919_);
  and _32954_ (_09921_, _09905_, _09538_);
  and _32955_ (_09922_, _09907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _32956_ (_12417_, _09922_, _09921_);
  and _32957_ (_09923_, _09814_, _09620_);
  and _32958_ (_09924_, _09923_, _09513_);
  not _32959_ (_09925_, _09923_);
  and _32960_ (_09926_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _32961_ (_12419_, _09926_, _09924_);
  and _32962_ (_09927_, _09923_, _09520_);
  and _32963_ (_09928_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _32964_ (_12420_, _09928_, _09927_);
  and _32965_ (_09929_, _09923_, _09523_);
  and _32966_ (_09930_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _32967_ (_12421_, _09930_, _09929_);
  and _32968_ (_09931_, _09923_, _09526_);
  and _32969_ (_09932_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _32970_ (_12423_, _09932_, _09931_);
  and _32971_ (_09933_, _09923_, _09529_);
  and _32972_ (_09934_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _32973_ (_12424_, _09934_, _09933_);
  and _32974_ (_09935_, _09923_, _09532_);
  and _32975_ (_09936_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _32976_ (_12425_, _09936_, _09935_);
  and _32977_ (_09937_, _09923_, _09535_);
  and _32978_ (_09938_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _32979_ (_12426_, _09938_, _09937_);
  and _32980_ (_09939_, _09923_, _09538_);
  and _32981_ (_09940_, _09925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _32982_ (_12427_, _09940_, _09939_);
  and _32983_ (_09941_, _09814_, _09639_);
  and _32984_ (_09942_, _09941_, _09513_);
  not _32985_ (_09943_, _09941_);
  and _32986_ (_09944_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or _32987_ (_12428_, _09944_, _09942_);
  and _32988_ (_09945_, _09941_, _09520_);
  and _32989_ (_09946_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or _32990_ (_12429_, _09946_, _09945_);
  and _32991_ (_09947_, _09941_, _09523_);
  and _32992_ (_09948_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or _32993_ (_12431_, _09948_, _09947_);
  and _32994_ (_09949_, _09941_, _09526_);
  and _32995_ (_09950_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or _32996_ (_12432_, _09950_, _09949_);
  and _32997_ (_09951_, _09941_, _09529_);
  and _32998_ (_09952_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or _32999_ (_12433_, _09952_, _09951_);
  and _33000_ (_09953_, _09941_, _09532_);
  and _33001_ (_09954_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or _33002_ (_12435_, _09954_, _09953_);
  and _33003_ (_09955_, _09941_, _09535_);
  and _33004_ (_09956_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or _33005_ (_12436_, _09956_, _09955_);
  and _33006_ (_09957_, _09941_, _09538_);
  and _33007_ (_09958_, _09943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or _33008_ (_12437_, _09958_, _09957_);
  and _33009_ (_09959_, _09814_, _09659_);
  and _33010_ (_09960_, _09959_, _09513_);
  not _33011_ (_09961_, _09959_);
  and _33012_ (_09962_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _33013_ (_12438_, _09962_, _09960_);
  and _33014_ (_09963_, _09959_, _09520_);
  and _33015_ (_09964_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _33016_ (_12439_, _09964_, _09963_);
  and _33017_ (_09965_, _09959_, _09523_);
  and _33018_ (_09966_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _33019_ (_12440_, _09966_, _09965_);
  and _33020_ (_09967_, _09959_, _09526_);
  and _33021_ (_09968_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _33022_ (_12441_, _09968_, _09967_);
  and _33023_ (_09969_, _09959_, _09529_);
  and _33024_ (_09970_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _33025_ (_12443_, _09970_, _09969_);
  and _33026_ (_09971_, _09959_, _09532_);
  and _33027_ (_09972_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _33028_ (_12444_, _09972_, _09971_);
  and _33029_ (_09973_, _09959_, _09535_);
  and _33030_ (_09974_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _33031_ (_12445_, _09974_, _09973_);
  and _33032_ (_09975_, _09959_, _09538_);
  and _33033_ (_09976_, _09961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _33034_ (_12446_, _09976_, _09975_);
  and _33035_ (_09977_, _09814_, _09678_);
  and _33036_ (_09978_, _09977_, _09513_);
  not _33037_ (_09979_, _09977_);
  and _33038_ (_09980_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or _33039_ (_12448_, _09980_, _09978_);
  and _33040_ (_09981_, _09977_, _09520_);
  and _33041_ (_09982_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or _33042_ (_12449_, _09982_, _09981_);
  and _33043_ (_09983_, _09977_, _09523_);
  and _33044_ (_09984_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or _33045_ (_12450_, _09984_, _09983_);
  and _33046_ (_09985_, _09977_, _09526_);
  and _33047_ (_09986_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or _33048_ (_12451_, _09986_, _09985_);
  and _33049_ (_09987_, _09977_, _09529_);
  and _33050_ (_09988_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or _33051_ (_12452_, _09988_, _09987_);
  and _33052_ (_09989_, _09977_, _09532_);
  and _33053_ (_09990_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or _33054_ (_12453_, _09990_, _09989_);
  and _33055_ (_09991_, _09977_, _09535_);
  and _33056_ (_09992_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or _33057_ (_12455_, _09992_, _09991_);
  and _33058_ (_09993_, _09977_, _09538_);
  and _33059_ (_09994_, _09979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or _33060_ (_12456_, _09994_, _09993_);
  and _33061_ (_09995_, _09814_, _09697_);
  and _33062_ (_09996_, _09995_, _09513_);
  not _33063_ (_09997_, _09995_);
  and _33064_ (_09998_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or _33065_ (_12457_, _09998_, _09996_);
  and _33066_ (_09999_, _09995_, _09520_);
  and _33067_ (_10000_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or _33068_ (_12459_, _10000_, _09999_);
  and _33069_ (_10001_, _09995_, _09523_);
  and _33070_ (_10002_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or _33071_ (_12460_, _10002_, _10001_);
  and _33072_ (_10003_, _09995_, _09526_);
  and _33073_ (_10004_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or _33074_ (_12461_, _10004_, _10003_);
  and _33075_ (_10005_, _09995_, _09529_);
  and _33076_ (_10006_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or _33077_ (_12462_, _10006_, _10005_);
  and _33078_ (_10007_, _09995_, _09532_);
  and _33079_ (_10008_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or _33080_ (_12463_, _10008_, _10007_);
  and _33081_ (_10009_, _09995_, _09535_);
  and _33082_ (_10010_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or _33083_ (_12464_, _10010_, _10009_);
  and _33084_ (_10011_, _09995_, _09538_);
  and _33085_ (_10012_, _09997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or _33086_ (_12465_, _10012_, _10011_);
  and _33087_ (_10013_, _09814_, _09716_);
  and _33088_ (_10014_, _10013_, _09513_);
  not _33089_ (_10015_, _10013_);
  and _33090_ (_10016_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _33091_ (_12467_, _10016_, _10014_);
  and _33092_ (_10017_, _10013_, _09520_);
  and _33093_ (_10018_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _33094_ (_12468_, _10018_, _10017_);
  and _33095_ (_10019_, _10013_, _09523_);
  and _33096_ (_10020_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _33097_ (_12469_, _10020_, _10019_);
  and _33098_ (_10021_, _10013_, _09526_);
  and _33099_ (_10022_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _33100_ (_12471_, _10022_, _10021_);
  and _33101_ (_10023_, _10013_, _09529_);
  and _33102_ (_10024_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _33103_ (_12472_, _10024_, _10023_);
  and _33104_ (_10025_, _10013_, _09532_);
  and _33105_ (_10026_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _33106_ (_12473_, _10026_, _10025_);
  and _33107_ (_10027_, _10013_, _09535_);
  and _33108_ (_10028_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _33109_ (_12474_, _10028_, _10027_);
  and _33110_ (_10029_, _10013_, _09538_);
  and _33111_ (_10030_, _10015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _33112_ (_12475_, _10030_, _10029_);
  and _33113_ (_10031_, _09814_, _09736_);
  and _33114_ (_10032_, _10031_, _09513_);
  not _33115_ (_10033_, _10031_);
  and _33116_ (_10034_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _33117_ (_12476_, _10034_, _10032_);
  and _33118_ (_10035_, _10031_, _09520_);
  and _33119_ (_10036_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _33120_ (_12477_, _10036_, _10035_);
  and _33121_ (_10037_, _10031_, _09523_);
  and _33122_ (_10038_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _33123_ (_12479_, _10038_, _10037_);
  and _33124_ (_10039_, _10031_, _09526_);
  and _33125_ (_10040_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _33126_ (_12480_, _10040_, _10039_);
  and _33127_ (_10041_, _10031_, _09529_);
  and _33128_ (_10042_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _33129_ (_12481_, _10042_, _10041_);
  and _33130_ (_10043_, _10031_, _09532_);
  and _33131_ (_10044_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _33132_ (_12483_, _10044_, _10043_);
  and _33133_ (_10045_, _10031_, _09535_);
  and _33134_ (_10046_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _33135_ (_12484_, _10046_, _10045_);
  and _33136_ (_10047_, _10031_, _09538_);
  and _33137_ (_10048_, _10033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _33138_ (_12485_, _10048_, _10047_);
  and _33139_ (_10049_, _09814_, _09755_);
  and _33140_ (_10050_, _10049_, _09513_);
  not _33141_ (_10051_, _10049_);
  and _33142_ (_10052_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or _33143_ (_12486_, _10052_, _10050_);
  and _33144_ (_10053_, _10049_, _09520_);
  and _33145_ (_10054_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or _33146_ (_12487_, _10054_, _10053_);
  and _33147_ (_10055_, _10049_, _09523_);
  and _33148_ (_10056_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or _33149_ (_12488_, _10056_, _10055_);
  and _33150_ (_10057_, _10049_, _09526_);
  and _33151_ (_10058_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or _33152_ (_12489_, _10058_, _10057_);
  and _33153_ (_10059_, _10049_, _09529_);
  and _33154_ (_10060_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or _33155_ (_12491_, _10060_, _10059_);
  and _33156_ (_10061_, _10049_, _09532_);
  and _33157_ (_10062_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or _33158_ (_12492_, _10062_, _10061_);
  and _33159_ (_10063_, _10049_, _09535_);
  and _33160_ (_10064_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or _33161_ (_12493_, _10064_, _10063_);
  and _33162_ (_10065_, _10049_, _09538_);
  and _33163_ (_10066_, _10051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or _33164_ (_12494_, _10066_, _10065_);
  and _33165_ (_10067_, _09814_, _09774_);
  and _33166_ (_10068_, _10067_, _09513_);
  not _33167_ (_10069_, _10067_);
  and _33168_ (_10070_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or _33169_ (_12496_, _10070_, _10068_);
  and _33170_ (_10071_, _10067_, _09520_);
  and _33171_ (_10072_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or _33172_ (_12497_, _10072_, _10071_);
  and _33173_ (_10073_, _10067_, _09523_);
  and _33174_ (_10074_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or _33175_ (_12498_, _10074_, _10073_);
  and _33176_ (_10075_, _10067_, _09526_);
  and _33177_ (_10076_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or _33178_ (_12499_, _10076_, _10075_);
  and _33179_ (_10077_, _10067_, _09529_);
  and _33180_ (_10078_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or _33181_ (_12500_, _10078_, _10077_);
  and _33182_ (_10079_, _10067_, _09532_);
  and _33183_ (_10080_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or _33184_ (_12501_, _10080_, _10079_);
  and _33185_ (_10081_, _10067_, _09535_);
  and _33186_ (_10082_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or _33187_ (_12503_, _10082_, _10081_);
  and _33188_ (_10083_, _10067_, _09538_);
  and _33189_ (_10084_, _10069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or _33190_ (_12504_, _10084_, _10083_);
  and _33191_ (_10085_, _09814_, _09793_);
  and _33192_ (_10086_, _10085_, _09513_);
  not _33193_ (_10087_, _10085_);
  and _33194_ (_10088_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _33195_ (_12505_, _10088_, _10086_);
  and _33196_ (_10089_, _10085_, _09520_);
  and _33197_ (_10090_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _33198_ (_12507_, _10090_, _10089_);
  and _33199_ (_10091_, _10085_, _09523_);
  and _33200_ (_10092_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _33201_ (_12508_, _10092_, _10091_);
  and _33202_ (_10093_, _10085_, _09526_);
  and _33203_ (_10094_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _33204_ (_12509_, _10094_, _10093_);
  and _33205_ (_10095_, _10085_, _09529_);
  and _33206_ (_10096_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _33207_ (_12510_, _10096_, _10095_);
  and _33208_ (_10097_, _10085_, _09532_);
  and _33209_ (_10098_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _33210_ (_12512_, _10098_, _10097_);
  and _33211_ (_10099_, _10085_, _09535_);
  and _33212_ (_10100_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _33213_ (_12513_, _10100_, _10099_);
  and _33214_ (_10101_, _10085_, _09538_);
  and _33215_ (_10102_, _10087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _33216_ (_12514_, _10102_, _10101_);
  and _33217_ (_10103_, _09253_, _05778_);
  and _33218_ (_10104_, _10103_, _09812_);
  and _33219_ (_10105_, _10104_, _09265_);
  and _33220_ (_10106_, _10105_, _09513_);
  not _33221_ (_10107_, _10105_);
  and _33222_ (_10108_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _33223_ (_12516_, _10108_, _10106_);
  and _33224_ (_10109_, _10105_, _09520_);
  and _33225_ (_10110_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _33226_ (_12517_, _10110_, _10109_);
  and _33227_ (_10111_, _10105_, _09523_);
  and _33228_ (_10112_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _33229_ (_12518_, _10112_, _10111_);
  and _33230_ (_10113_, _10105_, _09526_);
  and _33231_ (_10114_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _33232_ (_12519_, _10114_, _10113_);
  and _33233_ (_10115_, _10105_, _09529_);
  and _33234_ (_10116_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _33235_ (_12520_, _10116_, _10115_);
  and _33236_ (_10117_, _10105_, _09532_);
  and _33237_ (_10118_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _33238_ (_12522_, _10118_, _10117_);
  and _33239_ (_10119_, _10105_, _09535_);
  and _33240_ (_10120_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _33241_ (_12523_, _10120_, _10119_);
  and _33242_ (_10121_, _10105_, _09538_);
  and _33243_ (_10122_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _33244_ (_12524_, _10122_, _10121_);
  and _33245_ (_10123_, _10104_, _09515_);
  and _33246_ (_10124_, _10123_, _09513_);
  not _33247_ (_10125_, _10123_);
  and _33248_ (_10126_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or _33249_ (_12525_, _10126_, _10124_);
  and _33250_ (_10127_, _10123_, _09520_);
  and _33251_ (_10128_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or _33252_ (_12527_, _10128_, _10127_);
  and _33253_ (_10129_, _10123_, _09523_);
  and _33254_ (_10130_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or _33255_ (_12528_, _10130_, _10129_);
  and _33256_ (_10131_, _10123_, _09526_);
  and _33257_ (_10132_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or _33258_ (_12529_, _10132_, _10131_);
  and _33259_ (_10133_, _10123_, _09529_);
  and _33260_ (_10134_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or _33261_ (_12530_, _10134_, _10133_);
  and _33262_ (_10135_, _10123_, _09532_);
  and _33263_ (_10136_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or _33264_ (_12531_, _10136_, _10135_);
  and _33265_ (_10137_, _10123_, _09535_);
  and _33266_ (_10138_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or _33267_ (_12532_, _10138_, _10137_);
  and _33268_ (_10139_, _10123_, _09538_);
  and _33269_ (_10140_, _10125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or _33270_ (_12533_, _10140_, _10139_);
  and _33271_ (_10141_, _10104_, _09542_);
  and _33272_ (_10142_, _10141_, _09513_);
  not _33273_ (_10143_, _10141_);
  and _33274_ (_10144_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or _33275_ (_12535_, _10144_, _10142_);
  and _33276_ (_10145_, _10141_, _09520_);
  and _33277_ (_10146_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or _33278_ (_12536_, _10146_, _10145_);
  and _33279_ (_10147_, _10141_, _09523_);
  and _33280_ (_10148_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or _33281_ (_12537_, _10148_, _10147_);
  and _33282_ (_10149_, _10141_, _09526_);
  and _33283_ (_10150_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or _33284_ (_12539_, _10150_, _10149_);
  and _33285_ (_10151_, _10141_, _09529_);
  and _33286_ (_10152_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or _33287_ (_12540_, _10152_, _10151_);
  and _33288_ (_10153_, _10141_, _09532_);
  and _33289_ (_10154_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or _33290_ (_12541_, _10154_, _10153_);
  and _33291_ (_10155_, _10141_, _09535_);
  and _33292_ (_10156_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or _33293_ (_12542_, _10156_, _10155_);
  and _33294_ (_10157_, _10141_, _09538_);
  and _33295_ (_10158_, _10143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or _33296_ (_12543_, _10158_, _10157_);
  and _33297_ (_10159_, _10104_, _09562_);
  and _33298_ (_10160_, _10159_, _09513_);
  not _33299_ (_10161_, _10159_);
  and _33300_ (_10162_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _33301_ (_12544_, _10162_, _10160_);
  and _33302_ (_10163_, _10159_, _09520_);
  and _33303_ (_10164_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _33304_ (_12546_, _10164_, _10163_);
  and _33305_ (_10165_, _10159_, _09523_);
  and _33306_ (_10166_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _33307_ (_12547_, _10166_, _10165_);
  and _33308_ (_10167_, _10159_, _09526_);
  and _33309_ (_10168_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _33310_ (_12548_, _10168_, _10167_);
  and _33311_ (_10169_, _10159_, _09529_);
  and _33312_ (_10170_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _33313_ (_12549_, _10170_, _10169_);
  and _33314_ (_10171_, _10159_, _09532_);
  and _33315_ (_10172_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _33316_ (_12551_, _10172_, _10171_);
  and _33317_ (_10173_, _10159_, _09535_);
  and _33318_ (_10174_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _33319_ (_12552_, _10174_, _10173_);
  and _33320_ (_10175_, _10159_, _09538_);
  and _33321_ (_10176_, _10161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _33322_ (_12553_, _10176_, _10175_);
  and _33323_ (_10177_, _10104_, _09582_);
  and _33324_ (_10178_, _10177_, _09513_);
  not _33325_ (_10179_, _10177_);
  and _33326_ (_10180_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _33327_ (_12554_, _10180_, _10178_);
  and _33328_ (_10181_, _10177_, _09520_);
  and _33329_ (_10182_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _33330_ (_12555_, _10182_, _10181_);
  and _33331_ (_10183_, _10177_, _09523_);
  and _33332_ (_10184_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _33333_ (_12556_, _10184_, _10183_);
  and _33334_ (_10185_, _10177_, _09526_);
  and _33335_ (_10186_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _33336_ (_12558_, _10186_, _10185_);
  and _33337_ (_10187_, _10177_, _09529_);
  and _33338_ (_10188_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _33339_ (_12559_, _10188_, _10187_);
  and _33340_ (_10189_, _10177_, _09532_);
  and _33341_ (_10190_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _33342_ (_12560_, _10190_, _10189_);
  and _33343_ (_10191_, _10177_, _09535_);
  and _33344_ (_10192_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _33345_ (_12561_, _10192_, _10191_);
  and _33346_ (_10193_, _10177_, _09538_);
  and _33347_ (_10194_, _10179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _33348_ (_12563_, _10194_, _10193_);
  and _33349_ (_10195_, _10104_, _09601_);
  and _33350_ (_10196_, _10195_, _09513_);
  not _33351_ (_10197_, _10195_);
  and _33352_ (_10198_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or _33353_ (_12564_, _10198_, _10196_);
  and _33354_ (_10199_, _10195_, _09520_);
  and _33355_ (_10200_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or _33356_ (_12565_, _10200_, _10199_);
  and _33357_ (_10201_, _10195_, _09523_);
  and _33358_ (_10202_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or _33359_ (_12566_, _10202_, _10201_);
  and _33360_ (_10203_, _10195_, _09526_);
  and _33361_ (_10204_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or _33362_ (_12567_, _10204_, _10203_);
  and _33363_ (_10205_, _10195_, _09529_);
  and _33364_ (_10206_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or _33365_ (_12568_, _10206_, _10205_);
  and _33366_ (_10207_, _10195_, _09532_);
  and _33367_ (_10208_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or _33368_ (_12570_, _10208_, _10207_);
  and _33369_ (_10209_, _10195_, _09535_);
  and _33370_ (_10210_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or _33371_ (_12571_, _10210_, _10209_);
  and _33372_ (_10211_, _10195_, _09538_);
  and _33373_ (_10212_, _10197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or _33374_ (_12572_, _10212_, _10211_);
  and _33375_ (_10213_, _10104_, _09620_);
  and _33376_ (_10214_, _10213_, _09513_);
  not _33377_ (_10215_, _10213_);
  and _33378_ (_10216_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or _33379_ (_12573_, _10216_, _10214_);
  and _33380_ (_10217_, _10213_, _09520_);
  and _33381_ (_10218_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or _33382_ (_12575_, _10218_, _10217_);
  and _33383_ (_10219_, _10213_, _09523_);
  and _33384_ (_10220_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or _33385_ (_12576_, _10220_, _10219_);
  and _33386_ (_10221_, _10213_, _09526_);
  and _33387_ (_10222_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or _33388_ (_12577_, _10222_, _10221_);
  and _33389_ (_10223_, _10213_, _09529_);
  and _33390_ (_10224_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or _33391_ (_12578_, _10224_, _10223_);
  and _33392_ (_10225_, _10213_, _09532_);
  and _33393_ (_10226_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or _33394_ (_12579_, _10226_, _10225_);
  and _33395_ (_10227_, _10213_, _09535_);
  and _33396_ (_10228_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or _33397_ (_12580_, _10228_, _10227_);
  and _33398_ (_10229_, _10213_, _09538_);
  and _33399_ (_10230_, _10215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or _33400_ (_12581_, _10230_, _10229_);
  and _33401_ (_10231_, _10104_, _09639_);
  and _33402_ (_10232_, _10231_, _09513_);
  not _33403_ (_10233_, _10231_);
  and _33404_ (_10234_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _33405_ (_12583_, _10234_, _10232_);
  and _33406_ (_10235_, _10231_, _09520_);
  and _33407_ (_10236_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _33408_ (_12584_, _10236_, _10235_);
  and _33409_ (_10237_, _10231_, _09523_);
  and _33410_ (_10238_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _33411_ (_12585_, _10238_, _10237_);
  and _33412_ (_10239_, _10231_, _09526_);
  and _33413_ (_10240_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _33414_ (_12587_, _10240_, _10239_);
  and _33415_ (_10241_, _10231_, _09529_);
  and _33416_ (_10242_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _33417_ (_12588_, _10242_, _10241_);
  and _33418_ (_10243_, _10231_, _09532_);
  and _33419_ (_10244_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _33420_ (_12589_, _10244_, _10243_);
  and _33421_ (_10245_, _10231_, _09535_);
  and _33422_ (_10246_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _33423_ (_12590_, _10246_, _10245_);
  and _33424_ (_10247_, _10231_, _09538_);
  and _33425_ (_10248_, _10233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _33426_ (_12591_, _10248_, _10247_);
  and _33427_ (_10249_, _10104_, _09659_);
  and _33428_ (_10250_, _10249_, _09513_);
  not _33429_ (_10251_, _10249_);
  and _33430_ (_10252_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or _33431_ (_12592_, _10252_, _10250_);
  and _33432_ (_10253_, _10249_, _09520_);
  and _33433_ (_10254_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or _33434_ (_12594_, _10254_, _10253_);
  and _33435_ (_10255_, _10249_, _09523_);
  and _33436_ (_10256_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or _33437_ (_12595_, _10256_, _10255_);
  and _33438_ (_10257_, _10249_, _09526_);
  and _33439_ (_10258_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or _33440_ (_12596_, _10258_, _10257_);
  and _33441_ (_10259_, _10249_, _09529_);
  and _33442_ (_10260_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or _33443_ (_12597_, _10260_, _10259_);
  and _33444_ (_10261_, _10249_, _09532_);
  and _33445_ (_10262_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or _33446_ (_12599_, _10262_, _10261_);
  and _33447_ (_10263_, _10249_, _09535_);
  and _33448_ (_10264_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or _33449_ (_12600_, _10264_, _10263_);
  and _33450_ (_10265_, _10249_, _09538_);
  and _33451_ (_10266_, _10251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or _33452_ (_12601_, _10266_, _10265_);
  and _33453_ (_10267_, _10104_, _09678_);
  and _33454_ (_10268_, _10267_, _09513_);
  not _33455_ (_10269_, _10267_);
  and _33456_ (_10270_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _33457_ (_12602_, _10270_, _10268_);
  and _33458_ (_10271_, _10267_, _09520_);
  and _33459_ (_10272_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _33460_ (_12603_, _10272_, _10271_);
  and _33461_ (_10273_, _10267_, _09523_);
  and _33462_ (_10274_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _33463_ (_12604_, _10274_, _10273_);
  and _33464_ (_10275_, _10267_, _09526_);
  and _33465_ (_10276_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _33466_ (_12606_, _10276_, _10275_);
  and _33467_ (_10277_, _10267_, _09529_);
  and _33468_ (_10278_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _33469_ (_12607_, _10278_, _10277_);
  and _33470_ (_10279_, _10267_, _09532_);
  and _33471_ (_10280_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _33472_ (_12608_, _10280_, _10279_);
  and _33473_ (_10281_, _10267_, _09535_);
  and _33474_ (_10282_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _33475_ (_12609_, _10282_, _10281_);
  and _33476_ (_10283_, _10267_, _09538_);
  and _33477_ (_10284_, _10269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _33478_ (_12611_, _10284_, _10283_);
  and _33479_ (_10285_, _10104_, _09697_);
  and _33480_ (_10286_, _10285_, _09513_);
  not _33481_ (_10287_, _10285_);
  and _33482_ (_10288_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _33483_ (_12612_, _10288_, _10286_);
  and _33484_ (_10289_, _10285_, _09520_);
  and _33485_ (_10290_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _33486_ (_12613_, _10290_, _10289_);
  and _33487_ (_10291_, _10285_, _09523_);
  and _33488_ (_10292_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _33489_ (_12615_, _10292_, _10291_);
  and _33490_ (_10293_, _10285_, _09526_);
  and _33491_ (_10294_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _33492_ (_12616_, _10294_, _10293_);
  and _33493_ (_10295_, _10285_, _09529_);
  and _33494_ (_10296_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _33495_ (_12617_, _10296_, _10295_);
  and _33496_ (_10297_, _10285_, _09532_);
  and _33497_ (_10298_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _33498_ (_12619_, _10298_, _10297_);
  and _33499_ (_10299_, _10285_, _09535_);
  and _33500_ (_10300_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _33501_ (_12620_, _10300_, _10299_);
  and _33502_ (_10301_, _10285_, _09538_);
  and _33503_ (_10302_, _10287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _33504_ (_12621_, _10302_, _10301_);
  and _33505_ (_10303_, _10104_, _09716_);
  and _33506_ (_10304_, _10303_, _09513_);
  not _33507_ (_10305_, _10303_);
  and _33508_ (_10306_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or _33509_ (_12622_, _10306_, _10304_);
  and _33510_ (_10307_, _10303_, _09520_);
  and _33511_ (_10308_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or _33512_ (_12623_, _10308_, _10307_);
  and _33513_ (_10309_, _10303_, _09523_);
  and _33514_ (_10310_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or _33515_ (_12624_, _10310_, _10309_);
  and _33516_ (_10311_, _10303_, _09526_);
  and _33517_ (_10312_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or _33518_ (_12625_, _10312_, _10311_);
  and _33519_ (_10313_, _10303_, _09529_);
  and _33520_ (_10314_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or _33521_ (_12627_, _10314_, _10313_);
  and _33522_ (_10315_, _10303_, _09532_);
  and _33523_ (_10316_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or _33524_ (_12628_, _10316_, _10315_);
  and _33525_ (_10317_, _10303_, _09535_);
  and _33526_ (_10318_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or _33527_ (_12629_, _10318_, _10317_);
  and _33528_ (_10319_, _10303_, _09538_);
  and _33529_ (_10320_, _10305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or _33530_ (_12630_, _10320_, _10319_);
  and _33531_ (_10321_, _10104_, _09736_);
  and _33532_ (_10322_, _10321_, _09513_);
  not _33533_ (_10323_, _10321_);
  and _33534_ (_10324_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or _33535_ (_12632_, _10324_, _10322_);
  and _33536_ (_10325_, _10321_, _09520_);
  and _33537_ (_10326_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or _33538_ (_12633_, _10326_, _10325_);
  and _33539_ (_10327_, _10321_, _09523_);
  and _33540_ (_10328_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or _33541_ (_12634_, _10328_, _10327_);
  and _33542_ (_10329_, _10321_, _09526_);
  and _33543_ (_10330_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or _33544_ (_12635_, _10330_, _10329_);
  and _33545_ (_10331_, _10321_, _09529_);
  and _33546_ (_10332_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or _33547_ (_12636_, _10332_, _10331_);
  and _33548_ (_10333_, _10321_, _09532_);
  and _33549_ (_10334_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or _33550_ (_12637_, _10334_, _10333_);
  and _33551_ (_10335_, _10321_, _09535_);
  and _33552_ (_10336_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or _33553_ (_12639_, _10336_, _10335_);
  and _33554_ (_10337_, _10321_, _09538_);
  and _33555_ (_10338_, _10323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or _33556_ (_12640_, _10338_, _10337_);
  and _33557_ (_10339_, _10104_, _09755_);
  and _33558_ (_10340_, _10339_, _09513_);
  not _33559_ (_10341_, _10339_);
  and _33560_ (_10342_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _33561_ (_12641_, _10342_, _10340_);
  and _33562_ (_10343_, _10339_, _09520_);
  and _33563_ (_10344_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _33564_ (_12643_, _10344_, _10343_);
  and _33565_ (_10345_, _10339_, _09523_);
  and _33566_ (_10346_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _33567_ (_12644_, _10346_, _10345_);
  and _33568_ (_10347_, _10339_, _09526_);
  and _33569_ (_10348_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _33570_ (_12645_, _10348_, _10347_);
  and _33571_ (_10349_, _10339_, _09529_);
  and _33572_ (_10350_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _33573_ (_12646_, _10350_, _10349_);
  and _33574_ (_10351_, _10339_, _09532_);
  and _33575_ (_10352_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _33576_ (_12647_, _10352_, _10351_);
  and _33577_ (_10353_, _10339_, _09535_);
  and _33578_ (_10354_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _33579_ (_12648_, _10354_, _10353_);
  and _33580_ (_10355_, _10339_, _09538_);
  and _33581_ (_10356_, _10341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _33582_ (_12649_, _10356_, _10355_);
  and _33583_ (_10357_, _10104_, _09774_);
  and _33584_ (_10358_, _10357_, _09513_);
  not _33585_ (_10359_, _10357_);
  and _33586_ (_10360_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _33587_ (_12651_, _10360_, _10358_);
  and _33588_ (_10361_, _10357_, _09520_);
  and _33589_ (_10362_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _33590_ (_12652_, _10362_, _10361_);
  and _33591_ (_10363_, _10357_, _09523_);
  and _33592_ (_10364_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _33593_ (_12653_, _10364_, _10363_);
  and _33594_ (_10365_, _10357_, _09526_);
  and _33595_ (_10366_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _33596_ (_12655_, _10366_, _10365_);
  and _33597_ (_10367_, _10357_, _09529_);
  and _33598_ (_10368_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _33599_ (_12656_, _10368_, _10367_);
  and _33600_ (_10369_, _10357_, _09532_);
  and _33601_ (_10370_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _33602_ (_12657_, _10370_, _10369_);
  and _33603_ (_10371_, _10357_, _09535_);
  and _33604_ (_10372_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _33605_ (_12658_, _10372_, _10371_);
  and _33606_ (_10373_, _10357_, _09538_);
  and _33607_ (_10374_, _10359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _33608_ (_12659_, _10374_, _10373_);
  and _33609_ (_10375_, _10104_, _09793_);
  and _33610_ (_10376_, _10375_, _09513_);
  not _33611_ (_10377_, _10375_);
  and _33612_ (_10378_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or _33613_ (_12660_, _10378_, _10376_);
  and _33614_ (_10379_, _10375_, _09520_);
  and _33615_ (_10380_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or _33616_ (_12661_, _10380_, _10379_);
  and _33617_ (_10381_, _10375_, _09523_);
  and _33618_ (_10382_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or _33619_ (_12663_, _10382_, _10381_);
  and _33620_ (_10383_, _10375_, _09526_);
  and _33621_ (_10384_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or _33622_ (_12664_, _10384_, _10383_);
  and _33623_ (_10385_, _10375_, _09529_);
  and _33624_ (_10386_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or _33625_ (_12665_, _10386_, _10385_);
  and _33626_ (_10387_, _10375_, _09532_);
  and _33627_ (_10388_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or _33628_ (_12667_, _10388_, _10387_);
  and _33629_ (_10389_, _10375_, _09535_);
  and _33630_ (_10390_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or _33631_ (_12668_, _10390_, _10389_);
  and _33632_ (_10391_, _10375_, _09538_);
  and _33633_ (_10392_, _10377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or _33634_ (_12669_, _10392_, _10391_);
  and _33635_ (_10393_, _09252_, _05824_);
  and _33636_ (_10394_, _10393_, _09812_);
  and _33637_ (_10395_, _10394_, _09265_);
  and _33638_ (_10396_, _10395_, _09513_);
  not _33639_ (_10397_, _10395_);
  and _33640_ (_10398_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or _33641_ (_12670_, _10398_, _10396_);
  and _33642_ (_10399_, _10395_, _09520_);
  and _33643_ (_10400_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  or _33644_ (_12671_, _10400_, _10399_);
  and _33645_ (_10401_, _10395_, _09523_);
  and _33646_ (_10402_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or _33647_ (_12672_, _10402_, _10401_);
  and _33648_ (_10403_, _10395_, _09526_);
  and _33649_ (_10404_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  or _33650_ (_12674_, _10404_, _10403_);
  and _33651_ (_10405_, _10395_, _09529_);
  and _33652_ (_10406_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or _33653_ (_12675_, _10406_, _10405_);
  and _33654_ (_10407_, _10395_, _09532_);
  and _33655_ (_10408_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or _33656_ (_12676_, _10408_, _10407_);
  and _33657_ (_10409_, _10395_, _09535_);
  and _33658_ (_10410_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  or _33659_ (_12677_, _10410_, _10409_);
  and _33660_ (_10411_, _10395_, _09538_);
  and _33661_ (_10412_, _10397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  or _33662_ (_12679_, _10412_, _10411_);
  and _33663_ (_10413_, _10394_, _09515_);
  and _33664_ (_10414_, _10413_, _09513_);
  not _33665_ (_10415_, _10413_);
  and _33666_ (_10416_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _33667_ (_12680_, _10416_, _10414_);
  and _33668_ (_10417_, _10413_, _09520_);
  and _33669_ (_10418_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _33670_ (_12681_, _10418_, _10417_);
  and _33671_ (_10419_, _10413_, _09523_);
  and _33672_ (_10420_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _33673_ (_12682_, _10420_, _10419_);
  and _33674_ (_10421_, _10413_, _09526_);
  and _33675_ (_10422_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _33676_ (_12683_, _10422_, _10421_);
  and _33677_ (_10423_, _10413_, _09529_);
  and _33678_ (_10424_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _33679_ (_12684_, _10424_, _10423_);
  and _33680_ (_10425_, _10413_, _09532_);
  and _33681_ (_10426_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _33682_ (_12686_, _10426_, _10425_);
  and _33683_ (_10427_, _10413_, _09535_);
  and _33684_ (_10428_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _33685_ (_12687_, _10428_, _10427_);
  and _33686_ (_10429_, _10413_, _09538_);
  and _33687_ (_10430_, _10415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _33688_ (_12688_, _10430_, _10429_);
  and _33689_ (_10431_, _10394_, _09542_);
  and _33690_ (_10432_, _10431_, _09513_);
  not _33691_ (_10433_, _10431_);
  and _33692_ (_10434_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _33693_ (_12689_, _10434_, _10432_);
  and _33694_ (_10435_, _10431_, _09520_);
  and _33695_ (_10436_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _33696_ (_12691_, _10436_, _10435_);
  and _33697_ (_10437_, _10431_, _09523_);
  and _33698_ (_10438_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _33699_ (_12692_, _10438_, _10437_);
  and _33700_ (_10439_, _10431_, _09526_);
  and _33701_ (_10440_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _33702_ (_12693_, _10440_, _10439_);
  and _33703_ (_10441_, _10431_, _09529_);
  and _33704_ (_10442_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _33705_ (_12694_, _10442_, _10441_);
  and _33706_ (_10443_, _10431_, _09532_);
  and _33707_ (_10444_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _33708_ (_12695_, _10444_, _10443_);
  and _33709_ (_10445_, _10431_, _09535_);
  and _33710_ (_10446_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _33711_ (_12696_, _10446_, _10445_);
  and _33712_ (_10447_, _10431_, _09538_);
  and _33713_ (_10448_, _10433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _33714_ (_12697_, _10448_, _10447_);
  and _33715_ (_10449_, _10394_, _09562_);
  and _33716_ (_10450_, _10449_, _09513_);
  not _33717_ (_10451_, _10449_);
  and _33718_ (_10452_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or _33719_ (_12699_, _10452_, _10450_);
  and _33720_ (_10453_, _10449_, _09520_);
  and _33721_ (_10454_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or _33722_ (_12700_, _10454_, _10453_);
  and _33723_ (_10455_, _10449_, _09523_);
  and _33724_ (_10456_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or _33725_ (_12701_, _10456_, _10455_);
  and _33726_ (_10457_, _10449_, _09526_);
  and _33727_ (_10458_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or _33728_ (_12703_, _10458_, _10457_);
  and _33729_ (_10459_, _10449_, _09529_);
  and _33730_ (_10460_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or _33731_ (_12704_, _10460_, _10459_);
  and _33732_ (_10461_, _10449_, _09532_);
  and _33733_ (_10462_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or _33734_ (_12705_, _10462_, _10461_);
  and _33735_ (_10463_, _10449_, _09535_);
  and _33736_ (_10464_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or _33737_ (_12706_, _10464_, _10463_);
  and _33738_ (_10465_, _10449_, _09538_);
  and _33739_ (_10466_, _10451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or _33740_ (_12707_, _10466_, _10465_);
  and _33741_ (_10467_, _10394_, _09582_);
  and _33742_ (_10468_, _10467_, _09513_);
  not _33743_ (_10469_, _10467_);
  and _33744_ (_10470_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or _33745_ (_12708_, _10470_, _10468_);
  and _33746_ (_10471_, _10467_, _09520_);
  and _33747_ (_10472_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or _33748_ (_12710_, _10472_, _10471_);
  and _33749_ (_10473_, _10467_, _09523_);
  and _33750_ (_10474_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or _33751_ (_12711_, _10474_, _10473_);
  and _33752_ (_10475_, _10467_, _09526_);
  and _33753_ (_10476_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or _33754_ (_12712_, _10476_, _10475_);
  and _33755_ (_10477_, _10467_, _09529_);
  and _33756_ (_10478_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or _33757_ (_12713_, _10478_, _10477_);
  and _33758_ (_10479_, _10467_, _09532_);
  and _33759_ (_10480_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or _33760_ (_12715_, _10480_, _10479_);
  and _33761_ (_10481_, _10467_, _09535_);
  and _33762_ (_10482_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or _33763_ (_12716_, _10482_, _10481_);
  and _33764_ (_10483_, _10467_, _09538_);
  and _33765_ (_10484_, _10469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or _33766_ (_12717_, _10484_, _10483_);
  and _33767_ (_10485_, _10394_, _09601_);
  and _33768_ (_10486_, _10485_, _09513_);
  not _33769_ (_10487_, _10485_);
  and _33770_ (_10488_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _33771_ (_12719_, _10488_, _10486_);
  and _33772_ (_10489_, _10485_, _09520_);
  and _33773_ (_10490_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _33774_ (_12720_, _10490_, _10489_);
  and _33775_ (_10491_, _10485_, _09523_);
  and _33776_ (_10492_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _33777_ (_12721_, _10492_, _10491_);
  and _33778_ (_10493_, _10485_, _09526_);
  and _33779_ (_10494_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _33780_ (_12723_, _10494_, _10493_);
  and _33781_ (_10495_, _10485_, _09529_);
  and _33782_ (_10496_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _33783_ (_12724_, _10496_, _10495_);
  and _33784_ (_10497_, _10485_, _09532_);
  and _33785_ (_10498_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _33786_ (_12725_, _10498_, _10497_);
  and _33787_ (_10499_, _10485_, _09535_);
  and _33788_ (_10500_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _33789_ (_12726_, _10500_, _10499_);
  and _33790_ (_10501_, _10485_, _09538_);
  and _33791_ (_10502_, _10487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _33792_ (_12727_, _10502_, _10501_);
  and _33793_ (_10503_, _10394_, _09620_);
  and _33794_ (_10504_, _10503_, _09513_);
  not _33795_ (_10505_, _10503_);
  and _33796_ (_10506_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _33797_ (_12728_, _10506_, _10504_);
  and _33798_ (_10507_, _10503_, _09520_);
  and _33799_ (_10508_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _33800_ (_12729_, _10508_, _10507_);
  and _33801_ (_10509_, _10503_, _09523_);
  and _33802_ (_10510_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _33803_ (_12731_, _10510_, _10509_);
  and _33804_ (_10511_, _10503_, _09526_);
  and _33805_ (_10512_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _33806_ (_12732_, _10512_, _10511_);
  and _33807_ (_10513_, _10503_, _09529_);
  and _33808_ (_10514_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _33809_ (_12733_, _10514_, _10513_);
  and _33810_ (_10515_, _10503_, _09532_);
  and _33811_ (_10516_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _33812_ (_12735_, _10516_, _10515_);
  and _33813_ (_10517_, _10503_, _09535_);
  and _33814_ (_10518_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _33815_ (_12736_, _10518_, _10517_);
  and _33816_ (_10519_, _10503_, _09538_);
  and _33817_ (_10520_, _10505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _33818_ (_12737_, _10520_, _10519_);
  and _33819_ (_10521_, _10394_, _09639_);
  and _33820_ (_10522_, _10521_, _09513_);
  not _33821_ (_10523_, _10521_);
  and _33822_ (_10524_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or _33823_ (_12738_, _10524_, _10522_);
  and _33824_ (_10525_, _10521_, _09520_);
  and _33825_ (_10526_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or _33826_ (_12739_, _10526_, _10525_);
  and _33827_ (_10527_, _10521_, _09523_);
  and _33828_ (_10528_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or _33829_ (_12740_, _10528_, _10527_);
  and _33830_ (_10529_, _10521_, _09526_);
  and _33831_ (_10530_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or _33832_ (_12741_, _10530_, _10529_);
  and _33833_ (_10531_, _10521_, _09529_);
  and _33834_ (_10532_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or _33835_ (_12743_, _10532_, _10531_);
  and _33836_ (_10533_, _10521_, _09532_);
  and _33837_ (_10534_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or _33838_ (_12744_, _10534_, _10533_);
  and _33839_ (_10535_, _10521_, _09535_);
  and _33840_ (_10536_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or _33841_ (_12745_, _10536_, _10535_);
  and _33842_ (_10537_, _10521_, _09538_);
  and _33843_ (_10538_, _10523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or _33844_ (_12746_, _10538_, _10537_);
  and _33845_ (_10539_, _10394_, _09659_);
  and _33846_ (_10540_, _10539_, _09513_);
  not _33847_ (_10541_, _10539_);
  and _33848_ (_10542_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _33849_ (_12748_, _10542_, _10540_);
  and _33850_ (_10543_, _10539_, _09520_);
  and _33851_ (_10544_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _33852_ (_12749_, _10544_, _10543_);
  and _33853_ (_10545_, _10539_, _09523_);
  and _33854_ (_10546_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _33855_ (_12750_, _10546_, _10545_);
  and _33856_ (_10547_, _10539_, _09526_);
  and _33857_ (_10548_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _33858_ (_12751_, _10548_, _10547_);
  and _33859_ (_10549_, _10539_, _09529_);
  and _33860_ (_10550_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _33861_ (_12752_, _10550_, _10549_);
  and _33862_ (_10551_, _10539_, _09532_);
  and _33863_ (_10552_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _33864_ (_12753_, _10552_, _10551_);
  and _33865_ (_10553_, _10539_, _09535_);
  and _33866_ (_10554_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _33867_ (_12755_, _10554_, _10553_);
  and _33868_ (_10555_, _10539_, _09538_);
  and _33869_ (_10556_, _10541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _33870_ (_12756_, _10556_, _10555_);
  and _33871_ (_10557_, _10394_, _09678_);
  and _33872_ (_10558_, _10557_, _09513_);
  not _33873_ (_10559_, _10557_);
  and _33874_ (_10560_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or _33875_ (_12757_, _10560_, _10558_);
  and _33876_ (_10561_, _10557_, _09520_);
  and _33877_ (_10562_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or _33878_ (_12759_, _10562_, _10561_);
  and _33879_ (_10563_, _10557_, _09523_);
  and _33880_ (_10564_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or _33881_ (_12760_, _10564_, _10563_);
  and _33882_ (_10565_, _10557_, _09526_);
  and _33883_ (_10566_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or _33884_ (_12761_, _10566_, _10565_);
  and _33885_ (_10567_, _10557_, _09529_);
  and _33886_ (_10568_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or _33887_ (_12762_, _10568_, _10567_);
  and _33888_ (_10569_, _10557_, _09532_);
  and _33889_ (_10570_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or _33890_ (_12763_, _10570_, _10569_);
  and _33891_ (_10571_, _10557_, _09535_);
  and _33892_ (_10572_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or _33893_ (_12764_, _10572_, _10571_);
  and _33894_ (_10573_, _10557_, _09538_);
  and _33895_ (_10574_, _10559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or _33896_ (_12765_, _10574_, _10573_);
  and _33897_ (_10575_, _10394_, _09697_);
  and _33898_ (_10576_, _10575_, _09513_);
  not _33899_ (_10577_, _10575_);
  and _33900_ (_10578_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or _33901_ (_12767_, _10578_, _10576_);
  and _33902_ (_10579_, _10575_, _09520_);
  and _33903_ (_10580_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or _33904_ (_12768_, _10580_, _10579_);
  and _33905_ (_10581_, _10575_, _09523_);
  and _33906_ (_10582_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or _33907_ (_12769_, _10582_, _10581_);
  and _33908_ (_10583_, _10575_, _09526_);
  and _33909_ (_10584_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or _33910_ (_12771_, _10584_, _10583_);
  and _33911_ (_10585_, _10575_, _09529_);
  and _33912_ (_10586_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or _33913_ (_12772_, _10586_, _10585_);
  and _33914_ (_10587_, _10575_, _09532_);
  and _33915_ (_10588_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or _33916_ (_12773_, _10588_, _10587_);
  and _33917_ (_10589_, _10575_, _09535_);
  and _33918_ (_10590_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or _33919_ (_12774_, _10590_, _10589_);
  and _33920_ (_10591_, _10575_, _09538_);
  and _33921_ (_10592_, _10577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or _33922_ (_12775_, _10592_, _10591_);
  and _33923_ (_10593_, _10394_, _09716_);
  and _33924_ (_10594_, _10593_, _09513_);
  not _33925_ (_10595_, _10593_);
  and _33926_ (_10596_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _33927_ (_12776_, _10596_, _10594_);
  and _33928_ (_10597_, _10593_, _09520_);
  and _33929_ (_10598_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _33930_ (_12777_, _10598_, _10597_);
  and _33931_ (_10599_, _10593_, _09523_);
  and _33932_ (_10600_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _33933_ (_12779_, _10600_, _10599_);
  and _33934_ (_10601_, _10593_, _09526_);
  and _33935_ (_10602_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _33936_ (_12780_, _10602_, _10601_);
  and _33937_ (_10603_, _10593_, _09529_);
  and _33938_ (_10604_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _33939_ (_12781_, _10604_, _10603_);
  and _33940_ (_10605_, _10593_, _09532_);
  and _33941_ (_10606_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _33942_ (_12783_, _10606_, _10605_);
  and _33943_ (_10607_, _10593_, _09535_);
  and _33944_ (_10608_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _33945_ (_12784_, _10608_, _10607_);
  and _33946_ (_10609_, _10593_, _09538_);
  and _33947_ (_10610_, _10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _33948_ (_12785_, _10610_, _10609_);
  and _33949_ (_10611_, _10394_, _09736_);
  and _33950_ (_10612_, _10611_, _09513_);
  not _33951_ (_10613_, _10611_);
  and _33952_ (_10614_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _33953_ (_12786_, _10614_, _10612_);
  and _33954_ (_10615_, _10611_, _09520_);
  and _33955_ (_10616_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _33956_ (_12787_, _10616_, _10615_);
  and _33957_ (_10617_, _10611_, _09523_);
  and _33958_ (_10618_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _33959_ (_12788_, _10618_, _10617_);
  and _33960_ (_10619_, _10611_, _09526_);
  and _33961_ (_10620_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _33962_ (_12789_, _10620_, _10619_);
  and _33963_ (_10621_, _10611_, _09529_);
  and _33964_ (_10622_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _33965_ (_12791_, _10622_, _10621_);
  and _33966_ (_10623_, _10611_, _09532_);
  and _33967_ (_10624_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _33968_ (_12792_, _10624_, _10623_);
  and _33969_ (_10625_, _10611_, _09535_);
  and _33970_ (_10626_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _33971_ (_12793_, _10626_, _10625_);
  and _33972_ (_10627_, _10611_, _09538_);
  and _33973_ (_10628_, _10613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _33974_ (_12794_, _10628_, _10627_);
  and _33975_ (_10629_, _10394_, _09755_);
  and _33976_ (_10630_, _10629_, _09513_);
  not _33977_ (_10631_, _10629_);
  and _33978_ (_10632_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or _33979_ (_12796_, _10632_, _10630_);
  and _33980_ (_10633_, _10629_, _09520_);
  and _33981_ (_10634_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or _33982_ (_12797_, _10634_, _10633_);
  and _33983_ (_10635_, _10629_, _09523_);
  and _33984_ (_10636_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or _33985_ (_12798_, _10636_, _10635_);
  and _33986_ (_10637_, _10629_, _09526_);
  and _33987_ (_10638_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or _33988_ (_12799_, _10638_, _10637_);
  and _33989_ (_10639_, _10629_, _09529_);
  and _33990_ (_10640_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or _33991_ (_12800_, _10640_, _10639_);
  and _33992_ (_10641_, _10629_, _09532_);
  and _33993_ (_10642_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or _33994_ (_12801_, _10642_, _10641_);
  and _33995_ (_10643_, _10629_, _09535_);
  and _33996_ (_10644_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or _33997_ (_12803_, _10644_, _10643_);
  and _33998_ (_10645_, _10629_, _09538_);
  and _33999_ (_10646_, _10631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or _34000_ (_12804_, _10646_, _10645_);
  and _34001_ (_10647_, _10394_, _09774_);
  and _34002_ (_10648_, _10647_, _09513_);
  not _34003_ (_10649_, _10647_);
  and _34004_ (_10650_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or _34005_ (_12805_, _10650_, _10648_);
  and _34006_ (_10651_, _10647_, _09520_);
  and _34007_ (_10652_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or _34008_ (_12807_, _10652_, _10651_);
  and _34009_ (_10653_, _10647_, _09523_);
  and _34010_ (_10654_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or _34011_ (_12808_, _10654_, _10653_);
  and _34012_ (_10655_, _10647_, _09526_);
  and _34013_ (_10656_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or _34014_ (_12809_, _10656_, _10655_);
  and _34015_ (_10657_, _10647_, _09529_);
  and _34016_ (_10658_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or _34017_ (_12810_, _10658_, _10657_);
  and _34018_ (_10659_, _10647_, _09532_);
  and _34019_ (_10660_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or _34020_ (_12811_, _10660_, _10659_);
  and _34021_ (_10661_, _10647_, _09535_);
  and _34022_ (_10662_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or _34023_ (_12812_, _10662_, _10661_);
  and _34024_ (_10663_, _10647_, _09538_);
  and _34025_ (_10664_, _10649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or _34026_ (_12813_, _10664_, _10663_);
  and _34027_ (_10665_, _10394_, _09793_);
  and _34028_ (_10666_, _10665_, _09513_);
  not _34029_ (_10667_, _10665_);
  and _34030_ (_10668_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _34031_ (_12815_, _10668_, _10666_);
  and _34032_ (_10669_, _10665_, _09520_);
  and _34033_ (_10670_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _34034_ (_12816_, _10670_, _10669_);
  and _34035_ (_10671_, _10665_, _09523_);
  and _34036_ (_10672_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _34037_ (_12817_, _10672_, _10671_);
  and _34038_ (_10673_, _10665_, _09526_);
  and _34039_ (_10674_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _34040_ (_12819_, _10674_, _10673_);
  and _34041_ (_10675_, _10665_, _09529_);
  and _34042_ (_10676_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _34043_ (_12820_, _10676_, _10675_);
  and _34044_ (_10677_, _10665_, _09532_);
  and _34045_ (_10678_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _34046_ (_12821_, _10678_, _10677_);
  and _34047_ (_10679_, _10665_, _09535_);
  and _34048_ (_10680_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _34049_ (_12822_, _10680_, _10679_);
  and _34050_ (_10681_, _10665_, _09538_);
  and _34051_ (_10682_, _10667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _34052_ (_12824_, _10682_, _10681_);
  and _34053_ (_10683_, _01187_, _00906_);
  and _34054_ (_10684_, _10683_, _05869_);
  and _34055_ (_10685_, _10684_, _09254_);
  and _34056_ (_10686_, _10685_, _09265_);
  and _34057_ (_10687_, _10686_, _09513_);
  not _34058_ (_10688_, _10686_);
  and _34059_ (_10689_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _34060_ (_12825_, _10689_, _10687_);
  and _34061_ (_10690_, _10686_, _09520_);
  and _34062_ (_10691_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or _34063_ (_12827_, _10691_, _10690_);
  and _34064_ (_10692_, _10686_, _09523_);
  and _34065_ (_10693_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or _34066_ (_12828_, _10693_, _10692_);
  and _34067_ (_10694_, _10686_, _09526_);
  and _34068_ (_10695_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or _34069_ (_12829_, _10695_, _10694_);
  and _34070_ (_10696_, _10686_, _09529_);
  and _34071_ (_10697_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or _34072_ (_12830_, _10697_, _10696_);
  and _34073_ (_10698_, _10686_, _09532_);
  and _34074_ (_10699_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _34075_ (_12831_, _10699_, _10698_);
  and _34076_ (_10700_, _10686_, _09535_);
  and _34077_ (_10701_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _34078_ (_12832_, _10701_, _10700_);
  and _34079_ (_10702_, _10686_, _09538_);
  and _34080_ (_10703_, _10688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or _34081_ (_12833_, _10703_, _10702_);
  and _34082_ (_10704_, _10685_, _09515_);
  and _34083_ (_10705_, _10704_, _09513_);
  not _34084_ (_10706_, _10704_);
  and _34085_ (_10707_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or _34086_ (_12835_, _10707_, _10705_);
  and _34087_ (_10708_, _10704_, _09520_);
  and _34088_ (_10709_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or _34089_ (_12836_, _10709_, _10708_);
  and _34090_ (_10710_, _10704_, _09523_);
  and _34091_ (_10711_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or _34092_ (_12837_, _10711_, _10710_);
  and _34093_ (_10712_, _10704_, _09526_);
  and _34094_ (_10713_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or _34095_ (_12839_, _10713_, _10712_);
  and _34096_ (_10714_, _10704_, _09529_);
  and _34097_ (_10715_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or _34098_ (_12840_, _10715_, _10714_);
  and _34099_ (_10716_, _10704_, _09532_);
  and _34100_ (_10717_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or _34101_ (_12841_, _10717_, _10716_);
  and _34102_ (_10718_, _10704_, _09535_);
  and _34103_ (_10719_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or _34104_ (_12842_, _10719_, _10718_);
  and _34105_ (_10720_, _10704_, _09538_);
  and _34106_ (_10721_, _10706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or _34107_ (_12843_, _10721_, _10720_);
  and _34108_ (_10722_, _10685_, _09542_);
  and _34109_ (_10723_, _10722_, _09513_);
  not _34110_ (_10724_, _10722_);
  and _34111_ (_10725_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or _34112_ (_12844_, _10725_, _10723_);
  and _34113_ (_10726_, _10722_, _09520_);
  and _34114_ (_10727_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or _34115_ (_12846_, _10727_, _10726_);
  and _34116_ (_10728_, _10722_, _09523_);
  and _34117_ (_10729_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or _34118_ (_12847_, _10729_, _10728_);
  and _34119_ (_10730_, _10722_, _09526_);
  and _34120_ (_10731_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or _34121_ (_12848_, _10731_, _10730_);
  and _34122_ (_10732_, _10722_, _09529_);
  and _34123_ (_10733_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or _34124_ (_12849_, _10733_, _10732_);
  and _34125_ (_10734_, _10722_, _09532_);
  and _34126_ (_10735_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or _34127_ (_12851_, _10735_, _10734_);
  and _34128_ (_10736_, _10722_, _09535_);
  and _34129_ (_10737_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or _34130_ (_12852_, _10737_, _10736_);
  and _34131_ (_10738_, _10722_, _09538_);
  and _34132_ (_10739_, _10724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or _34133_ (_12853_, _10739_, _10738_);
  and _34134_ (_10740_, _10685_, _09562_);
  and _34135_ (_10741_, _10740_, _09513_);
  not _34136_ (_10742_, _10740_);
  and _34137_ (_10743_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _34138_ (_12854_, _10743_, _10741_);
  and _34139_ (_10744_, _10740_, _09520_);
  and _34140_ (_10745_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or _34141_ (_12855_, _10745_, _10744_);
  and _34142_ (_10746_, _10740_, _09523_);
  and _34143_ (_10747_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or _34144_ (_12856_, _10747_, _10746_);
  and _34145_ (_10748_, _10740_, _09526_);
  and _34146_ (_10749_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or _34147_ (_12858_, _10749_, _10748_);
  and _34148_ (_10750_, _10740_, _09529_);
  and _34149_ (_10751_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _34150_ (_12859_, _10751_, _10750_);
  and _34151_ (_10752_, _10740_, _09532_);
  and _34152_ (_10753_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _34153_ (_12860_, _10753_, _10752_);
  and _34154_ (_10755_, _10740_, _09535_);
  and _34155_ (_10756_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _34156_ (_12861_, _10756_, _10755_);
  and _34157_ (_10757_, _10740_, _09538_);
  and _34158_ (_10758_, _10742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _34159_ (_12863_, _10758_, _10757_);
  and _34160_ (_10759_, _10685_, _09582_);
  and _34161_ (_10760_, _10759_, _09513_);
  not _34162_ (_10761_, _10759_);
  and _34163_ (_10763_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _34164_ (_12864_, _10763_, _10760_);
  and _34165_ (_10764_, _10759_, _09520_);
  and _34166_ (_10765_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or _34167_ (_12865_, _10765_, _10764_);
  and _34168_ (_10766_, _10759_, _09523_);
  and _34169_ (_10767_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or _34170_ (_12866_, _10767_, _10766_);
  and _34171_ (_10768_, _10759_, _09526_);
  and _34172_ (_10769_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or _34173_ (_12867_, _10769_, _10768_);
  and _34174_ (_10771_, _10759_, _09529_);
  and _34175_ (_10772_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or _34176_ (_12868_, _10772_, _10771_);
  and _34177_ (_10773_, _10759_, _09532_);
  and _34178_ (_10774_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _34179_ (_12870_, _10774_, _10773_);
  and _34180_ (_10775_, _10759_, _09535_);
  and _34181_ (_10776_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _34182_ (_12871_, _10776_, _10775_);
  and _34183_ (_10778_, _10759_, _09538_);
  and _34184_ (_10779_, _10761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _34185_ (_12872_, _10779_, _10778_);
  and _34186_ (_10780_, _10685_, _09601_);
  and _34187_ (_10781_, _10780_, _09513_);
  not _34188_ (_10782_, _10780_);
  and _34189_ (_10783_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or _34190_ (_12873_, _10783_, _10781_);
  and _34191_ (_10784_, _10780_, _09520_);
  and _34192_ (_10785_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or _34193_ (_12875_, _10785_, _10784_);
  and _34194_ (_10787_, _10780_, _09523_);
  and _34195_ (_10788_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or _34196_ (_12876_, _10788_, _10787_);
  and _34197_ (_10789_, _10780_, _09526_);
  and _34198_ (_10790_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or _34199_ (_12877_, _10790_, _10789_);
  and _34200_ (_10791_, _10780_, _09529_);
  and _34201_ (_10792_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or _34202_ (_12878_, _10792_, _10791_);
  and _34203_ (_10794_, _10780_, _09532_);
  and _34204_ (_10795_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or _34205_ (_12879_, _10795_, _10794_);
  and _34206_ (_10796_, _10780_, _09535_);
  and _34207_ (_10797_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or _34208_ (_12880_, _10797_, _10796_);
  and _34209_ (_10798_, _10780_, _09538_);
  and _34210_ (_10799_, _10782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or _34211_ (_12881_, _10799_, _10798_);
  and _34212_ (_10800_, _10685_, _09620_);
  and _34213_ (_10802_, _10800_, _09513_);
  not _34214_ (_10803_, _10800_);
  and _34215_ (_10804_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or _34216_ (_12883_, _10804_, _10802_);
  and _34217_ (_10805_, _10800_, _09520_);
  and _34218_ (_10806_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or _34219_ (_12884_, _10806_, _10805_);
  and _34220_ (_10807_, _10800_, _09523_);
  and _34221_ (_10808_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or _34222_ (_12885_, _10808_, _10807_);
  and _34223_ (_10809_, _10800_, _09526_);
  and _34224_ (_10810_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or _34225_ (_12887_, _10810_, _10809_);
  and _34226_ (_10811_, _10800_, _09529_);
  and _34227_ (_10812_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or _34228_ (_12888_, _10812_, _10811_);
  and _34229_ (_10813_, _10800_, _09532_);
  and _34230_ (_10814_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or _34231_ (_12889_, _10814_, _10813_);
  and _34232_ (_10815_, _10800_, _09535_);
  and _34233_ (_10816_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or _34234_ (_12890_, _10816_, _10815_);
  and _34235_ (_10817_, _10800_, _09538_);
  and _34236_ (_10818_, _10803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or _34237_ (_12891_, _10818_, _10817_);
  and _34238_ (_10819_, _10685_, _09639_);
  and _34239_ (_10820_, _10819_, _09513_);
  not _34240_ (_10821_, _10819_);
  and _34241_ (_10822_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _34242_ (_12892_, _10822_, _10820_);
  and _34243_ (_10823_, _10819_, _09520_);
  and _34244_ (_10824_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or _34245_ (_12894_, _10824_, _10823_);
  and _34246_ (_10825_, _10819_, _09523_);
  and _34247_ (_10826_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or _34248_ (_12895_, _10826_, _10825_);
  and _34249_ (_10827_, _10819_, _09526_);
  and _34250_ (_10828_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or _34251_ (_12896_, _10828_, _10827_);
  and _34252_ (_10829_, _10819_, _09529_);
  and _34253_ (_10830_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or _34254_ (_12897_, _10830_, _10829_);
  and _34255_ (_10831_, _10819_, _09532_);
  and _34256_ (_10832_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _34257_ (_12899_, _10832_, _10831_);
  and _34258_ (_10833_, _10819_, _09535_);
  and _34259_ (_10834_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _34260_ (_12900_, _10834_, _10833_);
  and _34261_ (_10835_, _10819_, _09538_);
  and _34262_ (_10836_, _10821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _34263_ (_12901_, _10836_, _10835_);
  and _34264_ (_10837_, _10685_, _09659_);
  and _34265_ (_10838_, _10837_, _09513_);
  not _34266_ (_10839_, _10837_);
  and _34267_ (_10840_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or _34268_ (_12902_, _10840_, _10838_);
  and _34269_ (_10841_, _10837_, _09520_);
  and _34270_ (_10842_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or _34271_ (_12903_, _10842_, _10841_);
  and _34272_ (_10843_, _10837_, _09523_);
  and _34273_ (_10844_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or _34274_ (_12904_, _10844_, _10843_);
  and _34275_ (_10845_, _10837_, _09526_);
  and _34276_ (_10846_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or _34277_ (_12906_, _10846_, _10845_);
  and _34278_ (_10847_, _10837_, _09529_);
  and _34279_ (_10848_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or _34280_ (_12907_, _10848_, _10847_);
  and _34281_ (_10849_, _10837_, _09532_);
  and _34282_ (_10850_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or _34283_ (_12908_, _10850_, _10849_);
  and _34284_ (_10851_, _10837_, _09535_);
  and _34285_ (_10852_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or _34286_ (_12909_, _10852_, _10851_);
  and _34287_ (_10853_, _10837_, _09538_);
  and _34288_ (_10854_, _10839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or _34289_ (_12911_, _10854_, _10853_);
  and _34290_ (_10855_, _10685_, _09678_);
  and _34291_ (_10856_, _10855_, _09513_);
  not _34292_ (_10857_, _10855_);
  and _34293_ (_10858_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _34294_ (_12912_, _10858_, _10856_);
  and _34295_ (_10859_, _10855_, _09520_);
  and _34296_ (_10860_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or _34297_ (_12913_, _10860_, _10859_);
  and _34298_ (_10861_, _10855_, _09523_);
  and _34299_ (_10862_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or _34300_ (_12914_, _10862_, _10861_);
  and _34301_ (_10863_, _10855_, _09526_);
  and _34302_ (_10864_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or _34303_ (_12915_, _10864_, _10863_);
  and _34304_ (_10865_, _10855_, _09529_);
  and _34305_ (_10866_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or _34306_ (_12916_, _10866_, _10865_);
  and _34307_ (_10867_, _10855_, _09532_);
  and _34308_ (_10868_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _34309_ (_12918_, _10868_, _10867_);
  and _34310_ (_10869_, _10855_, _09535_);
  and _34311_ (_10870_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _34312_ (_12919_, _10870_, _10869_);
  and _34313_ (_10871_, _10855_, _09538_);
  and _34314_ (_10872_, _10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or _34315_ (_12920_, _10872_, _10871_);
  and _34316_ (_10873_, _10685_, _09697_);
  and _34317_ (_10874_, _10873_, _09513_);
  not _34318_ (_10875_, _10873_);
  and _34319_ (_10876_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _34320_ (_12921_, _10876_, _10874_);
  and _34321_ (_10877_, _10873_, _09520_);
  and _34322_ (_10878_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or _34323_ (_12923_, _10878_, _10877_);
  and _34324_ (_10879_, _10873_, _09523_);
  and _34325_ (_10880_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or _34326_ (_12924_, _10880_, _10879_);
  and _34327_ (_10881_, _10873_, _09526_);
  and _34328_ (_10882_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or _34329_ (_12925_, _10882_, _10881_);
  and _34330_ (_10883_, _10873_, _09529_);
  and _34331_ (_10884_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _34332_ (_12927_, _10884_, _10883_);
  and _34333_ (_10885_, _10873_, _09532_);
  and _34334_ (_10886_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or _34335_ (_12928_, _10886_, _10885_);
  and _34336_ (_10887_, _10873_, _09535_);
  and _34337_ (_10888_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _34338_ (_12929_, _10888_, _10887_);
  and _34339_ (_10889_, _10873_, _09538_);
  and _34340_ (_10890_, _10875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _34341_ (_12930_, _10890_, _10889_);
  and _34342_ (_10891_, _10685_, _09716_);
  and _34343_ (_10892_, _10891_, _09513_);
  not _34344_ (_10893_, _10891_);
  and _34345_ (_10894_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or _34346_ (_12932_, _10894_, _10892_);
  and _34347_ (_10895_, _10891_, _09520_);
  and _34348_ (_10896_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or _34349_ (_12933_, _10896_, _10895_);
  and _34350_ (_10897_, _10891_, _09523_);
  and _34351_ (_10898_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or _34352_ (_12934_, _10898_, _10897_);
  and _34353_ (_10899_, _10891_, _09526_);
  and _34354_ (_10900_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or _34355_ (_12935_, _10900_, _10899_);
  and _34356_ (_10901_, _10891_, _09529_);
  and _34357_ (_10902_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or _34358_ (_12936_, _10902_, _10901_);
  and _34359_ (_10903_, _10891_, _09532_);
  and _34360_ (_10904_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or _34361_ (_12937_, _10904_, _10903_);
  and _34362_ (_10905_, _10891_, _09535_);
  and _34363_ (_10906_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or _34364_ (_12939_, _10906_, _10905_);
  and _34365_ (_10907_, _10891_, _09538_);
  and _34366_ (_10908_, _10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or _34367_ (_12940_, _10908_, _10907_);
  and _34368_ (_10909_, _10685_, _09736_);
  and _34369_ (_10910_, _10909_, _09513_);
  not _34370_ (_10911_, _10909_);
  and _34371_ (_10912_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or _34372_ (_12941_, _10912_, _10910_);
  and _34373_ (_10913_, _10909_, _09520_);
  and _34374_ (_10914_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or _34375_ (_12943_, _10914_, _10913_);
  and _34376_ (_10915_, _10909_, _09523_);
  and _34377_ (_10916_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or _34378_ (_12944_, _10916_, _10915_);
  and _34379_ (_10917_, _10909_, _09526_);
  and _34380_ (_10918_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or _34381_ (_12945_, _10918_, _10917_);
  and _34382_ (_10919_, _10909_, _09529_);
  and _34383_ (_10920_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or _34384_ (_12946_, _10920_, _10919_);
  and _34385_ (_10921_, _10909_, _09532_);
  and _34386_ (_10922_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or _34387_ (_12947_, _10922_, _10921_);
  and _34388_ (_10923_, _10909_, _09535_);
  and _34389_ (_10924_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or _34390_ (_12948_, _10924_, _10923_);
  and _34391_ (_10925_, _10909_, _09538_);
  and _34392_ (_10926_, _10911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or _34393_ (_12949_, _10926_, _10925_);
  and _34394_ (_10927_, _10685_, _09755_);
  and _34395_ (_10928_, _10927_, _09513_);
  not _34396_ (_10929_, _10927_);
  and _34397_ (_10930_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _34398_ (_12951_, _10930_, _10928_);
  and _34399_ (_10931_, _10927_, _09520_);
  and _34400_ (_10932_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or _34401_ (_12952_, _10932_, _10931_);
  and _34402_ (_10933_, _10927_, _09523_);
  and _34403_ (_10934_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or _34404_ (_12953_, _10934_, _10933_);
  and _34405_ (_10935_, _10927_, _09526_);
  and _34406_ (_10936_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or _34407_ (_12955_, _10936_, _10935_);
  and _34408_ (_10937_, _10927_, _09529_);
  and _34409_ (_10938_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or _34410_ (_12956_, _10938_, _10937_);
  and _34411_ (_10939_, _10927_, _09532_);
  and _34412_ (_10940_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _34413_ (_12957_, _10940_, _10939_);
  and _34414_ (_10941_, _10927_, _09535_);
  and _34415_ (_10942_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _34416_ (_12958_, _10942_, _10941_);
  and _34417_ (_10943_, _10927_, _09538_);
  and _34418_ (_10944_, _10929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or _34419_ (_12959_, _10944_, _10943_);
  and _34420_ (_10945_, _10685_, _09774_);
  and _34421_ (_10946_, _10945_, _09513_);
  not _34422_ (_10947_, _10945_);
  and _34423_ (_10948_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _34424_ (_12960_, _10948_, _10946_);
  and _34425_ (_10949_, _10945_, _09520_);
  and _34426_ (_10950_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or _34427_ (_12961_, _10950_, _10949_);
  and _34428_ (_10951_, _10945_, _09523_);
  and _34429_ (_10952_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or _34430_ (_12963_, _10952_, _10951_);
  and _34431_ (_10953_, _10945_, _09526_);
  and _34432_ (_10954_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or _34433_ (_12964_, _10954_, _10953_);
  and _34434_ (_10955_, _10945_, _09529_);
  and _34435_ (_10956_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _34436_ (_12965_, _10956_, _10955_);
  and _34437_ (_10957_, _10945_, _09532_);
  and _34438_ (_10958_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or _34439_ (_12967_, _10958_, _10957_);
  and _34440_ (_10959_, _10945_, _09535_);
  and _34441_ (_10960_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _34442_ (_12968_, _10960_, _10959_);
  and _34443_ (_10961_, _10945_, _09538_);
  and _34444_ (_10962_, _10947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _34445_ (_12969_, _10962_, _10961_);
  and _34446_ (_10963_, _10685_, _09793_);
  and _34447_ (_10964_, _10963_, _09513_);
  not _34448_ (_10965_, _10963_);
  and _34449_ (_10966_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or _34450_ (_12970_, _10966_, _10964_);
  and _34451_ (_10967_, _10963_, _09520_);
  and _34452_ (_10968_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or _34453_ (_12971_, _10968_, _10967_);
  and _34454_ (_10969_, _10963_, _09523_);
  and _34455_ (_10970_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or _34456_ (_12972_, _10970_, _10969_);
  and _34457_ (_10971_, _10963_, _09526_);
  and _34458_ (_10972_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or _34459_ (_12973_, _10972_, _10971_);
  and _34460_ (_10973_, _10963_, _09529_);
  and _34461_ (_10974_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or _34462_ (_12975_, _10974_, _10973_);
  and _34463_ (_10975_, _10963_, _09532_);
  and _34464_ (_10976_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or _34465_ (_12976_, _10976_, _10975_);
  and _34466_ (_10977_, _10963_, _09535_);
  and _34467_ (_10978_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or _34468_ (_12977_, _10978_, _10977_);
  and _34469_ (_10979_, _10963_, _09538_);
  and _34470_ (_10980_, _10965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or _34471_ (_12978_, _10980_, _10979_);
  and _34472_ (_10981_, _10684_, _09813_);
  and _34473_ (_10982_, _10981_, _09265_);
  and _34474_ (_10983_, _10982_, _09513_);
  not _34475_ (_10984_, _10982_);
  and _34476_ (_10985_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or _34477_ (_12980_, _10985_, _10983_);
  and _34478_ (_10986_, _10982_, _09520_);
  and _34479_ (_10987_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or _34480_ (_12981_, _10987_, _10986_);
  and _34481_ (_10988_, _10982_, _09523_);
  and _34482_ (_10989_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or _34483_ (_12982_, _10989_, _10988_);
  and _34484_ (_10990_, _10982_, _09526_);
  and _34485_ (_10991_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or _34486_ (_12983_, _10991_, _10990_);
  and _34487_ (_10992_, _10982_, _09529_);
  and _34488_ (_10993_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or _34489_ (_12984_, _10993_, _10992_);
  and _34490_ (_10994_, _10982_, _09532_);
  and _34491_ (_10995_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or _34492_ (_12985_, _10995_, _10994_);
  and _34493_ (_10996_, _10982_, _09535_);
  and _34494_ (_10997_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or _34495_ (_12987_, _10997_, _10996_);
  and _34496_ (_10998_, _10982_, _09538_);
  and _34497_ (_10999_, _10984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or _34498_ (_12988_, _10999_, _10998_);
  and _34499_ (_11000_, _10981_, _09515_);
  and _34500_ (_11001_, _11000_, _09513_);
  not _34501_ (_11002_, _11000_);
  and _34502_ (_11003_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _34503_ (_12989_, _11003_, _11001_);
  and _34504_ (_11004_, _11000_, _09520_);
  and _34505_ (_11005_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _34506_ (_12991_, _11005_, _11004_);
  and _34507_ (_11006_, _11000_, _09523_);
  and _34508_ (_11007_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _34509_ (_12992_, _11007_, _11006_);
  and _34510_ (_11008_, _11000_, _09526_);
  and _34511_ (_11009_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _34512_ (_12993_, _11009_, _11008_);
  and _34513_ (_11010_, _11000_, _09529_);
  and _34514_ (_11011_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _34515_ (_12994_, _11011_, _11010_);
  and _34516_ (_11012_, _11000_, _09532_);
  and _34517_ (_11013_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _34518_ (_12995_, _11013_, _11012_);
  and _34519_ (_11014_, _11000_, _09535_);
  and _34520_ (_11015_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _34521_ (_12996_, _11015_, _11014_);
  and _34522_ (_11016_, _11000_, _09538_);
  and _34523_ (_11017_, _11002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _34524_ (_12997_, _11017_, _11016_);
  and _34525_ (_11018_, _10981_, _09542_);
  and _34526_ (_11019_, _11018_, _09513_);
  not _34527_ (_11020_, _11018_);
  and _34528_ (_11021_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _34529_ (_12999_, _11021_, _11019_);
  and _34530_ (_11022_, _11018_, _09520_);
  and _34531_ (_11023_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _34532_ (_13000_, _11023_, _11022_);
  and _34533_ (_11024_, _11018_, _09523_);
  and _34534_ (_11025_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _34535_ (_13001_, _11025_, _11024_);
  and _34536_ (_11026_, _11018_, _09526_);
  and _34537_ (_11027_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _34538_ (_13003_, _11027_, _11026_);
  and _34539_ (_11028_, _11018_, _09529_);
  and _34540_ (_11029_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _34541_ (_13004_, _11029_, _11028_);
  and _34542_ (_11030_, _11018_, _09532_);
  and _34543_ (_11031_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _34544_ (_13005_, _11031_, _11030_);
  and _34545_ (_11032_, _11018_, _09535_);
  and _34546_ (_11033_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _34547_ (_13006_, _11033_, _11032_);
  and _34548_ (_11034_, _11018_, _09538_);
  and _34549_ (_11035_, _11020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _34550_ (_13007_, _11035_, _11034_);
  and _34551_ (_11036_, _10981_, _09562_);
  and _34552_ (_11037_, _11036_, _09513_);
  not _34553_ (_11038_, _11036_);
  and _34554_ (_11039_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or _34555_ (_13008_, _11039_, _11037_);
  and _34556_ (_11040_, _11036_, _09520_);
  and _34557_ (_11041_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or _34558_ (_13009_, _11041_, _11040_);
  and _34559_ (_11042_, _11036_, _09523_);
  and _34560_ (_11043_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or _34561_ (_13011_, _11043_, _11042_);
  and _34562_ (_11044_, _11036_, _09526_);
  and _34563_ (_11045_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or _34564_ (_13012_, _11045_, _11044_);
  and _34565_ (_11046_, _11036_, _09529_);
  and _34566_ (_11047_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or _34567_ (_13013_, _11047_, _11046_);
  and _34568_ (_11048_, _11036_, _09532_);
  and _34569_ (_11049_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or _34570_ (_13015_, _11049_, _11048_);
  and _34571_ (_11050_, _11036_, _09535_);
  and _34572_ (_11051_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or _34573_ (_13016_, _11051_, _11050_);
  and _34574_ (_11052_, _11036_, _09538_);
  and _34575_ (_11053_, _11038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or _34576_ (_13017_, _11053_, _11052_);
  and _34577_ (_11054_, _10981_, _09582_);
  and _34578_ (_11055_, _11054_, _09513_);
  not _34579_ (_11056_, _11054_);
  and _34580_ (_11057_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or _34581_ (_13018_, _11057_, _11055_);
  and _34582_ (_11058_, _11054_, _09520_);
  and _34583_ (_11059_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or _34584_ (_13019_, _11059_, _11058_);
  and _34585_ (_11060_, _11054_, _09523_);
  and _34586_ (_11061_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or _34587_ (_13020_, _11061_, _11060_);
  and _34588_ (_11062_, _11054_, _09526_);
  and _34589_ (_11063_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or _34590_ (_13021_, _11063_, _11062_);
  and _34591_ (_11064_, _11054_, _09529_);
  and _34592_ (_11065_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or _34593_ (_13023_, _11065_, _11064_);
  and _34594_ (_11066_, _11054_, _09532_);
  and _34595_ (_11067_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or _34596_ (_13024_, _11067_, _11066_);
  and _34597_ (_11068_, _11054_, _09535_);
  and _34598_ (_11069_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or _34599_ (_13025_, _11069_, _11068_);
  and _34600_ (_11070_, _11054_, _09538_);
  and _34601_ (_11071_, _11056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or _34602_ (_13027_, _11071_, _11070_);
  and _34603_ (_11072_, _10981_, _09601_);
  and _34604_ (_11073_, _11072_, _09513_);
  not _34605_ (_11074_, _11072_);
  and _34606_ (_11075_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _34607_ (_13028_, _11075_, _11073_);
  and _34608_ (_11076_, _11072_, _09520_);
  and _34609_ (_11077_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _34610_ (_13029_, _11077_, _11076_);
  and _34611_ (_11078_, _11072_, _09523_);
  and _34612_ (_11079_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _34613_ (_13031_, _11079_, _11078_);
  and _34614_ (_11080_, _11072_, _09526_);
  and _34615_ (_11081_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _34616_ (_13032_, _11081_, _11080_);
  and _34617_ (_11082_, _11072_, _09529_);
  and _34618_ (_11083_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _34619_ (_13033_, _11083_, _11082_);
  and _34620_ (_11084_, _11072_, _09532_);
  and _34621_ (_11085_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _34622_ (_13034_, _11085_, _11084_);
  and _34623_ (_11086_, _11072_, _09535_);
  and _34624_ (_11087_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _34625_ (_13036_, _11087_, _11086_);
  and _34626_ (_11088_, _11072_, _09538_);
  and _34627_ (_11089_, _11074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _34628_ (_13037_, _11089_, _11088_);
  and _34629_ (_11090_, _10981_, _09620_);
  and _34630_ (_11091_, _11090_, _09513_);
  not _34631_ (_11092_, _11090_);
  and _34632_ (_11093_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _34633_ (_13038_, _11093_, _11091_);
  and _34634_ (_11094_, _11090_, _09520_);
  and _34635_ (_11095_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _34636_ (_13039_, _11095_, _11094_);
  and _34637_ (_11096_, _11090_, _09523_);
  and _34638_ (_11097_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _34639_ (_13040_, _11097_, _11096_);
  and _34640_ (_11098_, _11090_, _09526_);
  and _34641_ (_11099_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _34642_ (_13041_, _11099_, _11098_);
  and _34643_ (_11100_, _11090_, _09529_);
  and _34644_ (_11101_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _34645_ (_13043_, _11101_, _11100_);
  and _34646_ (_11102_, _11090_, _09532_);
  and _34647_ (_11103_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _34648_ (_13044_, _11103_, _11102_);
  and _34649_ (_11104_, _11090_, _09535_);
  and _34650_ (_11105_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _34651_ (_13045_, _11105_, _11104_);
  and _34652_ (_11106_, _11090_, _09538_);
  and _34653_ (_11107_, _11092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _34654_ (_13046_, _11107_, _11106_);
  and _34655_ (_11108_, _10981_, _09639_);
  and _34656_ (_11109_, _11108_, _09513_);
  not _34657_ (_11110_, _11108_);
  and _34658_ (_11111_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or _34659_ (_13048_, _11111_, _11109_);
  and _34660_ (_11112_, _11108_, _09520_);
  and _34661_ (_11113_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or _34662_ (_13049_, _11113_, _11112_);
  and _34663_ (_11114_, _11108_, _09523_);
  and _34664_ (_11115_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or _34665_ (_13050_, _11115_, _11114_);
  and _34666_ (_11116_, _11108_, _09526_);
  and _34667_ (_11117_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or _34668_ (_13051_, _11117_, _11116_);
  and _34669_ (_11118_, _11108_, _09529_);
  and _34670_ (_11119_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or _34671_ (_13052_, _11119_, _11118_);
  and _34672_ (_11120_, _11108_, _09532_);
  and _34673_ (_11121_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or _34674_ (_13053_, _11121_, _11120_);
  and _34675_ (_11122_, _11108_, _09535_);
  and _34676_ (_11123_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or _34677_ (_13055_, _11123_, _11122_);
  and _34678_ (_11124_, _11108_, _09538_);
  and _34679_ (_11125_, _11110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or _34680_ (_13056_, _11125_, _11124_);
  and _34681_ (_11126_, _10981_, _09659_);
  and _34682_ (_11127_, _11126_, _09513_);
  not _34683_ (_11128_, _11126_);
  and _34684_ (_11129_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _34685_ (_13057_, _11129_, _11127_);
  and _34686_ (_11130_, _11126_, _09520_);
  and _34687_ (_11131_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _34688_ (_13058_, _11131_, _11130_);
  and _34689_ (_11132_, _11126_, _09523_);
  and _34690_ (_11133_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _34691_ (_13060_, _11133_, _11132_);
  and _34692_ (_11134_, _11126_, _09526_);
  and _34693_ (_11135_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _34694_ (_13061_, _11135_, _11134_);
  and _34695_ (_11136_, _11126_, _09529_);
  and _34696_ (_11137_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _34697_ (_13062_, _11137_, _11136_);
  and _34698_ (_11138_, _11126_, _09532_);
  and _34699_ (_11139_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _34700_ (_13063_, _11139_, _11138_);
  and _34701_ (_11140_, _11126_, _09535_);
  and _34702_ (_11141_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _34703_ (_13064_, _11141_, _11140_);
  and _34704_ (_11142_, _11126_, _09538_);
  and _34705_ (_11143_, _11128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _34706_ (_13065_, _11143_, _11142_);
  and _34707_ (_11144_, _10981_, _09678_);
  and _34708_ (_11145_, _11144_, _09513_);
  not _34709_ (_11146_, _11144_);
  and _34710_ (_11147_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or _34711_ (_13067_, _11147_, _11145_);
  and _34712_ (_11148_, _11144_, _09520_);
  and _34713_ (_11149_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or _34714_ (_13068_, _11149_, _11148_);
  and _34715_ (_11150_, _11144_, _09523_);
  and _34716_ (_11151_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or _34717_ (_13069_, _11151_, _11150_);
  and _34718_ (_11152_, _11144_, _09526_);
  and _34719_ (_11153_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or _34720_ (_13070_, _11153_, _11152_);
  and _34721_ (_11154_, _11144_, _09529_);
  and _34722_ (_11155_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or _34723_ (_13072_, _11155_, _11154_);
  and _34724_ (_11156_, _11144_, _09532_);
  and _34725_ (_11157_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or _34726_ (_13073_, _11157_, _11156_);
  and _34727_ (_11158_, _11144_, _09535_);
  and _34728_ (_11159_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or _34729_ (_13074_, _11159_, _11158_);
  and _34730_ (_11160_, _11144_, _09538_);
  and _34731_ (_11161_, _11146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or _34732_ (_13075_, _11161_, _11160_);
  and _34733_ (_11162_, _10981_, _09697_);
  and _34734_ (_11163_, _11162_, _09513_);
  not _34735_ (_11164_, _11162_);
  and _34736_ (_11165_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or _34737_ (_13076_, _11165_, _11163_);
  and _34738_ (_11166_, _11162_, _09520_);
  and _34739_ (_11167_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or _34740_ (_13077_, _11167_, _11166_);
  and _34741_ (_11168_, _11162_, _09523_);
  and _34742_ (_11169_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or _34743_ (_13079_, _11169_, _11168_);
  and _34744_ (_11170_, _11162_, _09526_);
  and _34745_ (_11171_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or _34746_ (_13080_, _11171_, _11170_);
  and _34747_ (_11172_, _11162_, _09529_);
  and _34748_ (_11173_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or _34749_ (_13081_, _11173_, _11172_);
  and _34750_ (_11174_, _11162_, _09532_);
  and _34751_ (_11175_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or _34752_ (_13082_, _11175_, _11174_);
  and _34753_ (_11176_, _11162_, _09535_);
  and _34754_ (_11177_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or _34755_ (_13084_, _11177_, _11176_);
  and _34756_ (_11178_, _11162_, _09538_);
  and _34757_ (_11179_, _11164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or _34758_ (_13085_, _11179_, _11178_);
  and _34759_ (_11180_, _10981_, _09716_);
  and _34760_ (_11181_, _11180_, _09513_);
  not _34761_ (_11182_, _11180_);
  and _34762_ (_11183_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _34763_ (_13086_, _11183_, _11181_);
  and _34764_ (_11185_, _11180_, _09520_);
  and _34765_ (_11186_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _34766_ (_13087_, _11186_, _11185_);
  and _34767_ (_11187_, _11180_, _09523_);
  and _34768_ (_11188_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _34769_ (_13088_, _11188_, _11187_);
  and _34770_ (_11189_, _11180_, _09526_);
  and _34771_ (_11190_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _34772_ (_13089_, _11190_, _11189_);
  and _34773_ (_11191_, _11180_, _09529_);
  and _34774_ (_11192_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _34775_ (_13091_, _11192_, _11191_);
  and _34776_ (_11193_, _11180_, _09532_);
  and _34777_ (_11194_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _34778_ (_13092_, _11194_, _11193_);
  and _34779_ (_11195_, _11180_, _09535_);
  and _34780_ (_11196_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _34781_ (_13093_, _11196_, _11195_);
  and _34782_ (_11197_, _11180_, _09538_);
  and _34783_ (_11199_, _11182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _34784_ (_13094_, _11199_, _11197_);
  and _34785_ (_11200_, _10981_, _09736_);
  and _34786_ (_11201_, _11200_, _09513_);
  not _34787_ (_11202_, _11200_);
  and _34788_ (_11203_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _34789_ (_13096_, _11203_, _11201_);
  and _34790_ (_11204_, _11200_, _09520_);
  and _34791_ (_11205_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _34792_ (_13097_, _11205_, _11204_);
  and _34793_ (_11206_, _11200_, _09523_);
  and _34794_ (_11207_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _34795_ (_13098_, _11207_, _11206_);
  and _34796_ (_11208_, _11200_, _09526_);
  and _34797_ (_11209_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _34798_ (_13099_, _11209_, _11208_);
  and _34799_ (_11210_, _11200_, _09529_);
  and _34800_ (_11211_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _34801_ (_13100_, _11211_, _11210_);
  and _34802_ (_11212_, _11200_, _09532_);
  and _34803_ (_11213_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _34804_ (_13101_, _11213_, _11212_);
  and _34805_ (_11214_, _11200_, _09535_);
  and _34806_ (_11215_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _34807_ (_13103_, _11215_, _11214_);
  and _34808_ (_11216_, _11200_, _09538_);
  and _34809_ (_11217_, _11202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _34810_ (_13104_, _11217_, _11216_);
  and _34811_ (_11218_, _10981_, _09755_);
  and _34812_ (_11219_, _11218_, _09513_);
  not _34813_ (_11220_, _11218_);
  and _34814_ (_11221_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or _34815_ (_13105_, _11221_, _11219_);
  and _34816_ (_11222_, _11218_, _09520_);
  and _34817_ (_11223_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or _34818_ (_13106_, _11223_, _11222_);
  and _34819_ (_11224_, _11218_, _09523_);
  and _34820_ (_11225_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or _34821_ (_13108_, _11225_, _11224_);
  and _34822_ (_11226_, _11218_, _09526_);
  and _34823_ (_11227_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or _34824_ (_13109_, _11227_, _11226_);
  and _34825_ (_11228_, _11218_, _09529_);
  and _34826_ (_11229_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or _34827_ (_13110_, _11229_, _11228_);
  and _34828_ (_11230_, _11218_, _09532_);
  and _34829_ (_11231_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or _34830_ (_13111_, _11231_, _11230_);
  and _34831_ (_11232_, _11218_, _09535_);
  and _34832_ (_11233_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or _34833_ (_13112_, _11233_, _11232_);
  and _34834_ (_11234_, _11218_, _09538_);
  and _34835_ (_11235_, _11220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or _34836_ (_13113_, _11235_, _11234_);
  and _34837_ (_11236_, _10981_, _09774_);
  and _34838_ (_11237_, _11236_, _09513_);
  not _34839_ (_11238_, _11236_);
  and _34840_ (_11239_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or _34841_ (_13115_, _11239_, _11237_);
  and _34842_ (_11240_, _11236_, _09520_);
  and _34843_ (_11241_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or _34844_ (_13116_, _11241_, _11240_);
  and _34845_ (_11242_, _11236_, _09523_);
  and _34846_ (_11243_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or _34847_ (_13117_, _11243_, _11242_);
  and _34848_ (_11244_, _11236_, _09526_);
  and _34849_ (_11245_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or _34850_ (_13118_, _11245_, _11244_);
  and _34851_ (_11246_, _11236_, _09529_);
  and _34852_ (_11247_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or _34853_ (_13120_, _11247_, _11246_);
  and _34854_ (_11248_, _11236_, _09532_);
  and _34855_ (_11249_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or _34856_ (_13121_, _11249_, _11248_);
  and _34857_ (_11250_, _11236_, _09535_);
  and _34858_ (_11251_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or _34859_ (_13122_, _11251_, _11250_);
  and _34860_ (_11252_, _11236_, _09538_);
  and _34861_ (_11253_, _11238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or _34862_ (_13123_, _11253_, _11252_);
  and _34863_ (_11254_, _10981_, _09793_);
  and _34864_ (_11255_, _11254_, _09513_);
  not _34865_ (_11256_, _11254_);
  and _34866_ (_11257_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _34867_ (_13124_, _11257_, _11255_);
  and _34868_ (_11258_, _11254_, _09520_);
  and _34869_ (_11259_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _34870_ (_13125_, _11259_, _11258_);
  and _34871_ (_11260_, _11254_, _09523_);
  and _34872_ (_11261_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _34873_ (_13127_, _11261_, _11260_);
  and _34874_ (_11262_, _11254_, _09526_);
  and _34875_ (_11263_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _34876_ (_13128_, _11263_, _11262_);
  and _34877_ (_11264_, _11254_, _09529_);
  and _34878_ (_11265_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _34879_ (_13129_, _11265_, _11264_);
  and _34880_ (_11266_, _11254_, _09532_);
  and _34881_ (_11267_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _34882_ (_13130_, _11267_, _11266_);
  and _34883_ (_11268_, _11254_, _09535_);
  and _34884_ (_11269_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _34885_ (_13132_, _11269_, _11268_);
  and _34886_ (_11270_, _11254_, _09538_);
  and _34887_ (_11271_, _11256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _34888_ (_13133_, _11271_, _11270_);
  and _34889_ (_11272_, _10684_, _10103_);
  and _34890_ (_11273_, _11272_, _09265_);
  and _34891_ (_11274_, _11273_, _09513_);
  not _34892_ (_11275_, _11273_);
  and _34893_ (_11276_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _34894_ (_13134_, _11276_, _11274_);
  and _34895_ (_11277_, _11273_, _09520_);
  and _34896_ (_11278_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _34897_ (_13136_, _11278_, _11277_);
  and _34898_ (_11279_, _11273_, _09523_);
  and _34899_ (_11280_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _34900_ (_13137_, _11280_, _11279_);
  and _34901_ (_11281_, _11273_, _09526_);
  and _34902_ (_11282_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _34903_ (_13138_, _11282_, _11281_);
  and _34904_ (_11283_, _11273_, _09529_);
  and _34905_ (_11284_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _34906_ (_13140_, _11284_, _11283_);
  and _34907_ (_11285_, _11273_, _09532_);
  and _34908_ (_11286_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _34909_ (_13141_, _11286_, _11285_);
  and _34910_ (_11287_, _11273_, _09535_);
  and _34911_ (_11288_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _34912_ (_13142_, _11288_, _11287_);
  and _34913_ (_11289_, _11273_, _09538_);
  and _34914_ (_11290_, _11275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _34915_ (_13143_, _11290_, _11289_);
  and _34916_ (_11291_, _11272_, _09515_);
  and _34917_ (_11292_, _11291_, _09513_);
  not _34918_ (_11293_, _11291_);
  and _34919_ (_11294_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or _34920_ (_13144_, _11294_, _11292_);
  and _34921_ (_11295_, _11291_, _09520_);
  and _34922_ (_11296_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or _34923_ (_13145_, _11296_, _11295_);
  and _34924_ (_11297_, _11291_, _09523_);
  and _34925_ (_11298_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or _34926_ (_13146_, _11298_, _11297_);
  and _34927_ (_11299_, _11291_, _09526_);
  and _34928_ (_11300_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or _34929_ (_13148_, _11300_, _11299_);
  and _34930_ (_11301_, _11291_, _09529_);
  and _34931_ (_11302_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or _34932_ (_13149_, _11302_, _11301_);
  and _34933_ (_11303_, _11291_, _09532_);
  and _34934_ (_11304_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or _34935_ (_13150_, _11304_, _11303_);
  and _34936_ (_11305_, _11291_, _09535_);
  and _34937_ (_11306_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or _34938_ (_13152_, _11306_, _11305_);
  and _34939_ (_11307_, _11291_, _09538_);
  and _34940_ (_11308_, _11293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or _34941_ (_13153_, _11308_, _11307_);
  and _34942_ (_11309_, _11272_, _09542_);
  and _34943_ (_11310_, _11309_, _09513_);
  not _34944_ (_11311_, _11309_);
  and _34945_ (_11312_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or _34946_ (_13154_, _11312_, _11310_);
  and _34947_ (_11313_, _11309_, _09520_);
  and _34948_ (_11314_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or _34949_ (_13155_, _11314_, _11313_);
  and _34950_ (_11315_, _11309_, _09523_);
  and _34951_ (_11316_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or _34952_ (_13156_, _11316_, _11315_);
  and _34953_ (_11317_, _11309_, _09526_);
  and _34954_ (_11318_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or _34955_ (_13157_, _11318_, _11317_);
  and _34956_ (_11319_, _11309_, _09529_);
  and _34957_ (_11320_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or _34958_ (_13158_, _11320_, _11319_);
  and _34959_ (_11321_, _11309_, _09532_);
  and _34960_ (_11322_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or _34961_ (_13160_, _11322_, _11321_);
  and _34962_ (_11323_, _11309_, _09535_);
  and _34963_ (_11324_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or _34964_ (_13161_, _11324_, _11323_);
  and _34965_ (_11325_, _11309_, _09538_);
  and _34966_ (_11326_, _11311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or _34967_ (_13162_, _11326_, _11325_);
  and _34968_ (_11327_, _11272_, _09562_);
  and _34969_ (_11328_, _11327_, _09513_);
  not _34970_ (_11329_, _11327_);
  and _34971_ (_11330_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _34972_ (_13164_, _11330_, _11328_);
  and _34973_ (_11331_, _11327_, _09520_);
  and _34974_ (_11332_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _34975_ (_13165_, _11332_, _11331_);
  and _34976_ (_11333_, _11327_, _09523_);
  and _34977_ (_11334_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _34978_ (_13166_, _11334_, _11333_);
  and _34979_ (_11335_, _11327_, _09526_);
  and _34980_ (_11336_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _34981_ (_13167_, _11336_, _11335_);
  and _34982_ (_11337_, _11327_, _09529_);
  and _34983_ (_11338_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _34984_ (_13168_, _11338_, _11337_);
  and _34985_ (_11339_, _11327_, _09532_);
  and _34986_ (_11340_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _34987_ (_13169_, _11340_, _11339_);
  and _34988_ (_11341_, _11327_, _09535_);
  and _34989_ (_11342_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _34990_ (_13170_, _11342_, _11341_);
  and _34991_ (_11343_, _11327_, _09538_);
  and _34992_ (_11344_, _11329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _34993_ (_13172_, _11344_, _11343_);
  and _34994_ (_11345_, _11272_, _09582_);
  and _34995_ (_11346_, _11345_, _09513_);
  not _34996_ (_11347_, _11345_);
  and _34997_ (_11348_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _34998_ (_13173_, _11348_, _11346_);
  and _34999_ (_11349_, _11345_, _09520_);
  and _35000_ (_11350_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _35001_ (_13174_, _11350_, _11349_);
  and _35002_ (_11351_, _11345_, _09523_);
  and _35003_ (_11352_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _35004_ (_13176_, _11352_, _11351_);
  and _35005_ (_11353_, _11345_, _09526_);
  and _35006_ (_11354_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _35007_ (_13177_, _11354_, _11353_);
  and _35008_ (_11355_, _11345_, _09529_);
  and _35009_ (_11356_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _35010_ (_13178_, _11356_, _11355_);
  and _35011_ (_11357_, _11345_, _09532_);
  and _35012_ (_11358_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _35013_ (_13179_, _11358_, _11357_);
  and _35014_ (_11359_, _11345_, _09535_);
  and _35015_ (_11360_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _35016_ (_13180_, _11360_, _11359_);
  and _35017_ (_11361_, _11345_, _09538_);
  and _35018_ (_11362_, _11347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _35019_ (_13181_, _11362_, _11361_);
  and _35020_ (_11363_, _11272_, _09601_);
  and _35021_ (_11364_, _11363_, _09513_);
  not _35022_ (_11365_, _11363_);
  and _35023_ (_11366_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or _35024_ (_13182_, _11366_, _11364_);
  and _35025_ (_11367_, _11363_, _09520_);
  and _35026_ (_11368_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or _35027_ (_13184_, _11368_, _11367_);
  and _35028_ (_11369_, _11363_, _09523_);
  and _35029_ (_11370_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or _35030_ (_13185_, _11370_, _11369_);
  and _35031_ (_11371_, _11363_, _09526_);
  and _35032_ (_11372_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or _35033_ (_13186_, _11372_, _11371_);
  and _35034_ (_11373_, _11363_, _09529_);
  and _35035_ (_11374_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or _35036_ (_13188_, _11374_, _11373_);
  and _35037_ (_11375_, _11363_, _09532_);
  and _35038_ (_11376_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or _35039_ (_13189_, _11376_, _11375_);
  and _35040_ (_11377_, _11363_, _09535_);
  and _35041_ (_11378_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or _35042_ (_13190_, _11378_, _11377_);
  and _35043_ (_11379_, _11363_, _09538_);
  and _35044_ (_11380_, _11365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or _35045_ (_13191_, _11380_, _11379_);
  and _35046_ (_11381_, _11272_, _09620_);
  and _35047_ (_11382_, _11381_, _09513_);
  not _35048_ (_11383_, _11381_);
  and _35049_ (_11384_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or _35050_ (_13192_, _11384_, _11382_);
  and _35051_ (_11385_, _11381_, _09520_);
  and _35052_ (_11386_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or _35053_ (_13193_, _11386_, _11385_);
  and _35054_ (_11387_, _11381_, _09523_);
  and _35055_ (_11388_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or _35056_ (_13194_, _11388_, _11387_);
  and _35057_ (_11389_, _11381_, _09526_);
  and _35058_ (_11390_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or _35059_ (_13196_, _11390_, _11389_);
  and _35060_ (_11391_, _11381_, _09529_);
  and _35061_ (_11392_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or _35062_ (_13197_, _11392_, _11391_);
  and _35063_ (_11393_, _11381_, _09532_);
  and _35064_ (_11394_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or _35065_ (_13198_, _11394_, _11393_);
  and _35066_ (_11395_, _11381_, _09535_);
  and _35067_ (_11396_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or _35068_ (_13200_, _11396_, _11395_);
  and _35069_ (_11397_, _11381_, _09538_);
  and _35070_ (_11398_, _11383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or _35071_ (_13201_, _11398_, _11397_);
  and _35072_ (_11399_, _11272_, _09639_);
  and _35073_ (_11400_, _11399_, _09513_);
  not _35074_ (_11401_, _11399_);
  and _35075_ (_11402_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _35076_ (_13202_, _11402_, _11400_);
  and _35077_ (_11403_, _11399_, _09520_);
  and _35078_ (_11404_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _35079_ (_13203_, _11404_, _11403_);
  and _35080_ (_11405_, _11399_, _09523_);
  and _35081_ (_11406_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _35082_ (_13204_, _11406_, _11405_);
  and _35083_ (_11407_, _11399_, _09526_);
  and _35084_ (_11408_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _35085_ (_13205_, _11408_, _11407_);
  and _35086_ (_11409_, _11399_, _09529_);
  and _35087_ (_11410_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _35088_ (_13206_, _11410_, _11409_);
  and _35089_ (_11411_, _11399_, _09532_);
  and _35090_ (_11412_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _35091_ (_13208_, _11412_, _11411_);
  and _35092_ (_11413_, _11399_, _09535_);
  and _35093_ (_11414_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _35094_ (_13209_, _11414_, _11413_);
  and _35095_ (_11415_, _11399_, _09538_);
  and _35096_ (_11416_, _11401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _35097_ (_13210_, _11416_, _11415_);
  and _35098_ (_11417_, _11272_, _09659_);
  and _35099_ (_11418_, _11417_, _09513_);
  not _35100_ (_11419_, _11417_);
  and _35101_ (_11420_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or _35102_ (_13212_, _11420_, _11418_);
  and _35103_ (_11421_, _11417_, _09520_);
  and _35104_ (_11422_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or _35105_ (_13213_, _11422_, _11421_);
  and _35106_ (_11423_, _11417_, _09523_);
  and _35107_ (_11424_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or _35108_ (_13214_, _11424_, _11423_);
  and _35109_ (_11425_, _11417_, _09526_);
  and _35110_ (_11426_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or _35111_ (_13215_, _11426_, _11425_);
  and _35112_ (_11427_, _11417_, _09529_);
  and _35113_ (_11428_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or _35114_ (_13216_, _11428_, _11427_);
  and _35115_ (_11429_, _11417_, _09532_);
  and _35116_ (_11430_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or _35117_ (_13217_, _11430_, _11429_);
  and _35118_ (_11431_, _11417_, _09535_);
  and _35119_ (_11432_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or _35120_ (_13218_, _11432_, _11431_);
  and _35121_ (_11433_, _11417_, _09538_);
  and _35122_ (_11434_, _11419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or _35123_ (_13220_, _11434_, _11433_);
  and _35124_ (_11435_, _11272_, _09678_);
  and _35125_ (_11436_, _11435_, _09513_);
  not _35126_ (_11437_, _11435_);
  and _35127_ (_11438_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _35128_ (_13221_, _11438_, _11436_);
  and _35129_ (_11439_, _11435_, _09520_);
  and _35130_ (_11440_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _35131_ (_13222_, _11440_, _11439_);
  and _35132_ (_11441_, _11435_, _09523_);
  and _35133_ (_11442_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _35134_ (_13224_, _11442_, _11441_);
  and _35135_ (_11443_, _11435_, _09526_);
  and _35136_ (_11444_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _35137_ (_13225_, _11444_, _11443_);
  and _35138_ (_11445_, _11435_, _09529_);
  and _35139_ (_11446_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _35140_ (_13226_, _11446_, _11445_);
  and _35141_ (_11447_, _11435_, _09532_);
  and _35142_ (_11448_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _35143_ (_13227_, _11448_, _11447_);
  and _35144_ (_11449_, _11435_, _09535_);
  and _35145_ (_11450_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _35146_ (_13228_, _11450_, _11449_);
  and _35147_ (_11451_, _11435_, _09538_);
  and _35148_ (_11452_, _11437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _35149_ (_13229_, _11452_, _11451_);
  and _35150_ (_11453_, _11272_, _09697_);
  and _35151_ (_11454_, _11453_, _09513_);
  not _35152_ (_11455_, _11453_);
  and _35153_ (_11456_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _35154_ (_13230_, _11456_, _11454_);
  and _35155_ (_11457_, _11453_, _09520_);
  and _35156_ (_11458_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _35157_ (_13232_, _11458_, _11457_);
  and _35158_ (_11459_, _11453_, _09523_);
  and _35159_ (_11460_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _35160_ (_13233_, _11460_, _11459_);
  and _35161_ (_11461_, _11453_, _09526_);
  and _35162_ (_11462_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _35163_ (_13234_, _11462_, _11461_);
  and _35164_ (_11463_, _11453_, _09529_);
  and _35165_ (_11464_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _35166_ (_13236_, _11464_, _11463_);
  and _35167_ (_11465_, _11453_, _09532_);
  and _35168_ (_11466_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _35169_ (_13237_, _11466_, _11465_);
  and _35170_ (_11467_, _11453_, _09535_);
  and _35171_ (_11468_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _35172_ (_13238_, _11468_, _11467_);
  and _35173_ (_11469_, _11453_, _09538_);
  and _35174_ (_11470_, _11455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _35175_ (_13239_, _11470_, _11469_);
  and _35176_ (_11471_, _11272_, _09716_);
  and _35177_ (_11472_, _11471_, _09513_);
  not _35178_ (_11473_, _11471_);
  and _35179_ (_11474_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or _35180_ (_13241_, _11474_, _11472_);
  and _35181_ (_11475_, _11471_, _09520_);
  and _35182_ (_11476_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or _35183_ (_13242_, _11476_, _11475_);
  and _35184_ (_11477_, _11471_, _09523_);
  and _35185_ (_11478_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or _35186_ (_13243_, _11478_, _11477_);
  and _35187_ (_11479_, _11471_, _09526_);
  and _35188_ (_11480_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or _35189_ (_13245_, _11480_, _11479_);
  and _35190_ (_11481_, _11471_, _09529_);
  and _35191_ (_11482_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or _35192_ (_13246_, _11482_, _11481_);
  and _35193_ (_11483_, _11471_, _09532_);
  and _35194_ (_11484_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or _35195_ (_13247_, _11484_, _11483_);
  and _35196_ (_11485_, _11471_, _09535_);
  and _35197_ (_11486_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or _35198_ (_13248_, _11486_, _11485_);
  and _35199_ (_11487_, _11471_, _09538_);
  and _35200_ (_11488_, _11473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or _35201_ (_13249_, _11488_, _11487_);
  and _35202_ (_11489_, _11272_, _09736_);
  and _35203_ (_11490_, _11489_, _09513_);
  not _35204_ (_11491_, _11489_);
  and _35205_ (_11492_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or _35206_ (_13250_, _11492_, _11490_);
  and _35207_ (_11493_, _11489_, _09520_);
  and _35208_ (_11494_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or _35209_ (_13252_, _11494_, _11493_);
  and _35210_ (_11495_, _11489_, _09523_);
  and _35211_ (_11496_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or _35212_ (_13253_, _11496_, _11495_);
  and _35213_ (_11497_, _11489_, _09526_);
  and _35214_ (_11498_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or _35215_ (_13254_, _11498_, _11497_);
  and _35216_ (_11499_, _11489_, _09529_);
  and _35217_ (_11500_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or _35218_ (_13255_, _11500_, _11499_);
  and _35219_ (_11501_, _11489_, _09532_);
  and _35220_ (_11502_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or _35221_ (_13257_, _11502_, _11501_);
  and _35222_ (_11503_, _11489_, _09535_);
  and _35223_ (_11504_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or _35224_ (_13258_, _11504_, _11503_);
  and _35225_ (_11505_, _11489_, _09538_);
  and _35226_ (_11506_, _11491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or _35227_ (_13259_, _11506_, _11505_);
  and _35228_ (_11507_, _11272_, _09755_);
  and _35229_ (_11508_, _11507_, _09513_);
  not _35230_ (_11509_, _11507_);
  and _35231_ (_11510_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _35232_ (_13260_, _11510_, _11508_);
  and _35233_ (_11511_, _11507_, _09520_);
  and _35234_ (_11512_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _35235_ (_13261_, _11512_, _11511_);
  and _35236_ (_11513_, _11507_, _09523_);
  and _35237_ (_11514_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _35238_ (_13262_, _11514_, _11513_);
  and _35239_ (_11515_, _11507_, _09526_);
  and _35240_ (_11516_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _35241_ (_13264_, _11516_, _11515_);
  and _35242_ (_11517_, _11507_, _09529_);
  and _35243_ (_11518_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _35244_ (_13265_, _11518_, _11517_);
  and _35245_ (_11519_, _11507_, _09532_);
  and _35246_ (_11520_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _35247_ (_13266_, _11520_, _11519_);
  and _35248_ (_11521_, _11507_, _09535_);
  and _35249_ (_11522_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _35250_ (_13267_, _11522_, _11521_);
  and _35251_ (_11523_, _11507_, _09538_);
  and _35252_ (_11524_, _11509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _35253_ (_13269_, _11524_, _11523_);
  and _35254_ (_11525_, _11272_, _09774_);
  and _35255_ (_11526_, _11525_, _09513_);
  not _35256_ (_11527_, _11525_);
  and _35257_ (_11528_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _35258_ (_13270_, _11528_, _11526_);
  and _35259_ (_11529_, _11525_, _09520_);
  and _35260_ (_11530_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _35261_ (_13271_, _11530_, _11529_);
  and _35262_ (_11531_, _11525_, _09523_);
  and _35263_ (_11532_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _35264_ (_13272_, _11532_, _11531_);
  and _35265_ (_11533_, _11525_, _09526_);
  and _35266_ (_11534_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _35267_ (_13273_, _11534_, _11533_);
  and _35268_ (_11535_, _11525_, _09529_);
  and _35269_ (_11536_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _35270_ (_13274_, _11536_, _11535_);
  and _35271_ (_11537_, _11525_, _09532_);
  and _35272_ (_11538_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _35273_ (_13276_, _11538_, _11537_);
  and _35274_ (_11539_, _11525_, _09535_);
  and _35275_ (_11540_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _35276_ (_13277_, _11540_, _11539_);
  and _35277_ (_11541_, _11525_, _09538_);
  and _35278_ (_11542_, _11527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _35279_ (_13278_, _11542_, _11541_);
  and _35280_ (_11543_, _11272_, _09793_);
  and _35281_ (_11544_, _11543_, _09513_);
  not _35282_ (_11545_, _11543_);
  and _35283_ (_11546_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or _35284_ (_13279_, _11546_, _11544_);
  and _35285_ (_11547_, _11543_, _09520_);
  and _35286_ (_11548_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or _35287_ (_13281_, _11548_, _11547_);
  and _35288_ (_11549_, _11543_, _09523_);
  and _35289_ (_11550_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or _35290_ (_13282_, _11550_, _11549_);
  and _35291_ (_11551_, _11543_, _09526_);
  and _35292_ (_11552_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or _35293_ (_13283_, _11552_, _11551_);
  and _35294_ (_11553_, _11543_, _09529_);
  and _35295_ (_11554_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or _35296_ (_13284_, _11554_, _11553_);
  and _35297_ (_11555_, _11543_, _09532_);
  and _35298_ (_11556_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or _35299_ (_13285_, _11556_, _11555_);
  and _35300_ (_11557_, _11543_, _09535_);
  and _35301_ (_11558_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or _35302_ (_13286_, _11558_, _11557_);
  and _35303_ (_11559_, _11543_, _09538_);
  and _35304_ (_11560_, _11545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or _35305_ (_13287_, _11560_, _11559_);
  and _35306_ (_11561_, _10684_, _10393_);
  and _35307_ (_11562_, _11561_, _09265_);
  and _35308_ (_11563_, _11562_, _09513_);
  not _35309_ (_11564_, _11562_);
  and _35310_ (_11565_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or _35311_ (_13289_, _11565_, _11563_);
  and _35312_ (_11566_, _11562_, _09520_);
  and _35313_ (_11567_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or _35314_ (_13290_, _11567_, _11566_);
  and _35315_ (_11568_, _11562_, _09523_);
  and _35316_ (_11569_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or _35317_ (_13292_, _11569_, _11568_);
  and _35318_ (_11570_, _11562_, _09526_);
  and _35319_ (_11571_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or _35320_ (_13293_, _11571_, _11570_);
  and _35321_ (_11572_, _11562_, _09529_);
  and _35322_ (_11573_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or _35323_ (_13294_, _11573_, _11572_);
  and _35324_ (_11574_, _11562_, _09532_);
  and _35325_ (_11575_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or _35326_ (_13295_, _11575_, _11574_);
  and _35327_ (_11576_, _11562_, _09535_);
  and _35328_ (_11577_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or _35329_ (_13296_, _11577_, _11576_);
  and _35330_ (_11578_, _11562_, _09538_);
  and _35331_ (_11579_, _11564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or _35332_ (_13297_, _11579_, _11578_);
  and _35333_ (_11580_, _11561_, _09515_);
  and _35334_ (_11581_, _11580_, _09513_);
  not _35335_ (_11582_, _11580_);
  and _35336_ (_11583_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _35337_ (_13298_, _11583_, _11581_);
  and _35338_ (_11584_, _11580_, _09520_);
  and _35339_ (_11585_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _35340_ (_13300_, _11585_, _11584_);
  and _35341_ (_11586_, _11580_, _09523_);
  and _35342_ (_11587_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _35343_ (_13301_, _11587_, _11586_);
  and _35344_ (_11588_, _11580_, _09526_);
  and _35345_ (_11589_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _35346_ (_13302_, _11589_, _11588_);
  and _35347_ (_11590_, _11580_, _09529_);
  and _35348_ (_11591_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _35349_ (_13304_, _11591_, _11590_);
  and _35350_ (_11592_, _11580_, _09532_);
  and _35351_ (_11593_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _35352_ (_13305_, _11593_, _11592_);
  and _35353_ (_11594_, _11580_, _09535_);
  and _35354_ (_11595_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _35355_ (_13306_, _11595_, _11594_);
  and _35356_ (_11596_, _11580_, _09538_);
  and _35357_ (_11597_, _11582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _35358_ (_13307_, _11597_, _11596_);
  and _35359_ (_11598_, _11561_, _09542_);
  and _35360_ (_11599_, _11598_, _09513_);
  not _35361_ (_11600_, _11598_);
  and _35362_ (_11601_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _35363_ (_13308_, _11601_, _11599_);
  and _35364_ (_11602_, _11598_, _09520_);
  and _35365_ (_11603_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _35366_ (_13309_, _11603_, _11602_);
  and _35367_ (_11604_, _11598_, _09523_);
  and _35368_ (_11605_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _35369_ (_13310_, _11605_, _11604_);
  and _35370_ (_11606_, _11598_, _09526_);
  and _35371_ (_11607_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _35372_ (_13312_, _11607_, _11606_);
  and _35373_ (_11608_, _11598_, _09529_);
  and _35374_ (_11609_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _35375_ (_13313_, _11609_, _11608_);
  and _35376_ (_11610_, _11598_, _09532_);
  and _35377_ (_11611_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _35378_ (_13314_, _11611_, _11610_);
  and _35379_ (_11612_, _11598_, _09535_);
  and _35380_ (_11613_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _35381_ (_13316_, _11613_, _11612_);
  and _35382_ (_11614_, _11598_, _09538_);
  and _35383_ (_11615_, _11600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _35384_ (_13317_, _11615_, _11614_);
  and _35385_ (_11616_, _11561_, _09562_);
  and _35386_ (_11617_, _11616_, _09513_);
  not _35387_ (_11618_, _11616_);
  and _35388_ (_11619_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or _35389_ (_13318_, _11619_, _11617_);
  and _35390_ (_11620_, _11616_, _09520_);
  and _35391_ (_11621_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or _35392_ (_13319_, _11621_, _11620_);
  and _35393_ (_11622_, _11616_, _09523_);
  and _35394_ (_11623_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or _35395_ (_13320_, _11623_, _11622_);
  and _35396_ (_11624_, _11616_, _09526_);
  and _35397_ (_11625_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or _35398_ (_13321_, _11625_, _11624_);
  and _35399_ (_11626_, _11616_, _09529_);
  and _35400_ (_11627_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or _35401_ (_13322_, _11627_, _11626_);
  and _35402_ (_11628_, _11616_, _09532_);
  and _35403_ (_11629_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or _35404_ (_13324_, _11629_, _11628_);
  and _35405_ (_11630_, _11616_, _09535_);
  and _35406_ (_11631_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or _35407_ (_13325_, _11631_, _11630_);
  and _35408_ (_11632_, _11616_, _09538_);
  and _35409_ (_11633_, _11618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or _35410_ (_13326_, _11633_, _11632_);
  and _35411_ (_11634_, _11561_, _09582_);
  and _35412_ (_11635_, _11634_, _09513_);
  not _35413_ (_11636_, _11634_);
  and _35414_ (_11637_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or _35415_ (_13328_, _11637_, _11635_);
  and _35416_ (_11638_, _11634_, _09520_);
  and _35417_ (_11639_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or _35418_ (_13329_, _11639_, _11638_);
  and _35419_ (_11640_, _11634_, _09523_);
  and _35420_ (_11641_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or _35421_ (_13330_, _11641_, _11640_);
  and _35422_ (_11642_, _11634_, _09526_);
  and _35423_ (_11643_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or _35424_ (_13331_, _11643_, _11642_);
  and _35425_ (_11644_, _11634_, _09529_);
  and _35426_ (_11645_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or _35427_ (_13332_, _11645_, _11644_);
  and _35428_ (_11646_, _11634_, _09532_);
  and _35429_ (_11647_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or _35430_ (_13333_, _11647_, _11646_);
  and _35431_ (_11648_, _11634_, _09535_);
  and _35432_ (_11649_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or _35433_ (_13334_, _11649_, _11648_);
  and _35434_ (_11650_, _11634_, _09538_);
  and _35435_ (_11651_, _11636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or _35436_ (_13336_, _11651_, _11650_);
  and _35437_ (_11652_, _11561_, _09601_);
  and _35438_ (_11653_, _11652_, _09513_);
  not _35439_ (_11654_, _11652_);
  and _35440_ (_11655_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _35441_ (_13337_, _11655_, _11653_);
  and _35442_ (_11656_, _11652_, _09520_);
  and _35443_ (_11657_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _35444_ (_13338_, _11657_, _11656_);
  and _35445_ (_11658_, _11652_, _09523_);
  and _35446_ (_11659_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _35447_ (_13340_, _11659_, _11658_);
  and _35448_ (_11660_, _11652_, _09526_);
  and _35449_ (_11661_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _35450_ (_13341_, _11661_, _11660_);
  and _35451_ (_11662_, _11652_, _09529_);
  and _35452_ (_11663_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _35453_ (_13342_, _11663_, _11662_);
  and _35454_ (_11664_, _11652_, _09532_);
  and _35455_ (_11665_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _35456_ (_13343_, _11665_, _11664_);
  and _35457_ (_11666_, _11652_, _09535_);
  and _35458_ (_11667_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _35459_ (_13345_, _11667_, _11666_);
  and _35460_ (_11668_, _11652_, _09538_);
  and _35461_ (_11669_, _11654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _35462_ (_13346_, _11669_, _11668_);
  and _35463_ (_11670_, _11561_, _09620_);
  and _35464_ (_11671_, _11670_, _09513_);
  not _35465_ (_11672_, _11670_);
  and _35466_ (_11673_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _35467_ (_13347_, _11673_, _11671_);
  and _35468_ (_11674_, _11670_, _09520_);
  and _35469_ (_11675_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _35470_ (_13349_, _11675_, _11674_);
  and _35471_ (_11676_, _11670_, _09523_);
  and _35472_ (_11677_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _35473_ (_13350_, _11677_, _11676_);
  and _35474_ (_11678_, _11670_, _09526_);
  and _35475_ (_11679_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _35476_ (_13351_, _11679_, _11678_);
  and _35477_ (_11680_, _11670_, _09529_);
  and _35478_ (_11681_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _35479_ (_13352_, _11681_, _11680_);
  and _35480_ (_11682_, _11670_, _09532_);
  and _35481_ (_11683_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _35482_ (_13353_, _11683_, _11682_);
  and _35483_ (_11684_, _11670_, _09535_);
  and _35484_ (_11685_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _35485_ (_13354_, _11685_, _11684_);
  and _35486_ (_11686_, _11670_, _09538_);
  and _35487_ (_11687_, _11672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _35488_ (_13355_, _11687_, _11686_);
  and _35489_ (_11688_, _11561_, _09639_);
  and _35490_ (_11689_, _11688_, _09513_);
  not _35491_ (_11690_, _11688_);
  and _35492_ (_11691_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or _35493_ (_13357_, _11691_, _11689_);
  and _35494_ (_11692_, _11688_, _09520_);
  and _35495_ (_11693_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or _35496_ (_13358_, _11693_, _11692_);
  and _35497_ (_11694_, _11688_, _09523_);
  and _35498_ (_11695_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or _35499_ (_13359_, _11695_, _11694_);
  and _35500_ (_11696_, _11688_, _09526_);
  and _35501_ (_11697_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or _35502_ (_13361_, _11697_, _11696_);
  and _35503_ (_11698_, _11688_, _09529_);
  and _35504_ (_11699_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or _35505_ (_13362_, _11699_, _11698_);
  and _35506_ (_11700_, _11688_, _09532_);
  and _35507_ (_11701_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or _35508_ (_13363_, _11701_, _11700_);
  and _35509_ (_11702_, _11688_, _09535_);
  and _35510_ (_11703_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or _35511_ (_13364_, _11703_, _11702_);
  and _35512_ (_11704_, _11688_, _09538_);
  and _35513_ (_11705_, _11690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or _35514_ (_13365_, _11705_, _11704_);
  and _35515_ (_11706_, _11561_, _09659_);
  and _35516_ (_11707_, _11706_, _09513_);
  not _35517_ (_11708_, _11706_);
  and _35518_ (_11709_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _35519_ (_13366_, _11709_, _11707_);
  and _35520_ (_11710_, _11706_, _09520_);
  and _35521_ (_11711_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _35522_ (_13367_, _11711_, _11710_);
  and _35523_ (_11712_, _11706_, _09523_);
  and _35524_ (_11713_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _35525_ (_13369_, _11713_, _11712_);
  and _35526_ (_11714_, _11706_, _09526_);
  and _35527_ (_11715_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _35528_ (_13370_, _11715_, _11714_);
  and _35529_ (_11716_, _11706_, _09529_);
  and _35530_ (_11717_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _35531_ (_13371_, _11717_, _11716_);
  and _35532_ (_11718_, _11706_, _09532_);
  and _35533_ (_11719_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _35534_ (_13373_, _11719_, _11718_);
  and _35535_ (_11720_, _11706_, _09535_);
  and _35536_ (_11721_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _35537_ (_13374_, _11721_, _11720_);
  and _35538_ (_11722_, _11706_, _09538_);
  and _35539_ (_11723_, _11708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _35540_ (_13375_, _11723_, _11722_);
  and _35541_ (_11724_, _11561_, _09678_);
  and _35542_ (_11725_, _11724_, _09513_);
  not _35543_ (_11726_, _11724_);
  and _35544_ (_11727_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or _35545_ (_13376_, _11727_, _11725_);
  and _35546_ (_11728_, _11724_, _09520_);
  and _35547_ (_11729_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or _35548_ (_13377_, _11729_, _11728_);
  and _35549_ (_11730_, _11724_, _09523_);
  and _35550_ (_11731_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or _35551_ (_13378_, _11731_, _11730_);
  and _35552_ (_11732_, _11724_, _09526_);
  and _35553_ (_11733_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or _35554_ (_13379_, _11733_, _11732_);
  and _35555_ (_11734_, _11724_, _09529_);
  and _35556_ (_11735_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or _35557_ (_13381_, _11735_, _11734_);
  and _35558_ (_11736_, _11724_, _09532_);
  and _35559_ (_11737_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or _35560_ (_13382_, _11737_, _11736_);
  and _35561_ (_11738_, _11724_, _09535_);
  and _35562_ (_11739_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or _35563_ (_13383_, _11739_, _11738_);
  and _35564_ (_11740_, _11724_, _09538_);
  and _35565_ (_11741_, _11726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or _35566_ (_13385_, _11741_, _11740_);
  and _35567_ (_11742_, _11561_, _09697_);
  and _35568_ (_11743_, _11742_, _09513_);
  not _35569_ (_11744_, _11742_);
  and _35570_ (_11745_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or _35571_ (_13386_, _11745_, _11743_);
  and _35572_ (_11746_, _11742_, _09520_);
  and _35573_ (_11747_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or _35574_ (_13387_, _11747_, _11746_);
  and _35575_ (_11748_, _11742_, _09523_);
  and _35576_ (_11749_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or _35577_ (_13388_, _11749_, _11748_);
  and _35578_ (_11750_, _11742_, _09526_);
  and _35579_ (_11751_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or _35580_ (_13389_, _11751_, _11750_);
  and _35581_ (_11752_, _11742_, _09529_);
  and _35582_ (_11753_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or _35583_ (_13390_, _11753_, _11752_);
  and _35584_ (_11754_, _11742_, _09532_);
  and _35585_ (_11755_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or _35586_ (_13391_, _11755_, _11754_);
  and _35587_ (_11756_, _11742_, _09535_);
  and _35588_ (_11757_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or _35589_ (_13393_, _11757_, _11756_);
  and _35590_ (_11758_, _11742_, _09538_);
  and _35591_ (_11759_, _11744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or _35592_ (_13394_, _11759_, _11758_);
  and _35593_ (_11760_, _11561_, _09716_);
  and _35594_ (_11761_, _11760_, _09513_);
  not _35595_ (_11762_, _11760_);
  and _35596_ (_11763_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _35597_ (_13395_, _11763_, _11761_);
  and _35598_ (_11764_, _11760_, _09520_);
  and _35599_ (_11765_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _35600_ (_13397_, _11765_, _11764_);
  and _35601_ (_11766_, _11760_, _09523_);
  and _35602_ (_11767_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _35603_ (_13398_, _11767_, _11766_);
  and _35604_ (_11768_, _11760_, _09526_);
  and _35605_ (_11769_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _35606_ (_13399_, _11769_, _11768_);
  and _35607_ (_11770_, _11760_, _09529_);
  and _35608_ (_11771_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _35609_ (_13400_, _11771_, _11770_);
  and _35610_ (_11772_, _11760_, _09532_);
  and _35611_ (_11773_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _35612_ (_13401_, _11773_, _11772_);
  and _35613_ (_11774_, _11760_, _09535_);
  and _35614_ (_11775_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _35615_ (_13402_, _11775_, _11774_);
  and _35616_ (_11776_, _11760_, _09538_);
  and _35617_ (_11777_, _11762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _35618_ (_13403_, _11777_, _11776_);
  and _35619_ (_11778_, _11561_, _09736_);
  and _35620_ (_11779_, _11778_, _09513_);
  not _35621_ (_11780_, _11778_);
  and _35622_ (_11781_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _35623_ (_13405_, _11781_, _11779_);
  and _35624_ (_11782_, _11778_, _09520_);
  and _35625_ (_11783_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _35626_ (_13406_, _11783_, _11782_);
  and _35627_ (_11784_, _11778_, _09523_);
  and _35628_ (_11785_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _35629_ (_13407_, _11785_, _11784_);
  and _35630_ (_11786_, _11778_, _09526_);
  and _35631_ (_11787_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _35632_ (_13409_, _11787_, _11786_);
  and _35633_ (_11788_, _11778_, _09529_);
  and _35634_ (_11789_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _35635_ (_13410_, _11789_, _11788_);
  and _35636_ (_11790_, _11778_, _09532_);
  and _35637_ (_11791_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _35638_ (_13411_, _11791_, _11790_);
  and _35639_ (_11792_, _11778_, _09535_);
  and _35640_ (_11793_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _35641_ (_13412_, _11793_, _11792_);
  and _35642_ (_11794_, _11778_, _09538_);
  and _35643_ (_11795_, _11780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _35644_ (_13413_, _11795_, _11794_);
  and _35645_ (_11796_, _11561_, _09755_);
  and _35646_ (_11797_, _11796_, _09513_);
  not _35647_ (_11798_, _11796_);
  and _35648_ (_11799_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or _35649_ (_13414_, _11799_, _11797_);
  and _35650_ (_11800_, _11796_, _09520_);
  and _35651_ (_11801_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or _35652_ (_13415_, _11801_, _11800_);
  and _35653_ (_11802_, _11796_, _09523_);
  and _35654_ (_11803_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or _35655_ (_13417_, _11803_, _11802_);
  and _35656_ (_11804_, _11796_, _09526_);
  and _35657_ (_11805_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or _35658_ (_13418_, _11805_, _11804_);
  and _35659_ (_11806_, _11796_, _09529_);
  and _35660_ (_11807_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or _35661_ (_13419_, _11807_, _11806_);
  and _35662_ (_11808_, _11796_, _09532_);
  and _35663_ (_11809_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or _35664_ (_13421_, _11809_, _11808_);
  and _35665_ (_11810_, _11796_, _09535_);
  and _35666_ (_11811_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or _35667_ (_13422_, _11811_, _11810_);
  and _35668_ (_11812_, _11796_, _09538_);
  and _35669_ (_11813_, _11798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or _35670_ (_13423_, _11813_, _11812_);
  and _35671_ (_11814_, _11561_, _09774_);
  and _35672_ (_11815_, _11814_, _09513_);
  not _35673_ (_11816_, _11814_);
  and _35674_ (_11817_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or _35675_ (_13424_, _11817_, _11815_);
  and _35676_ (_11818_, _11814_, _09520_);
  and _35677_ (_11819_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or _35678_ (_13425_, _11819_, _11818_);
  and _35679_ (_11820_, _11814_, _09523_);
  and _35680_ (_11821_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or _35681_ (_13426_, _11821_, _11820_);
  and _35682_ (_11822_, _11814_, _09526_);
  and _35683_ (_11823_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or _35684_ (_13427_, _11823_, _11822_);
  and _35685_ (_11824_, _11814_, _09529_);
  and _35686_ (_11825_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or _35687_ (_13429_, _11825_, _11824_);
  and _35688_ (_11826_, _11814_, _09532_);
  and _35689_ (_11827_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or _35690_ (_13430_, _11827_, _11826_);
  and _35691_ (_11828_, _11814_, _09535_);
  and _35692_ (_11829_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or _35693_ (_13431_, _11829_, _11828_);
  and _35694_ (_11830_, _11814_, _09538_);
  and _35695_ (_11831_, _11816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or _35696_ (_13433_, _11831_, _11830_);
  and _35697_ (_11832_, _11561_, _09793_);
  and _35698_ (_11833_, _11832_, _09513_);
  not _35699_ (_11834_, _11832_);
  and _35700_ (_11835_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _35701_ (_13434_, _11835_, _11833_);
  and _35702_ (_11836_, _11832_, _09520_);
  and _35703_ (_11837_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _35704_ (_13435_, _11837_, _11836_);
  and _35705_ (_11838_, _11832_, _09523_);
  and _35706_ (_11839_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _35707_ (_13436_, _11839_, _11838_);
  and _35708_ (_11840_, _11832_, _09526_);
  and _35709_ (_11841_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _35710_ (_13437_, _11841_, _11840_);
  and _35711_ (_11842_, _11832_, _09529_);
  and _35712_ (_11843_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _35713_ (_13438_, _11843_, _11842_);
  and _35714_ (_11844_, _11832_, _09532_);
  and _35715_ (_11845_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _35716_ (_13439_, _11845_, _11844_);
  and _35717_ (_11846_, _11832_, _09535_);
  and _35718_ (_11847_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _35719_ (_13441_, _11847_, _11846_);
  and _35720_ (_11848_, _11832_, _09538_);
  and _35721_ (_11849_, _11834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _35722_ (_13442_, _11849_, _11848_);
  not _35723_ (_11850_, _09265_);
  and _35724_ (_11851_, _06008_, _02161_);
  nand _35725_ (_11852_, _11851_, _09254_);
  or _35726_ (_11853_, _11852_, _11850_);
  and _35727_ (_11854_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  and _35728_ (_11855_, _09254_, _02161_);
  and _35729_ (_11856_, _11855_, _09266_);
  and _35730_ (_11857_, _11856_, _09334_);
  or _35731_ (_13444_, _11857_, _11854_);
  and _35732_ (_11858_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and _35733_ (_11859_, _11856_, _09453_);
  or _35734_ (_13445_, _11859_, _11858_);
  and _35735_ (_11860_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and _35736_ (_11861_, _11856_, _09463_);
  or _35737_ (_13446_, _11861_, _11860_);
  and _35738_ (_11862_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  and _35739_ (_11863_, _11856_, _09472_);
  or _35740_ (_13448_, _11863_, _11862_);
  and _35741_ (_11864_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and _35742_ (_11865_, _11856_, _09482_);
  or _35743_ (_13449_, _11865_, _11864_);
  and _35744_ (_11866_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and _35745_ (_11867_, _11856_, _09492_);
  or _35746_ (_13450_, _11867_, _11866_);
  and _35747_ (_11868_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and _35748_ (_11869_, _11856_, _09502_);
  or _35749_ (_13452_, _11869_, _11868_);
  and _35750_ (_11870_, _11853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  and _35751_ (_11871_, _11856_, _09510_);
  or _35752_ (_13453_, _11871_, _11870_);
  not _35753_ (_11872_, _09515_);
  or _35754_ (_11873_, _11852_, _11872_);
  and _35755_ (_11874_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _35756_ (_11875_, _11855_, _06008_);
  and _35757_ (_11876_, _11875_, _09515_);
  and _35758_ (_11877_, _11876_, _09334_);
  or _35759_ (_13454_, _11877_, _11874_);
  and _35760_ (_11878_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and _35761_ (_11879_, _11876_, _09453_);
  or _35762_ (_13455_, _11879_, _11878_);
  and _35763_ (_11880_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and _35764_ (_11881_, _11876_, _09463_);
  or _35765_ (_13456_, _11881_, _11880_);
  and _35766_ (_11882_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _35767_ (_11883_, _11876_, _09472_);
  or _35768_ (_13457_, _11883_, _11882_);
  and _35769_ (_11884_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and _35770_ (_11885_, _11876_, _09482_);
  or _35771_ (_13458_, _11885_, _11884_);
  and _35772_ (_11886_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _35773_ (_11887_, _11876_, _09492_);
  or _35774_ (_13460_, _11887_, _11886_);
  and _35775_ (_11888_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and _35776_ (_11889_, _11876_, _09502_);
  or _35777_ (_13461_, _11889_, _11888_);
  and _35778_ (_11890_, _11873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and _35779_ (_11891_, _11876_, _09510_);
  or _35780_ (_13462_, _11891_, _11890_);
  not _35781_ (_11892_, _09542_);
  or _35782_ (_11893_, _11852_, _11892_);
  and _35783_ (_11894_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _35784_ (_11895_, _11875_, _09542_);
  and _35785_ (_11896_, _11895_, _09334_);
  or _35786_ (_13464_, _11896_, _11894_);
  and _35787_ (_11897_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _35788_ (_11898_, _11895_, _09453_);
  or _35789_ (_13465_, _11898_, _11897_);
  and _35790_ (_11899_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and _35791_ (_11900_, _11895_, _09463_);
  or _35792_ (_13466_, _11900_, _11899_);
  and _35793_ (_11901_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _35794_ (_11902_, _11895_, _09472_);
  or _35795_ (_13467_, _11902_, _11901_);
  and _35796_ (_11903_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and _35797_ (_11904_, _11895_, _09482_);
  or _35798_ (_13468_, _11904_, _11903_);
  and _35799_ (_11905_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _35800_ (_11906_, _11895_, _09492_);
  or _35801_ (_13469_, _11906_, _11905_);
  and _35802_ (_11907_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and _35803_ (_11908_, _11895_, _09502_);
  or _35804_ (_13470_, _11908_, _11907_);
  and _35805_ (_11909_, _11893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and _35806_ (_11910_, _11895_, _09510_);
  or _35807_ (_13472_, _11910_, _11909_);
  not _35808_ (_11911_, _09562_);
  or _35809_ (_11912_, _11852_, _11911_);
  and _35810_ (_11913_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  and _35811_ (_11914_, _11875_, _09562_);
  and _35812_ (_11915_, _11914_, _09334_);
  or _35813_ (_13473_, _11915_, _11913_);
  and _35814_ (_11916_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  and _35815_ (_11917_, _11914_, _09453_);
  or _35816_ (_13474_, _11917_, _11916_);
  and _35817_ (_11918_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and _35818_ (_11919_, _11914_, _09463_);
  or _35819_ (_13476_, _11919_, _11918_);
  and _35820_ (_11920_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  and _35821_ (_11921_, _11914_, _09472_);
  or _35822_ (_13477_, _11921_, _11920_);
  and _35823_ (_11922_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and _35824_ (_11923_, _11914_, _09482_);
  or _35825_ (_13478_, _11923_, _11922_);
  and _35826_ (_11924_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  and _35827_ (_11925_, _11914_, _09492_);
  or _35828_ (_13479_, _11925_, _11924_);
  and _35829_ (_11926_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  and _35830_ (_11927_, _11914_, _09502_);
  or _35831_ (_13480_, _11927_, _11926_);
  and _35832_ (_11928_, _11912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  and _35833_ (_11929_, _11914_, _09510_);
  or _35834_ (_13481_, _11929_, _11928_);
  not _35835_ (_11930_, _09582_);
  or _35836_ (_11931_, _11852_, _11930_);
  and _35837_ (_11932_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and _35838_ (_11933_, _11875_, _09582_);
  and _35839_ (_11934_, _11933_, _09334_);
  or _35840_ (_13482_, _11934_, _11932_);
  and _35841_ (_11935_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and _35842_ (_11936_, _11933_, _09453_);
  or _35843_ (_13484_, _11936_, _11935_);
  and _35844_ (_11937_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and _35845_ (_11938_, _11933_, _09463_);
  or _35846_ (_13485_, _11938_, _11937_);
  and _35847_ (_11939_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  and _35848_ (_11940_, _11933_, _09472_);
  or _35849_ (_13486_, _11940_, _11939_);
  and _35850_ (_11941_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and _35851_ (_11942_, _11933_, _09482_);
  or _35852_ (_13488_, _11942_, _11941_);
  and _35853_ (_11943_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and _35854_ (_11944_, _11933_, _09492_);
  or _35855_ (_13489_, _11944_, _11943_);
  and _35856_ (_11945_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  and _35857_ (_11946_, _11933_, _09502_);
  or _35858_ (_13490_, _11946_, _11945_);
  and _35859_ (_11947_, _11931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and _35860_ (_11948_, _11933_, _09510_);
  or _35861_ (_13491_, _11948_, _11947_);
  not _35862_ (_11949_, _09601_);
  or _35863_ (_11950_, _11852_, _11949_);
  and _35864_ (_11951_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _35865_ (_11952_, _11875_, _09601_);
  and _35866_ (_11953_, _11952_, _09334_);
  or _35867_ (_13492_, _11953_, _11951_);
  and _35868_ (_11954_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and _35869_ (_11955_, _11952_, _09453_);
  or _35870_ (_13493_, _11955_, _11954_);
  and _35871_ (_11956_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and _35872_ (_11957_, _11952_, _09463_);
  or _35873_ (_13494_, _11957_, _11956_);
  and _35874_ (_11958_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _35875_ (_11959_, _11952_, _09472_);
  or _35876_ (_13496_, _11959_, _11958_);
  and _35877_ (_11960_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and _35878_ (_11961_, _11952_, _09482_);
  or _35879_ (_13497_, _11961_, _11960_);
  and _35880_ (_11962_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _35881_ (_11963_, _11952_, _09492_);
  or _35882_ (_13498_, _11963_, _11962_);
  and _35883_ (_11964_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and _35884_ (_11965_, _11952_, _09502_);
  or _35885_ (_13500_, _11965_, _11964_);
  and _35886_ (_11966_, _11950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and _35887_ (_11967_, _11952_, _09510_);
  or _35888_ (_13501_, _11967_, _11966_);
  not _35889_ (_11968_, _09620_);
  or _35890_ (_11969_, _11852_, _11968_);
  and _35891_ (_11970_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _35892_ (_11971_, _11875_, _09620_);
  and _35893_ (_11972_, _11971_, _09334_);
  or _35894_ (_13502_, _11972_, _11970_);
  and _35895_ (_11973_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and _35896_ (_11974_, _11971_, _09453_);
  or _35897_ (_13503_, _11974_, _11973_);
  and _35898_ (_11975_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _35899_ (_11976_, _11971_, _09463_);
  or _35900_ (_13504_, _11976_, _11975_);
  and _35901_ (_11977_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _35902_ (_11978_, _11971_, _09472_);
  or _35903_ (_13505_, _11978_, _11977_);
  and _35904_ (_11979_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _35905_ (_11980_, _11971_, _09482_);
  or _35906_ (_13506_, _11980_, _11979_);
  and _35907_ (_11981_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _35908_ (_11982_, _11971_, _09492_);
  or _35909_ (_13508_, _11982_, _11981_);
  and _35910_ (_11983_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and _35911_ (_11984_, _11971_, _09502_);
  or _35912_ (_13509_, _11984_, _11983_);
  and _35913_ (_11986_, _11969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and _35914_ (_11987_, _11971_, _09510_);
  or _35915_ (_13510_, _11987_, _11986_);
  not _35916_ (_11988_, _09639_);
  or _35917_ (_11989_, _11852_, _11988_);
  and _35918_ (_11990_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  and _35919_ (_11991_, _11875_, _09639_);
  and _35920_ (_11992_, _11991_, _09334_);
  or _35921_ (_13512_, _11992_, _11990_);
  and _35922_ (_11993_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and _35923_ (_11995_, _11991_, _09453_);
  or _35924_ (_13513_, _11995_, _11993_);
  and _35925_ (_11996_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and _35926_ (_11997_, _11991_, _09463_);
  or _35927_ (_13514_, _11997_, _11996_);
  and _35928_ (_11998_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  and _35929_ (_11999_, _11991_, _09472_);
  or _35930_ (_13515_, _11999_, _11998_);
  and _35931_ (_12000_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and _35932_ (_12001_, _11991_, _09482_);
  or _35933_ (_13516_, _12001_, _12000_);
  and _35934_ (_12003_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and _35935_ (_12004_, _11991_, _09492_);
  or _35936_ (_13517_, _12004_, _12003_);
  and _35937_ (_12005_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and _35938_ (_12006_, _11991_, _09502_);
  or _35939_ (_13518_, _12006_, _12005_);
  and _35940_ (_12007_, _11989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and _35941_ (_12008_, _11991_, _09510_);
  or _35942_ (_13520_, _12008_, _12007_);
  not _35943_ (_12010_, _09659_);
  or _35944_ (_12011_, _11852_, _12010_);
  and _35945_ (_12012_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _35946_ (_12013_, _11875_, _09659_);
  and _35947_ (_12014_, _12013_, _09334_);
  or _35948_ (_13521_, _12014_, _12012_);
  and _35949_ (_12015_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and _35950_ (_12016_, _12013_, _09453_);
  or _35951_ (_13522_, _12016_, _12015_);
  and _35952_ (_12017_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and _35953_ (_12019_, _12013_, _09463_);
  or _35954_ (_13524_, _12019_, _12017_);
  and _35955_ (_12020_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _35956_ (_12021_, _12013_, _09472_);
  or _35957_ (_13525_, _12021_, _12020_);
  and _35958_ (_12022_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and _35959_ (_12023_, _12013_, _09482_);
  or _35960_ (_13526_, _12023_, _12022_);
  and _35961_ (_12024_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and _35962_ (_12025_, _12013_, _09492_);
  or _35963_ (_13527_, _12025_, _12024_);
  and _35964_ (_12027_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and _35965_ (_12028_, _12013_, _09502_);
  or _35966_ (_13528_, _12028_, _12027_);
  and _35967_ (_12029_, _12011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and _35968_ (_12030_, _12013_, _09510_);
  or _35969_ (_13529_, _12030_, _12029_);
  not _35970_ (_12031_, _09678_);
  or _35971_ (_12032_, _11852_, _12031_);
  and _35972_ (_12033_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  and _35973_ (_12035_, _11875_, _09678_);
  and _35974_ (_12036_, _12035_, _09334_);
  or _35975_ (_13530_, _12036_, _12033_);
  and _35976_ (_12037_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  and _35977_ (_12038_, _12035_, _09453_);
  or _35978_ (_13532_, _12038_, _12037_);
  and _35979_ (_12039_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  and _35980_ (_12040_, _12035_, _09463_);
  or _35981_ (_13533_, _12040_, _12039_);
  and _35982_ (_12041_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  and _35983_ (_12042_, _12035_, _09472_);
  or _35984_ (_13534_, _12042_, _12041_);
  and _35985_ (_12043_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and _35986_ (_12044_, _12035_, _09482_);
  or _35987_ (_13536_, _12044_, _12043_);
  and _35988_ (_12045_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  and _35989_ (_12046_, _12035_, _09492_);
  or _35990_ (_13537_, _12046_, _12045_);
  and _35991_ (_12047_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  and _35992_ (_12048_, _12035_, _09502_);
  or _35993_ (_13538_, _12048_, _12047_);
  and _35994_ (_12049_, _12032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and _35995_ (_12050_, _12035_, _09510_);
  or _35996_ (_13539_, _12050_, _12049_);
  not _35997_ (_12051_, _09697_);
  or _35998_ (_12052_, _11852_, _12051_);
  and _35999_ (_12053_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  and _36000_ (_12054_, _11875_, _09697_);
  and _36001_ (_12055_, _12054_, _09334_);
  or _36002_ (_13540_, _12055_, _12053_);
  and _36003_ (_12056_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and _36004_ (_12057_, _12054_, _09453_);
  or _36005_ (_13541_, _12057_, _12056_);
  and _36006_ (_12058_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and _36007_ (_12059_, _12054_, _09463_);
  or _36008_ (_13542_, _12059_, _12058_);
  and _36009_ (_12060_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and _36010_ (_12061_, _12054_, _09472_);
  or _36011_ (_13544_, _12061_, _12060_);
  and _36012_ (_12062_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and _36013_ (_12063_, _12054_, _09482_);
  or _36014_ (_13545_, _12063_, _12062_);
  and _36015_ (_12064_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  and _36016_ (_12065_, _12054_, _09492_);
  or _36017_ (_13546_, _12065_, _12064_);
  and _36018_ (_12066_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and _36019_ (_12067_, _12054_, _09502_);
  or _36020_ (_13548_, _12067_, _12066_);
  and _36021_ (_12068_, _12052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and _36022_ (_12069_, _12054_, _09510_);
  or _36023_ (_13549_, _12069_, _12068_);
  not _36024_ (_12070_, _09716_);
  or _36025_ (_12071_, _11852_, _12070_);
  and _36026_ (_12072_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _36027_ (_12073_, _11875_, _09716_);
  and _36028_ (_12074_, _12073_, _09334_);
  or _36029_ (_13550_, _12074_, _12072_);
  and _36030_ (_12075_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and _36031_ (_12076_, _12073_, _09453_);
  or _36032_ (_13552_, _12076_, _12075_);
  and _36033_ (_12077_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and _36034_ (_12078_, _12073_, _09463_);
  or _36035_ (_13553_, _12078_, _12077_);
  and _36036_ (_12079_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _36037_ (_12080_, _12073_, _09472_);
  or _36038_ (_13554_, _12080_, _12079_);
  and _36039_ (_12081_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and _36040_ (_12082_, _12073_, _09482_);
  or _36041_ (_13555_, _12082_, _12081_);
  and _36042_ (_12083_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _36043_ (_12084_, _12073_, _09492_);
  or _36044_ (_13557_, _12084_, _12083_);
  and _36045_ (_12085_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and _36046_ (_12086_, _12073_, _09502_);
  or _36047_ (_13558_, _12086_, _12085_);
  and _36048_ (_12087_, _12071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _36049_ (_12088_, _12073_, _09510_);
  or _36050_ (_13559_, _12088_, _12087_);
  not _36051_ (_12089_, _09736_);
  or _36052_ (_12090_, _11852_, _12089_);
  and _36053_ (_12091_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _36054_ (_12092_, _11875_, _09736_);
  and _36055_ (_12093_, _12092_, _09334_);
  or _36056_ (_13560_, _12093_, _12091_);
  and _36057_ (_12094_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and _36058_ (_12095_, _12092_, _09453_);
  or _36059_ (_13561_, _12095_, _12094_);
  and _36060_ (_12096_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _36061_ (_12097_, _12092_, _09463_);
  or _36062_ (_13562_, _12097_, _12096_);
  and _36063_ (_12098_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and _36064_ (_12099_, _12092_, _09472_);
  or _36065_ (_13564_, _12099_, _12098_);
  and _36066_ (_12100_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and _36067_ (_12101_, _12092_, _09482_);
  or _36068_ (_13565_, _12101_, _12100_);
  and _36069_ (_12102_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _36070_ (_12103_, _12092_, _09492_);
  or _36071_ (_13566_, _12103_, _12102_);
  and _36072_ (_12104_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and _36073_ (_12105_, _12092_, _09502_);
  or _36074_ (_13567_, _12105_, _12104_);
  and _36075_ (_12106_, _12090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and _36076_ (_12107_, _12092_, _09510_);
  or _36077_ (_13569_, _12107_, _12106_);
  not _36078_ (_12108_, _09755_);
  or _36079_ (_12109_, _11852_, _12108_);
  and _36080_ (_12110_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  and _36081_ (_12111_, _11875_, _09755_);
  and _36082_ (_12112_, _12111_, _09334_);
  or _36083_ (_13570_, _12112_, _12110_);
  and _36084_ (_12113_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and _36085_ (_12114_, _12111_, _09453_);
  or _36086_ (_13571_, _12114_, _12113_);
  and _36087_ (_12115_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and _36088_ (_12116_, _12111_, _09463_);
  or _36089_ (_13572_, _12116_, _12115_);
  and _36090_ (_12117_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  and _36091_ (_12118_, _12111_, _09472_);
  or _36092_ (_13573_, _12118_, _12117_);
  and _36093_ (_12119_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and _36094_ (_12120_, _12111_, _09482_);
  or _36095_ (_13574_, _12120_, _12119_);
  and _36096_ (_12121_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and _36097_ (_12122_, _12111_, _09492_);
  or _36098_ (_13576_, _12122_, _12121_);
  and _36099_ (_12123_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  and _36100_ (_12124_, _12111_, _09502_);
  or _36101_ (_13577_, _12124_, _12123_);
  and _36102_ (_12125_, _12109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and _36103_ (_12126_, _12111_, _09510_);
  or _36104_ (_13578_, _12126_, _12125_);
  not _36105_ (_12127_, _09774_);
  or _36106_ (_12128_, _11852_, _12127_);
  and _36107_ (_12129_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  and _36108_ (_12130_, _11875_, _09774_);
  and _36109_ (_12131_, _12130_, _09334_);
  or _36110_ (_13579_, _12131_, _12129_);
  and _36111_ (_12132_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and _36112_ (_12133_, _12130_, _09453_);
  or _36113_ (_13581_, _12133_, _12132_);
  and _36114_ (_12134_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and _36115_ (_12135_, _12130_, _09463_);
  or _36116_ (_13582_, _12135_, _12134_);
  and _36117_ (_12136_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and _36118_ (_12137_, _12130_, _09472_);
  or _36119_ (_13583_, _12137_, _12136_);
  and _36120_ (_12138_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  and _36121_ (_12139_, _12130_, _09482_);
  or _36122_ (_13584_, _12139_, _12138_);
  and _36123_ (_12140_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  and _36124_ (_12141_, _12130_, _09492_);
  or _36125_ (_13585_, _12141_, _12140_);
  and _36126_ (_12142_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  and _36127_ (_12143_, _12130_, _09502_);
  or _36128_ (_13586_, _12143_, _12142_);
  and _36129_ (_12144_, _12128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and _36130_ (_12145_, _12130_, _09510_);
  or _36131_ (_13587_, _12145_, _12144_);
  not _36132_ (_12146_, _09793_);
  or _36133_ (_12147_, _11852_, _12146_);
  and _36134_ (_12148_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _36135_ (_12149_, _11875_, _09793_);
  and _36136_ (_12150_, _12149_, _09334_);
  or _36137_ (_13589_, _12150_, _12148_);
  and _36138_ (_12151_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and _36139_ (_12152_, _12149_, _09453_);
  or _36140_ (_13590_, _12152_, _12151_);
  and _36141_ (_12153_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and _36142_ (_12154_, _12149_, _09463_);
  or _36143_ (_13591_, _12154_, _12153_);
  and _36144_ (_12155_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _36145_ (_12156_, _12149_, _09472_);
  or _36146_ (_13593_, _12156_, _12155_);
  and _36147_ (_12157_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and _36148_ (_12158_, _12149_, _09482_);
  or _36149_ (_13594_, _12158_, _12157_);
  and _36150_ (_12159_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _36151_ (_12160_, _12149_, _09492_);
  or _36152_ (_13595_, _12160_, _12159_);
  and _36153_ (_12161_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and _36154_ (_12162_, _12149_, _09502_);
  or _36155_ (_13596_, _12162_, _12161_);
  and _36156_ (_12163_, _12147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and _36157_ (_12164_, _12149_, _09510_);
  or _36158_ (_13597_, _12164_, _12163_);
  and _36159_ (_12165_, _09813_, _02161_);
  and _36160_ (_12166_, _12165_, _09265_);
  and _36161_ (_12167_, _12166_, _09513_);
  not _36162_ (_12168_, _12166_);
  and _36163_ (_12169_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or _36164_ (_13598_, _12169_, _12167_);
  and _36165_ (_12170_, _12166_, _09520_);
  and _36166_ (_12171_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  or _36167_ (_13600_, _12171_, _12170_);
  and _36168_ (_12172_, _12166_, _09523_);
  and _36169_ (_12173_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  or _36170_ (_13601_, _12173_, _12172_);
  and _36171_ (_12174_, _12166_, _09526_);
  and _36172_ (_12175_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  or _36173_ (_13602_, _12175_, _12174_);
  and _36174_ (_12176_, _12166_, _09529_);
  and _36175_ (_12177_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  or _36176_ (_13604_, _12177_, _12176_);
  and _36177_ (_12178_, _12166_, _09532_);
  and _36178_ (_12179_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or _36179_ (_13605_, _12179_, _12178_);
  and _36180_ (_12180_, _12166_, _09535_);
  and _36181_ (_12181_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  or _36182_ (_13606_, _12181_, _12180_);
  and _36183_ (_12182_, _12166_, _09538_);
  and _36184_ (_12183_, _12168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or _36185_ (_13607_, _12183_, _12182_);
  and _36186_ (_12184_, _12165_, _09515_);
  and _36187_ (_12185_, _12184_, _09513_);
  not _36188_ (_12186_, _12184_);
  and _36189_ (_12187_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _36190_ (_13608_, _12187_, _12185_);
  and _36191_ (_12188_, _12184_, _09520_);
  and _36192_ (_12189_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _36193_ (_13609_, _12189_, _12188_);
  and _36194_ (_12190_, _12184_, _09523_);
  and _36195_ (_12191_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _36196_ (_13610_, _12191_, _12190_);
  and _36197_ (_12192_, _12184_, _09526_);
  and _36198_ (_12193_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _36199_ (_13612_, _12193_, _12192_);
  and _36200_ (_12194_, _12184_, _09529_);
  and _36201_ (_12195_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _36202_ (_13613_, _12195_, _12194_);
  and _36203_ (_12196_, _12184_, _09532_);
  and _36204_ (_12197_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _36205_ (_13614_, _12197_, _12196_);
  and _36206_ (_12198_, _12184_, _09535_);
  and _36207_ (_12199_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _36208_ (_13616_, _12199_, _12198_);
  and _36209_ (_12200_, _12184_, _09538_);
  and _36210_ (_12201_, _12186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _36211_ (_13617_, _12201_, _12200_);
  and _36212_ (_12203_, _12165_, _09542_);
  and _36213_ (_12206_, _12203_, _09513_);
  not _36214_ (_12209_, _12203_);
  and _36215_ (_12212_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _36216_ (_13618_, _12212_, _12206_);
  and _36217_ (_12218_, _12203_, _09520_);
  and _36218_ (_12223_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _36219_ (_13619_, _12223_, _12218_);
  and _36220_ (_12229_, _12203_, _09523_);
  and _36221_ (_12233_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _36222_ (_13620_, _12233_, _12229_);
  and _36223_ (_12240_, _12203_, _09526_);
  and _36224_ (_12243_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _36225_ (_13621_, _12243_, _12240_);
  and _36226_ (_12251_, _12203_, _09529_);
  and _36227_ (_12255_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _36228_ (_13622_, _12255_, _12251_);
  and _36229_ (_12262_, _12203_, _09532_);
  and _36230_ (_12267_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _36231_ (_13624_, _12267_, _12262_);
  and _36232_ (_12274_, _12203_, _09535_);
  and _36233_ (_12278_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _36234_ (_13625_, _12278_, _12274_);
  and _36235_ (_12285_, _12203_, _09538_);
  and _36236_ (_12289_, _12209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _36237_ (_13626_, _12289_, _12285_);
  and _36238_ (_12296_, _12165_, _09562_);
  and _36239_ (_12301_, _12296_, _09513_);
  not _36240_ (_12305_, _12296_);
  and _36241_ (_12309_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or _36242_ (_13628_, _12309_, _12301_);
  and _36243_ (_12316_, _12296_, _09520_);
  and _36244_ (_12321_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  or _36245_ (_13629_, _12321_, _12316_);
  and _36246_ (_12328_, _12296_, _09523_);
  and _36247_ (_12332_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  or _36248_ (_13630_, _12332_, _12328_);
  and _36249_ (_12340_, _12296_, _09526_);
  and _36250_ (_12343_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  or _36251_ (_13631_, _12343_, _12340_);
  and _36252_ (_12351_, _12296_, _09529_);
  and _36253_ (_12355_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or _36254_ (_13632_, _12355_, _12351_);
  and _36255_ (_12361_, _12296_, _09532_);
  and _36256_ (_12366_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or _36257_ (_13633_, _12366_, _12361_);
  and _36258_ (_12373_, _12296_, _09535_);
  and _36259_ (_12378_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or _36260_ (_13634_, _12378_, _12373_);
  and _36261_ (_12385_, _12296_, _09538_);
  and _36262_ (_12390_, _12305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  or _36263_ (_13636_, _12390_, _12385_);
  and _36264_ (_12398_, _12165_, _09582_);
  and _36265_ (_12402_, _12398_, _09513_);
  not _36266_ (_12406_, _12398_);
  and _36267_ (_12410_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  or _36268_ (_13637_, _12410_, _12402_);
  and _36269_ (_12418_, _12398_, _09520_);
  and _36270_ (_12422_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or _36271_ (_13638_, _12422_, _12418_);
  and _36272_ (_12430_, _12398_, _09523_);
  and _36273_ (_12434_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or _36274_ (_13640_, _12434_, _12430_);
  and _36275_ (_12442_, _12398_, _09526_);
  and _36276_ (_12447_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or _36277_ (_13641_, _12447_, _12442_);
  and _36278_ (_12454_, _12398_, _09529_);
  and _36279_ (_12458_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  or _36280_ (_13642_, _12458_, _12454_);
  and _36281_ (_12466_, _12398_, _09532_);
  and _36282_ (_12470_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or _36283_ (_13643_, _12470_, _12466_);
  and _36284_ (_12478_, _12398_, _09535_);
  and _36285_ (_12482_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  or _36286_ (_13644_, _12482_, _12478_);
  and _36287_ (_12490_, _12398_, _09538_);
  and _36288_ (_12495_, _12406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or _36289_ (_13645_, _12495_, _12490_);
  and _36290_ (_12502_, _12165_, _09601_);
  and _36291_ (_12506_, _12502_, _09513_);
  not _36292_ (_12511_, _12502_);
  and _36293_ (_12515_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _36294_ (_13646_, _12515_, _12506_);
  and _36295_ (_12521_, _12502_, _09520_);
  and _36296_ (_12526_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _36297_ (_13648_, _12526_, _12521_);
  and _36298_ (_12534_, _12502_, _09523_);
  and _36299_ (_12538_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _36300_ (_13649_, _12538_, _12534_);
  and _36301_ (_12545_, _12502_, _09526_);
  and _36302_ (_12550_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _36303_ (_13650_, _12550_, _12545_);
  and _36304_ (_12557_, _12502_, _09529_);
  and _36305_ (_12562_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _36306_ (_13652_, _12562_, _12557_);
  and _36307_ (_12569_, _12502_, _09532_);
  and _36308_ (_12574_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _36309_ (_13653_, _12574_, _12569_);
  and _36310_ (_12582_, _12502_, _09535_);
  and _36311_ (_12586_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _36312_ (_13654_, _12586_, _12582_);
  and _36313_ (_12593_, _12502_, _09538_);
  and _36314_ (_12598_, _12511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _36315_ (_13655_, _12598_, _12593_);
  and _36316_ (_12605_, _12165_, _09620_);
  and _36317_ (_12610_, _12605_, _09513_);
  not _36318_ (_12614_, _12605_);
  and _36319_ (_12618_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _36320_ (_13657_, _12618_, _12610_);
  and _36321_ (_12626_, _12605_, _09520_);
  and _36322_ (_12631_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _36323_ (_13658_, _12631_, _12626_);
  and _36324_ (_12638_, _12605_, _09523_);
  and _36325_ (_12642_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _36326_ (_13659_, _12642_, _12638_);
  and _36327_ (_12650_, _12605_, _09526_);
  and _36328_ (_12654_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _36329_ (_13661_, _12654_, _12650_);
  and _36330_ (_12662_, _12605_, _09529_);
  and _36331_ (_12666_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _36332_ (_13662_, _12666_, _12662_);
  and _36333_ (_12673_, _12605_, _09532_);
  and _36334_ (_12678_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _36335_ (_13663_, _12678_, _12673_);
  and _36336_ (_12685_, _12605_, _09535_);
  and _36337_ (_12690_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _36338_ (_13665_, _12690_, _12685_);
  and _36339_ (_12698_, _12605_, _09538_);
  and _36340_ (_12702_, _12614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _36341_ (_13666_, _12702_, _12698_);
  and _36342_ (_12709_, _12165_, _09639_);
  and _36343_ (_12714_, _12709_, _09513_);
  not _36344_ (_12718_, _12709_);
  and _36345_ (_12722_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or _36346_ (_13667_, _12722_, _12714_);
  and _36347_ (_12730_, _12709_, _09520_);
  and _36348_ (_12734_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or _36349_ (_13668_, _12734_, _12730_);
  and _36350_ (_12742_, _12709_, _09523_);
  and _36351_ (_12747_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or _36352_ (_13669_, _12747_, _12742_);
  and _36353_ (_12754_, _12709_, _09526_);
  and _36354_ (_12758_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  or _36355_ (_13670_, _12758_, _12754_);
  and _36356_ (_12766_, _12709_, _09529_);
  and _36357_ (_12770_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  or _36358_ (_13671_, _12770_, _12766_);
  and _36359_ (_12778_, _12709_, _09532_);
  and _36360_ (_12782_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  or _36361_ (_13673_, _12782_, _12778_);
  and _36362_ (_12790_, _12709_, _09535_);
  and _36363_ (_12795_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or _36364_ (_13674_, _12795_, _12790_);
  and _36365_ (_12802_, _12709_, _09538_);
  and _36366_ (_12806_, _12718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or _36367_ (_13675_, _12806_, _12802_);
  and _36368_ (_12814_, _12165_, _09659_);
  and _36369_ (_12818_, _12814_, _09513_);
  not _36370_ (_12823_, _12814_);
  and _36371_ (_12826_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _36372_ (_13677_, _12826_, _12818_);
  and _36373_ (_12834_, _12814_, _09520_);
  and _36374_ (_12838_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _36375_ (_13678_, _12838_, _12834_);
  and _36376_ (_12845_, _12814_, _09523_);
  and _36377_ (_12850_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _36378_ (_13679_, _12850_, _12845_);
  and _36379_ (_12857_, _12814_, _09526_);
  and _36380_ (_12862_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _36381_ (_13680_, _12862_, _12857_);
  and _36382_ (_12869_, _12814_, _09529_);
  and _36383_ (_12874_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _36384_ (_13681_, _12874_, _12869_);
  and _36385_ (_12882_, _12814_, _09532_);
  and _36386_ (_12886_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _36387_ (_13682_, _12886_, _12882_);
  and _36388_ (_12893_, _12814_, _09535_);
  and _36389_ (_12898_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _36390_ (_13683_, _12898_, _12893_);
  and _36391_ (_12905_, _12814_, _09538_);
  and _36392_ (_12910_, _12823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _36393_ (_13685_, _12910_, _12905_);
  and _36394_ (_12917_, _12165_, _09678_);
  and _36395_ (_12922_, _12917_, _09513_);
  not _36396_ (_12926_, _12917_);
  and _36397_ (_12931_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  or _36398_ (_13686_, _12931_, _12922_);
  and _36399_ (_12938_, _12917_, _09520_);
  and _36400_ (_12942_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  or _36401_ (_13687_, _12942_, _12938_);
  and _36402_ (_12950_, _12917_, _09523_);
  and _36403_ (_12954_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  or _36404_ (_13689_, _12954_, _12950_);
  and _36405_ (_12962_, _12917_, _09526_);
  and _36406_ (_12966_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  or _36407_ (_13690_, _12966_, _12962_);
  and _36408_ (_12974_, _12917_, _09529_);
  and _36409_ (_12979_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or _36410_ (_13691_, _12979_, _12974_);
  and _36411_ (_12986_, _12917_, _09532_);
  and _36412_ (_12990_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  or _36413_ (_13692_, _12990_, _12986_);
  and _36414_ (_12998_, _12917_, _09535_);
  and _36415_ (_13002_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  or _36416_ (_13693_, _13002_, _12998_);
  and _36417_ (_13010_, _12917_, _09538_);
  and _36418_ (_13014_, _12926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or _36419_ (_13694_, _13014_, _13010_);
  and _36420_ (_13022_, _12165_, _09697_);
  and _36421_ (_13026_, _13022_, _09513_);
  not _36422_ (_13030_, _13022_);
  and _36423_ (_13035_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or _36424_ (_13695_, _13035_, _13026_);
  and _36425_ (_13042_, _13022_, _09520_);
  and _36426_ (_13047_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or _36427_ (_13697_, _13047_, _13042_);
  and _36428_ (_13054_, _13022_, _09523_);
  and _36429_ (_13059_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or _36430_ (_13698_, _13059_, _13054_);
  and _36431_ (_13066_, _13022_, _09526_);
  and _36432_ (_13071_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or _36433_ (_13699_, _13071_, _13066_);
  and _36434_ (_13078_, _13022_, _09529_);
  and _36435_ (_13083_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  or _36436_ (_13701_, _13083_, _13078_);
  and _36437_ (_13090_, _13022_, _09532_);
  and _36438_ (_13095_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or _36439_ (_13702_, _13095_, _13090_);
  and _36440_ (_13102_, _13022_, _09535_);
  and _36441_ (_13107_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or _36442_ (_13703_, _13107_, _13102_);
  and _36443_ (_13114_, _13022_, _09538_);
  and _36444_ (_13119_, _13030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  or _36445_ (_13704_, _13119_, _13114_);
  and _36446_ (_13126_, _12165_, _09716_);
  and _36447_ (_13131_, _13126_, _09513_);
  not _36448_ (_13135_, _13126_);
  and _36449_ (_13139_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _36450_ (_13705_, _13139_, _13131_);
  and _36451_ (_13147_, _13126_, _09520_);
  and _36452_ (_13151_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _36453_ (_13706_, _13151_, _13147_);
  and _36454_ (_13159_, _13126_, _09523_);
  and _36455_ (_13163_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _36456_ (_13707_, _13163_, _13159_);
  and _36457_ (_13171_, _13126_, _09526_);
  and _36458_ (_13175_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _36459_ (_13709_, _13175_, _13171_);
  and _36460_ (_13183_, _13126_, _09529_);
  and _36461_ (_13187_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _36462_ (_13710_, _13187_, _13183_);
  and _36463_ (_13195_, _13126_, _09532_);
  and _36464_ (_13199_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _36465_ (_13711_, _13199_, _13195_);
  and _36466_ (_13207_, _13126_, _09535_);
  and _36467_ (_13211_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _36468_ (_13713_, _13211_, _13207_);
  and _36469_ (_13219_, _13126_, _09538_);
  and _36470_ (_13223_, _13135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _36471_ (_13714_, _13223_, _13219_);
  and _36472_ (_13231_, _12165_, _09736_);
  and _36473_ (_13235_, _13231_, _09513_);
  not _36474_ (_13240_, _13231_);
  and _36475_ (_13244_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _36476_ (_13715_, _13244_, _13235_);
  and _36477_ (_13251_, _13231_, _09520_);
  and _36478_ (_13256_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _36479_ (_13716_, _13256_, _13251_);
  and _36480_ (_13263_, _13231_, _09523_);
  and _36481_ (_13268_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _36482_ (_13717_, _13268_, _13263_);
  and _36483_ (_13275_, _13231_, _09526_);
  and _36484_ (_13280_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _36485_ (_13718_, _13280_, _13275_);
  and _36486_ (_13288_, _13231_, _09529_);
  and _36487_ (_13291_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _36488_ (_13719_, _13291_, _13288_);
  and _36489_ (_13299_, _13231_, _09532_);
  and _36490_ (_13303_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _36491_ (_13721_, _13303_, _13299_);
  and _36492_ (_13311_, _13231_, _09535_);
  and _36493_ (_13315_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _36494_ (_13722_, _13315_, _13311_);
  and _36495_ (_13323_, _13231_, _09538_);
  and _36496_ (_13327_, _13240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _36497_ (_13723_, _13327_, _13323_);
  and _36498_ (_13335_, _12165_, _09755_);
  and _36499_ (_13339_, _13335_, _09513_);
  not _36500_ (_13344_, _13335_);
  and _36501_ (_13348_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or _36502_ (_13725_, _13348_, _13339_);
  and _36503_ (_13356_, _13335_, _09520_);
  and _36504_ (_13360_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  or _36505_ (_13726_, _13360_, _13356_);
  and _36506_ (_13368_, _13335_, _09523_);
  and _36507_ (_13372_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or _36508_ (_13727_, _13372_, _13368_);
  and _36509_ (_13380_, _13335_, _09526_);
  and _36510_ (_13384_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or _36511_ (_13728_, _13384_, _13380_);
  and _36512_ (_13392_, _13335_, _09529_);
  and _36513_ (_13396_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or _36514_ (_13729_, _13396_, _13392_);
  and _36515_ (_13404_, _13335_, _09532_);
  and _36516_ (_13408_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  or _36517_ (_13730_, _13408_, _13404_);
  and _36518_ (_13416_, _13335_, _09535_);
  and _36519_ (_13420_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  or _36520_ (_13731_, _13420_, _13416_);
  and _36521_ (_13428_, _13335_, _09538_);
  and _36522_ (_13432_, _13344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  or _36523_ (_13733_, _13432_, _13428_);
  and _36524_ (_13440_, _12165_, _09774_);
  and _36525_ (_13443_, _13440_, _09513_);
  not _36526_ (_13447_, _13440_);
  and _36527_ (_13451_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  or _36528_ (_13734_, _13451_, _13443_);
  and _36529_ (_13459_, _13440_, _09520_);
  and _36530_ (_13463_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or _36531_ (_13735_, _13463_, _13459_);
  and _36532_ (_13471_, _13440_, _09523_);
  and _36533_ (_13475_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  or _36534_ (_13737_, _13475_, _13471_);
  and _36535_ (_13483_, _13440_, _09526_);
  and _36536_ (_13487_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  or _36537_ (_13738_, _13487_, _13483_);
  and _36538_ (_13495_, _13440_, _09529_);
  and _36539_ (_13499_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  or _36540_ (_13739_, _13499_, _13495_);
  and _36541_ (_13507_, _13440_, _09532_);
  and _36542_ (_13511_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or _36543_ (_13740_, _13511_, _13507_);
  and _36544_ (_13519_, _13440_, _09535_);
  and _36545_ (_13523_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or _36546_ (_13741_, _13523_, _13519_);
  and _36547_ (_13531_, _13440_, _09538_);
  and _36548_ (_13535_, _13447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or _36549_ (_13742_, _13535_, _13531_);
  and _36550_ (_13543_, _12165_, _09793_);
  and _36551_ (_13547_, _13543_, _09513_);
  not _36552_ (_13551_, _13543_);
  and _36553_ (_13556_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _36554_ (_13743_, _13556_, _13547_);
  and _36555_ (_13563_, _13543_, _09520_);
  and _36556_ (_13568_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _36557_ (_13745_, _13568_, _13563_);
  and _36558_ (_13575_, _13543_, _09523_);
  and _36559_ (_13580_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _36560_ (_13746_, _13580_, _13575_);
  and _36561_ (_13588_, _13543_, _09526_);
  and _36562_ (_13592_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _36563_ (_13747_, _13592_, _13588_);
  and _36564_ (_13599_, _13543_, _09529_);
  and _36565_ (_13603_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _36566_ (_13749_, _13603_, _13599_);
  and _36567_ (_13611_, _13543_, _09532_);
  and _36568_ (_13615_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _36569_ (_13750_, _13615_, _13611_);
  and _36570_ (_13623_, _13543_, _09535_);
  and _36571_ (_13627_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _36572_ (_13751_, _13627_, _13623_);
  and _36573_ (_13635_, _13543_, _09538_);
  and _36574_ (_13639_, _13551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _36575_ (_13752_, _13639_, _13635_);
  and _36576_ (_13647_, _10103_, _02161_);
  and _36577_ (_13651_, _13647_, _09265_);
  and _36578_ (_13656_, _13651_, _09513_);
  not _36579_ (_13660_, _13651_);
  and _36580_ (_13664_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _36581_ (_13753_, _13664_, _13656_);
  and _36582_ (_13672_, _13651_, _09520_);
  and _36583_ (_13676_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or _36584_ (_13754_, _13676_, _13672_);
  and _36585_ (_13684_, _13651_, _09523_);
  and _36586_ (_13688_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _36587_ (_13755_, _13688_, _13684_);
  and _36588_ (_13696_, _13651_, _09526_);
  and _36589_ (_13700_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _36590_ (_13757_, _13700_, _13696_);
  and _36591_ (_13708_, _13651_, _09529_);
  and _36592_ (_13712_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or _36593_ (_13758_, _13712_, _13708_);
  and _36594_ (_13720_, _13651_, _09532_);
  and _36595_ (_13724_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _36596_ (_13759_, _13724_, _13720_);
  and _36597_ (_13732_, _13651_, _09535_);
  and _36598_ (_13736_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _36599_ (_13761_, _13736_, _13732_);
  and _36600_ (_13744_, _13651_, _09538_);
  and _36601_ (_13748_, _13660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _36602_ (_13762_, _13748_, _13744_);
  and _36603_ (_13756_, _13647_, _09515_);
  and _36604_ (_13760_, _13756_, _09513_);
  not _36605_ (_13764_, _13756_);
  and _36606_ (_13769_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  or _36607_ (_13763_, _13769_, _13760_);
  and _36608_ (_13776_, _13756_, _09520_);
  and _36609_ (_13781_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  or _36610_ (_13765_, _13781_, _13776_);
  and _36611_ (_13788_, _13756_, _09523_);
  and _36612_ (_13793_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  or _36613_ (_13766_, _13793_, _13788_);
  and _36614_ (_13801_, _13756_, _09526_);
  and _36615_ (_13805_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  or _36616_ (_13767_, _13805_, _13801_);
  and _36617_ (_13812_, _13756_, _09529_);
  and _36618_ (_13817_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  or _36619_ (_13768_, _13817_, _13812_);
  and _36620_ (_13824_, _13756_, _09532_);
  and _36621_ (_13829_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  or _36622_ (_13770_, _13829_, _13824_);
  and _36623_ (_13836_, _13756_, _09535_);
  and _36624_ (_13841_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  or _36625_ (_13771_, _13841_, _13836_);
  and _36626_ (_13849_, _13756_, _09538_);
  and _36627_ (_13853_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  or _36628_ (_13772_, _13853_, _13849_);
  and _36629_ (_13860_, _13647_, _09542_);
  and _36630_ (_13865_, _13860_, _09513_);
  not _36631_ (_13869_, _13860_);
  and _36632_ (_13873_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  or _36633_ (_13773_, _13873_, _13865_);
  and _36634_ (_13881_, _13860_, _09520_);
  and _36635_ (_13885_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  or _36636_ (_13774_, _13885_, _13881_);
  and _36637_ (_13893_, _13860_, _09523_);
  and _36638_ (_13898_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  or _36639_ (_13775_, _13898_, _13893_);
  and _36640_ (_13905_, _13860_, _09526_);
  and _36641_ (_13909_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  or _36642_ (_13777_, _13909_, _13905_);
  and _36643_ (_13917_, _13860_, _09529_);
  and _36644_ (_13921_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  or _36645_ (_13778_, _13921_, _13917_);
  and _36646_ (_13929_, _13860_, _09532_);
  and _36647_ (_13933_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  or _36648_ (_13779_, _13933_, _13929_);
  and _36649_ (_13941_, _13860_, _09535_);
  and _36650_ (_13945_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  or _36651_ (_13780_, _13945_, _13941_);
  and _36652_ (_13953_, _13860_, _09538_);
  and _36653_ (_13957_, _13869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  or _36654_ (_13782_, _13957_, _13953_);
  and _36655_ (_13965_, _13647_, _09562_);
  and _36656_ (_13969_, _13965_, _09513_);
  not _36657_ (_13973_, _13965_);
  and _36658_ (_13978_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _36659_ (_13783_, _13978_, _13969_);
  and _36660_ (_13985_, _13965_, _09520_);
  and _36661_ (_13990_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or _36662_ (_13784_, _13990_, _13985_);
  and _36663_ (_13997_, _13965_, _09523_);
  and _36664_ (_14002_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _36665_ (_13785_, _14002_, _13997_);
  and _36666_ (_14009_, _13965_, _09526_);
  and _36667_ (_14014_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or _36668_ (_13786_, _14014_, _14009_);
  and _36669_ (_14021_, _13965_, _09529_);
  and _36670_ (_14026_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or _36671_ (_13787_, _14026_, _14021_);
  and _36672_ (_14033_, _13965_, _09532_);
  and _36673_ (_14038_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or _36674_ (_13789_, _14038_, _14033_);
  and _36675_ (_14045_, _13965_, _09535_);
  and _36676_ (_14050_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or _36677_ (_13790_, _14050_, _14045_);
  and _36678_ (_14057_, _13965_, _09538_);
  and _36679_ (_14062_, _13973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _36680_ (_13791_, _14062_, _14057_);
  and _36681_ (_14069_, _13647_, _09582_);
  and _36682_ (_14073_, _14069_, _09513_);
  not _36683_ (_14077_, _14069_);
  and _36684_ (_14082_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or _36685_ (_13792_, _14082_, _14073_);
  and _36686_ (_14089_, _14069_, _09520_);
  and _36687_ (_14094_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _36688_ (_13794_, _14094_, _14089_);
  and _36689_ (_14101_, _14069_, _09523_);
  and _36690_ (_14106_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or _36691_ (_13795_, _14106_, _14101_);
  and _36692_ (_14113_, _14069_, _09526_);
  and _36693_ (_14118_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _36694_ (_13796_, _14118_, _14113_);
  and _36695_ (_14125_, _14069_, _09529_);
  and _36696_ (_14130_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _36697_ (_13797_, _14130_, _14125_);
  and _36698_ (_14137_, _14069_, _09532_);
  and _36699_ (_14142_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _36700_ (_13798_, _14142_, _14137_);
  and _36701_ (_14149_, _14069_, _09535_);
  and _36702_ (_14154_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _36703_ (_13799_, _14154_, _14149_);
  and _36704_ (_14161_, _14069_, _09538_);
  and _36705_ (_14166_, _14077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _36706_ (_13800_, _14166_, _14161_);
  and _36707_ (_14173_, _13647_, _09601_);
  and _36708_ (_14178_, _14173_, _09513_);
  not _36709_ (_14182_, _14173_);
  and _36710_ (_14186_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  or _36711_ (_13802_, _14186_, _14178_);
  and _36712_ (_14194_, _14173_, _09520_);
  and _36713_ (_14198_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  or _36714_ (_13803_, _14198_, _14194_);
  and _36715_ (_14206_, _14173_, _09523_);
  and _36716_ (_14210_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  or _36717_ (_13804_, _14210_, _14206_);
  and _36718_ (_14218_, _14173_, _09526_);
  and _36719_ (_14222_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  or _36720_ (_13806_, _14222_, _14218_);
  and _36721_ (_14230_, _14173_, _09529_);
  and _36722_ (_14234_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  or _36723_ (_13807_, _14234_, _14230_);
  and _36724_ (_14242_, _14173_, _09532_);
  and _36725_ (_14246_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  or _36726_ (_13808_, _14246_, _14242_);
  and _36727_ (_14254_, _14173_, _09535_);
  and _36728_ (_14258_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  or _36729_ (_13809_, _14258_, _14254_);
  and _36730_ (_14266_, _14173_, _09538_);
  and _36731_ (_14270_, _14182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  or _36732_ (_13810_, _14270_, _14266_);
  and _36733_ (_14278_, _13647_, _09620_);
  and _36734_ (_14282_, _14278_, _09513_);
  not _36735_ (_14286_, _14278_);
  and _36736_ (_14291_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  or _36737_ (_13811_, _14291_, _14282_);
  and _36738_ (_14298_, _14278_, _09520_);
  and _36739_ (_14303_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  or _36740_ (_13813_, _14303_, _14298_);
  and _36741_ (_14310_, _14278_, _09523_);
  and _36742_ (_14315_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  or _36743_ (_13814_, _14315_, _14310_);
  and _36744_ (_14323_, _14278_, _09526_);
  and _36745_ (_14327_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  or _36746_ (_13815_, _14327_, _14323_);
  and _36747_ (_14334_, _14278_, _09529_);
  and _36748_ (_14339_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  or _36749_ (_13816_, _14339_, _14334_);
  and _36750_ (_14346_, _14278_, _09532_);
  and _36751_ (_14351_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  or _36752_ (_13818_, _14351_, _14346_);
  and _36753_ (_14358_, _14278_, _09535_);
  and _36754_ (_14363_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  or _36755_ (_13819_, _14363_, _14358_);
  and _36756_ (_14371_, _14278_, _09538_);
  and _36757_ (_14374_, _14286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  or _36758_ (_13820_, _14374_, _14371_);
  and _36759_ (_14382_, _13647_, _09639_);
  and _36760_ (_14386_, _14382_, _09513_);
  not _36761_ (_14391_, _14382_);
  and _36762_ (_14395_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _36763_ (_13821_, _14395_, _14386_);
  and _36764_ (_14403_, _14382_, _09520_);
  and _36765_ (_14407_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _36766_ (_13822_, _14407_, _14403_);
  and _36767_ (_14415_, _14382_, _09523_);
  and _36768_ (_14419_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _36769_ (_13823_, _14419_, _14415_);
  and _36770_ (_14427_, _14382_, _09526_);
  and _36771_ (_14431_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _36772_ (_13825_, _14431_, _14427_);
  and _36773_ (_14439_, _14382_, _09529_);
  and _36774_ (_14443_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or _36775_ (_13826_, _14443_, _14439_);
  and _36776_ (_14451_, _14382_, _09532_);
  and _36777_ (_14455_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _36778_ (_13827_, _14455_, _14451_);
  and _36779_ (_14463_, _14382_, _09535_);
  and _36780_ (_14467_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or _36781_ (_13828_, _14467_, _14463_);
  and _36782_ (_14475_, _14382_, _09538_);
  and _36783_ (_14479_, _14391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _36784_ (_13830_, _14479_, _14475_);
  and _36785_ (_14487_, _13647_, _09659_);
  and _36786_ (_14491_, _14487_, _09513_);
  not _36787_ (_14495_, _14487_);
  and _36788_ (_14500_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  or _36789_ (_13831_, _14500_, _14491_);
  and _36790_ (_14507_, _14487_, _09520_);
  and _36791_ (_14512_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  or _36792_ (_13832_, _14512_, _14507_);
  and _36793_ (_14519_, _14487_, _09523_);
  and _36794_ (_14524_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  or _36795_ (_13833_, _14524_, _14519_);
  and _36796_ (_14531_, _14487_, _09526_);
  and _36797_ (_14536_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  or _36798_ (_13834_, _14536_, _14531_);
  and _36799_ (_14543_, _14487_, _09529_);
  and _36800_ (_14547_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  or _36801_ (_13835_, _14547_, _14543_);
  and _36802_ (_14555_, _14487_, _09532_);
  and _36803_ (_14559_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  or _36804_ (_13837_, _14559_, _14555_);
  and _36805_ (_14567_, _14487_, _09535_);
  and _36806_ (_14571_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  or _36807_ (_13838_, _14571_, _14567_);
  and _36808_ (_14579_, _14487_, _09538_);
  and _36809_ (_14584_, _14495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  or _36810_ (_13839_, _14584_, _14579_);
  and _36811_ (_14591_, _13647_, _09678_);
  and _36812_ (_14595_, _14591_, _09513_);
  not _36813_ (_14600_, _14591_);
  and _36814_ (_14604_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _36815_ (_13840_, _14604_, _14595_);
  and _36816_ (_14612_, _14591_, _09520_);
  and _36817_ (_14616_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _36818_ (_13842_, _14616_, _14612_);
  and _36819_ (_14624_, _14591_, _09523_);
  and _36820_ (_14628_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _36821_ (_13843_, _14628_, _14624_);
  and _36822_ (_14636_, _14591_, _09526_);
  and _36823_ (_14640_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _36824_ (_13844_, _14640_, _14636_);
  and _36825_ (_14648_, _14591_, _09529_);
  and _36826_ (_14652_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _36827_ (_13845_, _14652_, _14648_);
  and _36828_ (_14660_, _14591_, _09532_);
  and _36829_ (_14664_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or _36830_ (_13846_, _14664_, _14660_);
  and _36831_ (_14672_, _14591_, _09535_);
  and _36832_ (_14676_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or _36833_ (_13847_, _14676_, _14672_);
  and _36834_ (_14682_, _14591_, _09538_);
  and _36835_ (_14686_, _14600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or _36836_ (_13848_, _14686_, _14682_);
  and _36837_ (_14690_, _13647_, _09697_);
  and _36838_ (_14691_, _14690_, _09513_);
  not _36839_ (_14692_, _14690_);
  and _36840_ (_14693_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or _36841_ (_13850_, _14693_, _14691_);
  and _36842_ (_14694_, _14690_, _09520_);
  and _36843_ (_14695_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or _36844_ (_13851_, _14695_, _14694_);
  and _36845_ (_14696_, _14690_, _09523_);
  and _36846_ (_14697_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or _36847_ (_13852_, _14697_, _14696_);
  and _36848_ (_14698_, _14690_, _09526_);
  and _36849_ (_14699_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or _36850_ (_13854_, _14699_, _14698_);
  and _36851_ (_14700_, _14690_, _09529_);
  and _36852_ (_14701_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or _36853_ (_13855_, _14701_, _14700_);
  and _36854_ (_14702_, _14690_, _09532_);
  and _36855_ (_14703_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _36856_ (_13856_, _14703_, _14702_);
  and _36857_ (_14704_, _14690_, _09535_);
  and _36858_ (_14705_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _36859_ (_13857_, _14705_, _14704_);
  and _36860_ (_14706_, _14690_, _09538_);
  and _36861_ (_14707_, _14692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _36862_ (_13858_, _14707_, _14706_);
  and _36863_ (_14708_, _13647_, _09716_);
  and _36864_ (_14709_, _14708_, _09513_);
  not _36865_ (_14710_, _14708_);
  and _36866_ (_14711_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  or _36867_ (_13859_, _14711_, _14709_);
  and _36868_ (_14712_, _14708_, _09520_);
  and _36869_ (_14713_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  or _36870_ (_13861_, _14713_, _14712_);
  and _36871_ (_14714_, _14708_, _09523_);
  and _36872_ (_14715_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  or _36873_ (_13862_, _14715_, _14714_);
  and _36874_ (_14716_, _14708_, _09526_);
  and _36875_ (_14717_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  or _36876_ (_13863_, _14717_, _14716_);
  and _36877_ (_14718_, _14708_, _09529_);
  and _36878_ (_14719_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  or _36879_ (_13864_, _14719_, _14718_);
  and _36880_ (_14720_, _14708_, _09532_);
  and _36881_ (_14721_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  or _36882_ (_13866_, _14721_, _14720_);
  and _36883_ (_14722_, _14708_, _09535_);
  and _36884_ (_14723_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  or _36885_ (_13867_, _14723_, _14722_);
  and _36886_ (_14724_, _14708_, _09538_);
  and _36887_ (_14725_, _14710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  or _36888_ (_13868_, _14725_, _14724_);
  and _36889_ (_14726_, _13647_, _09736_);
  and _36890_ (_14727_, _14726_, _09513_);
  not _36891_ (_14728_, _14726_);
  and _36892_ (_14729_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  or _36893_ (_13870_, _14729_, _14727_);
  and _36894_ (_14730_, _14726_, _09520_);
  and _36895_ (_14731_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  or _36896_ (_13871_, _14731_, _14730_);
  and _36897_ (_14732_, _14726_, _09523_);
  and _36898_ (_14733_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  or _36899_ (_13872_, _14733_, _14732_);
  and _36900_ (_14734_, _14726_, _09526_);
  and _36901_ (_14735_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  or _36902_ (_13874_, _14735_, _14734_);
  and _36903_ (_14736_, _14726_, _09529_);
  and _36904_ (_14737_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  or _36905_ (_13875_, _14737_, _14736_);
  and _36906_ (_14738_, _14726_, _09532_);
  and _36907_ (_14739_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  or _36908_ (_13876_, _14739_, _14738_);
  and _36909_ (_14740_, _14726_, _09535_);
  and _36910_ (_14741_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  or _36911_ (_13877_, _14741_, _14740_);
  and _36912_ (_14742_, _14726_, _09538_);
  and _36913_ (_14743_, _14728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  or _36914_ (_13878_, _14743_, _14742_);
  and _36915_ (_14744_, _13647_, _09755_);
  and _36916_ (_14745_, _14744_, _09513_);
  not _36917_ (_14746_, _14744_);
  and _36918_ (_14747_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or _36919_ (_13879_, _14747_, _14745_);
  and _36920_ (_14748_, _14744_, _09520_);
  and _36921_ (_14749_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _36922_ (_13880_, _14749_, _14748_);
  and _36923_ (_14750_, _14744_, _09523_);
  and _36924_ (_14751_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or _36925_ (_13882_, _14751_, _14750_);
  and _36926_ (_14752_, _14744_, _09526_);
  and _36927_ (_14753_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or _36928_ (_13883_, _14753_, _14752_);
  and _36929_ (_14754_, _14744_, _09529_);
  and _36930_ (_14755_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _36931_ (_13884_, _14755_, _14754_);
  and _36932_ (_14756_, _14744_, _09532_);
  and _36933_ (_14757_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or _36934_ (_13886_, _14757_, _14756_);
  and _36935_ (_14758_, _14744_, _09535_);
  and _36936_ (_14759_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or _36937_ (_13887_, _14759_, _14758_);
  and _36938_ (_14760_, _14744_, _09538_);
  and _36939_ (_14761_, _14746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _36940_ (_13888_, _14761_, _14760_);
  and _36941_ (_14762_, _13647_, _09774_);
  and _36942_ (_14763_, _14762_, _09513_);
  not _36943_ (_14764_, _14762_);
  and _36944_ (_14765_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _36945_ (_13889_, _14765_, _14763_);
  and _36946_ (_14766_, _14762_, _09520_);
  and _36947_ (_14767_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or _36948_ (_13890_, _14767_, _14766_);
  and _36949_ (_14768_, _14762_, _09523_);
  and _36950_ (_14769_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _36951_ (_13891_, _14769_, _14768_);
  and _36952_ (_14770_, _14762_, _09526_);
  and _36953_ (_14771_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _36954_ (_13892_, _14771_, _14770_);
  and _36955_ (_14772_, _14762_, _09529_);
  and _36956_ (_14773_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or _36957_ (_13894_, _14773_, _14772_);
  and _36958_ (_14774_, _14762_, _09532_);
  and _36959_ (_14775_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _36960_ (_13895_, _14775_, _14774_);
  and _36961_ (_14776_, _14762_, _09535_);
  and _36962_ (_14777_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _36963_ (_13896_, _14777_, _14776_);
  and _36964_ (_14778_, _14762_, _09538_);
  and _36965_ (_14779_, _14764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or _36966_ (_13897_, _14779_, _14778_);
  and _36967_ (_14780_, _13647_, _09793_);
  and _36968_ (_14781_, _14780_, _09513_);
  not _36969_ (_14782_, _14780_);
  and _36970_ (_14783_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  or _36971_ (_13899_, _14783_, _14781_);
  and _36972_ (_14784_, _14780_, _09520_);
  and _36973_ (_14785_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  or _36974_ (_13900_, _14785_, _14784_);
  and _36975_ (_14786_, _14780_, _09523_);
  and _36976_ (_14787_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  or _36977_ (_13901_, _14787_, _14786_);
  and _36978_ (_14788_, _14780_, _09526_);
  and _36979_ (_14789_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  or _36980_ (_13902_, _14789_, _14788_);
  and _36981_ (_14790_, _14780_, _09529_);
  and _36982_ (_14791_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  or _36983_ (_13903_, _14791_, _14790_);
  and _36984_ (_14792_, _14780_, _09532_);
  and _36985_ (_14793_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  or _36986_ (_13904_, _14793_, _14792_);
  and _36987_ (_14794_, _14780_, _09535_);
  and _36988_ (_14795_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  or _36989_ (_13906_, _14795_, _14794_);
  and _36990_ (_14796_, _14780_, _09538_);
  and _36991_ (_14797_, _14782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  or _36992_ (_13907_, _14797_, _14796_);
  and _36993_ (_14798_, _10393_, _02161_);
  and _36994_ (_14799_, _14798_, _09265_);
  and _36995_ (_14800_, _14799_, _09513_);
  not _36996_ (_14801_, _14799_);
  and _36997_ (_14802_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or _36998_ (_13908_, _14802_, _14800_);
  and _36999_ (_14810_, _14799_, _09520_);
  and _37000_ (_14811_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or _37001_ (_13910_, _14811_, _14810_);
  and _37002_ (_14812_, _14799_, _09523_);
  and _37003_ (_14813_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or _37004_ (_13911_, _14813_, _14812_);
  and _37005_ (_14814_, _14799_, _09526_);
  and _37006_ (_14815_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or _37007_ (_13912_, _14815_, _14814_);
  and _37008_ (_14816_, _14799_, _09529_);
  and _37009_ (_14817_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or _37010_ (_13913_, _14817_, _14816_);
  and _37011_ (_14818_, _14799_, _09532_);
  and _37012_ (_14819_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or _37013_ (_13914_, _14819_, _14818_);
  and _37014_ (_14820_, _14799_, _09535_);
  and _37015_ (_14821_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or _37016_ (_13915_, _14821_, _14820_);
  and _37017_ (_14822_, _14799_, _09538_);
  and _37018_ (_14823_, _14801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or _37019_ (_13916_, _14823_, _14822_);
  and _37020_ (_14824_, _14798_, _09515_);
  and _37021_ (_14825_, _14824_, _09513_);
  not _37022_ (_14826_, _14824_);
  and _37023_ (_14827_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _37024_ (_13918_, _14827_, _14825_);
  and _37025_ (_14828_, _14824_, _09520_);
  and _37026_ (_14829_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _37027_ (_13919_, _14829_, _14828_);
  and _37028_ (_14830_, _14824_, _09523_);
  and _37029_ (_14831_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _37030_ (_13920_, _14831_, _14830_);
  and _37031_ (_14832_, _14824_, _09526_);
  and _37032_ (_14833_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _37033_ (_13922_, _14833_, _14832_);
  and _37034_ (_14834_, _14824_, _09529_);
  and _37035_ (_14835_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _37036_ (_13923_, _14835_, _14834_);
  and _37037_ (_14836_, _14824_, _09532_);
  and _37038_ (_14837_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _37039_ (_13924_, _14837_, _14836_);
  and _37040_ (_14838_, _14824_, _09535_);
  and _37041_ (_14839_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _37042_ (_13925_, _14839_, _14838_);
  and _37043_ (_14840_, _14824_, _09538_);
  and _37044_ (_14841_, _14826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _37045_ (_13926_, _14841_, _14840_);
  and _37046_ (_14842_, _14798_, _09542_);
  and _37047_ (_14843_, _14842_, _09513_);
  not _37048_ (_14844_, _14842_);
  and _37049_ (_14845_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _37050_ (_13927_, _14845_, _14843_);
  and _37051_ (_14846_, _14842_, _09520_);
  and _37052_ (_14847_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _37053_ (_13928_, _14847_, _14846_);
  and _37054_ (_14848_, _14842_, _09523_);
  and _37055_ (_14849_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _37056_ (_13930_, _14849_, _14848_);
  and _37057_ (_14850_, _14842_, _09526_);
  and _37058_ (_14851_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _37059_ (_13931_, _14851_, _14850_);
  and _37060_ (_14852_, _14842_, _09529_);
  and _37061_ (_14853_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _37062_ (_13932_, _14853_, _14852_);
  and _37063_ (_14854_, _14842_, _09532_);
  and _37064_ (_14855_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _37065_ (_13934_, _14855_, _14854_);
  and _37066_ (_14856_, _14842_, _09535_);
  and _37067_ (_14857_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _37068_ (_13935_, _14857_, _14856_);
  and _37069_ (_14858_, _14842_, _09538_);
  and _37070_ (_14859_, _14844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _37071_ (_13936_, _14859_, _14858_);
  and _37072_ (_14860_, _14798_, _09562_);
  and _37073_ (_14861_, _14860_, _09513_);
  not _37074_ (_14862_, _14860_);
  and _37075_ (_14863_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or _37076_ (_13937_, _14863_, _14861_);
  and _37077_ (_14864_, _14860_, _09520_);
  and _37078_ (_14865_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or _37079_ (_13938_, _14865_, _14864_);
  and _37080_ (_14866_, _14860_, _09523_);
  and _37081_ (_14867_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or _37082_ (_13939_, _14867_, _14866_);
  and _37083_ (_14868_, _14860_, _09526_);
  and _37084_ (_14869_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or _37085_ (_13940_, _14869_, _14868_);
  and _37086_ (_14870_, _14860_, _09529_);
  and _37087_ (_14871_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or _37088_ (_13942_, _14871_, _14870_);
  and _37089_ (_14872_, _14860_, _09532_);
  and _37090_ (_14873_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or _37091_ (_13943_, _14873_, _14872_);
  and _37092_ (_14874_, _14860_, _09535_);
  and _37093_ (_14875_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or _37094_ (_13944_, _14875_, _14874_);
  and _37095_ (_14876_, _14860_, _09538_);
  and _37096_ (_14877_, _14862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or _37097_ (_13946_, _14877_, _14876_);
  and _37098_ (_14878_, _14798_, _09582_);
  and _37099_ (_14879_, _14878_, _09513_);
  not _37100_ (_14880_, _14878_);
  and _37101_ (_14881_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or _37102_ (_13947_, _14881_, _14879_);
  and _37103_ (_14882_, _14878_, _09520_);
  and _37104_ (_14883_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or _37105_ (_13948_, _14883_, _14882_);
  and _37106_ (_14884_, _14878_, _09523_);
  and _37107_ (_14885_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or _37108_ (_13949_, _14885_, _14884_);
  and _37109_ (_14886_, _14878_, _09526_);
  and _37110_ (_14887_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or _37111_ (_13950_, _14887_, _14886_);
  and _37112_ (_14888_, _14878_, _09529_);
  and _37113_ (_14889_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or _37114_ (_13951_, _14889_, _14888_);
  and _37115_ (_14890_, _14878_, _09532_);
  and _37116_ (_14891_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or _37117_ (_13952_, _14891_, _14890_);
  and _37118_ (_14892_, _14878_, _09535_);
  and _37119_ (_14893_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or _37120_ (_13954_, _14893_, _14892_);
  and _37121_ (_14894_, _14878_, _09538_);
  and _37122_ (_14895_, _14880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or _37123_ (_13955_, _14895_, _14894_);
  and _37124_ (_14896_, _14798_, _09601_);
  and _37125_ (_14897_, _14896_, _09513_);
  not _37126_ (_14898_, _14896_);
  and _37127_ (_14899_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _37128_ (_13956_, _14899_, _14897_);
  and _37129_ (_14900_, _14896_, _09520_);
  and _37130_ (_14901_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _37131_ (_13958_, _14901_, _14900_);
  and _37132_ (_14902_, _14896_, _09523_);
  and _37133_ (_14903_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _37134_ (_13959_, _14903_, _14902_);
  and _37135_ (_14904_, _14896_, _09526_);
  and _37136_ (_14905_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _37137_ (_13960_, _14905_, _14904_);
  and _37138_ (_14906_, _14896_, _09529_);
  and _37139_ (_14907_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _37140_ (_13961_, _14907_, _14906_);
  and _37141_ (_14908_, _14896_, _09532_);
  and _37142_ (_14909_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _37143_ (_13962_, _14909_, _14908_);
  and _37144_ (_14910_, _14896_, _09535_);
  and _37145_ (_14911_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _37146_ (_13963_, _14911_, _14910_);
  and _37147_ (_14912_, _14896_, _09538_);
  and _37148_ (_14913_, _14898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _37149_ (_13964_, _14913_, _14912_);
  and _37150_ (_14914_, _14798_, _09620_);
  and _37151_ (_14915_, _14914_, _09513_);
  not _37152_ (_14916_, _14914_);
  and _37153_ (_14917_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _37154_ (_13966_, _14917_, _14915_);
  and _37155_ (_14918_, _14914_, _09520_);
  and _37156_ (_14919_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _37157_ (_13967_, _14919_, _14918_);
  and _37158_ (_14920_, _14914_, _09523_);
  and _37159_ (_14921_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _37160_ (_13968_, _14921_, _14920_);
  and _37161_ (_14922_, _14914_, _09526_);
  and _37162_ (_14923_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _37163_ (_13970_, _14923_, _14922_);
  and _37164_ (_14924_, _14914_, _09529_);
  and _37165_ (_14925_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _37166_ (_13971_, _14925_, _14924_);
  and _37167_ (_14926_, _14914_, _09532_);
  and _37168_ (_14927_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _37169_ (_13972_, _14927_, _14926_);
  and _37170_ (_14928_, _14914_, _09535_);
  and _37171_ (_14929_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _37172_ (_13974_, _14929_, _14928_);
  and _37173_ (_14930_, _14914_, _09538_);
  and _37174_ (_14931_, _14916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _37175_ (_13975_, _14931_, _14930_);
  and _37176_ (_14932_, _14798_, _09639_);
  and _37177_ (_14933_, _14932_, _09513_);
  not _37178_ (_14934_, _14932_);
  and _37179_ (_14935_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or _37180_ (_13976_, _14935_, _14933_);
  and _37181_ (_14936_, _14932_, _09520_);
  and _37182_ (_14937_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or _37183_ (_13977_, _14937_, _14936_);
  and _37184_ (_14938_, _14932_, _09523_);
  and _37185_ (_14939_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or _37186_ (_13979_, _14939_, _14938_);
  and _37187_ (_14940_, _14932_, _09526_);
  and _37188_ (_14941_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or _37189_ (_13980_, _14941_, _14940_);
  and _37190_ (_14942_, _14932_, _09529_);
  and _37191_ (_14943_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or _37192_ (_13981_, _14943_, _14942_);
  and _37193_ (_14944_, _14932_, _09532_);
  and _37194_ (_14945_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or _37195_ (_13982_, _14945_, _14944_);
  and _37196_ (_14946_, _14932_, _09535_);
  and _37197_ (_14947_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or _37198_ (_13983_, _14947_, _14946_);
  and _37199_ (_14948_, _14932_, _09538_);
  and _37200_ (_14949_, _14934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or _37201_ (_13984_, _14949_, _14948_);
  and _37202_ (_14950_, _14798_, _09659_);
  and _37203_ (_14951_, _14950_, _09513_);
  not _37204_ (_14952_, _14950_);
  and _37205_ (_14953_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _37206_ (_13986_, _14953_, _14951_);
  and _37207_ (_14954_, _14950_, _09520_);
  and _37208_ (_14955_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _37209_ (_13987_, _14955_, _14954_);
  and _37210_ (_14956_, _14950_, _09523_);
  and _37211_ (_14957_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _37212_ (_13988_, _14957_, _14956_);
  and _37213_ (_14958_, _14950_, _09526_);
  and _37214_ (_14959_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _37215_ (_13989_, _14959_, _14958_);
  and _37216_ (_14960_, _14950_, _09529_);
  and _37217_ (_14961_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _37218_ (_13991_, _14961_, _14960_);
  and _37219_ (_14962_, _14950_, _09532_);
  and _37220_ (_14963_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _37221_ (_13992_, _14963_, _14962_);
  and _37222_ (_14964_, _14950_, _09535_);
  and _37223_ (_14965_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _37224_ (_13993_, _14965_, _14964_);
  and _37225_ (_14966_, _14950_, _09538_);
  and _37226_ (_14967_, _14952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _37227_ (_13994_, _14967_, _14966_);
  and _37228_ (_14968_, _14798_, _09678_);
  and _37229_ (_14969_, _14968_, _09513_);
  not _37230_ (_14970_, _14968_);
  and _37231_ (_14971_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or _37232_ (_13995_, _14971_, _14969_);
  and _37233_ (_14972_, _14968_, _09520_);
  and _37234_ (_14973_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or _37235_ (_13996_, _14973_, _14972_);
  and _37236_ (_14974_, _14968_, _09523_);
  and _37237_ (_14975_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or _37238_ (_13998_, _14975_, _14974_);
  and _37239_ (_14976_, _14968_, _09526_);
  and _37240_ (_14977_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or _37241_ (_13999_, _14977_, _14976_);
  and _37242_ (_14978_, _14968_, _09529_);
  and _37243_ (_14979_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or _37244_ (_14000_, _14979_, _14978_);
  and _37245_ (_14980_, _14968_, _09532_);
  and _37246_ (_14981_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or _37247_ (_14001_, _14981_, _14980_);
  and _37248_ (_14982_, _14968_, _09535_);
  and _37249_ (_14983_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or _37250_ (_14003_, _14983_, _14982_);
  and _37251_ (_14984_, _14968_, _09538_);
  and _37252_ (_14985_, _14970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or _37253_ (_14004_, _14985_, _14984_);
  and _37254_ (_14986_, _14798_, _09697_);
  and _37255_ (_14987_, _14986_, _09513_);
  not _37256_ (_14988_, _14986_);
  and _37257_ (_14989_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or _37258_ (_14005_, _14989_, _14987_);
  and _37259_ (_14990_, _14986_, _09520_);
  and _37260_ (_14991_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or _37261_ (_14006_, _14991_, _14990_);
  and _37262_ (_14992_, _14986_, _09523_);
  and _37263_ (_14993_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or _37264_ (_14007_, _14993_, _14992_);
  and _37265_ (_14994_, _14986_, _09526_);
  and _37266_ (_14995_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or _37267_ (_14008_, _14995_, _14994_);
  and _37268_ (_14996_, _14986_, _09529_);
  and _37269_ (_14997_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or _37270_ (_14010_, _14997_, _14996_);
  and _37271_ (_14998_, _14986_, _09532_);
  and _37272_ (_14999_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or _37273_ (_14011_, _14999_, _14998_);
  and _37274_ (_15000_, _14986_, _09535_);
  and _37275_ (_15001_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or _37276_ (_14012_, _15001_, _15000_);
  and _37277_ (_15002_, _14986_, _09538_);
  and _37278_ (_15003_, _14988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or _37279_ (_14013_, _15003_, _15002_);
  and _37280_ (_15004_, _14798_, _09716_);
  and _37281_ (_15005_, _15004_, _09513_);
  not _37282_ (_15006_, _15004_);
  and _37283_ (_15007_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _37284_ (_14015_, _15007_, _15005_);
  and _37285_ (_15008_, _15004_, _09520_);
  and _37286_ (_15009_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _37287_ (_14016_, _15009_, _15008_);
  and _37288_ (_15010_, _15004_, _09523_);
  and _37289_ (_15011_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _37290_ (_14017_, _15011_, _15010_);
  and _37291_ (_15012_, _15004_, _09526_);
  and _37292_ (_15013_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _37293_ (_14018_, _15013_, _15012_);
  and _37294_ (_15014_, _15004_, _09529_);
  and _37295_ (_15015_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _37296_ (_14019_, _15015_, _15014_);
  and _37297_ (_15016_, _15004_, _09532_);
  and _37298_ (_15017_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _37299_ (_14020_, _15017_, _15016_);
  and _37300_ (_15018_, _15004_, _09535_);
  and _37301_ (_15019_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _37302_ (_14022_, _15019_, _15018_);
  and _37303_ (_15020_, _15004_, _09538_);
  and _37304_ (_15021_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _37305_ (_14023_, _15021_, _15020_);
  and _37306_ (_15022_, _14798_, _09736_);
  and _37307_ (_15023_, _15022_, _09513_);
  not _37308_ (_15024_, _15022_);
  and _37309_ (_15025_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _37310_ (_14024_, _15025_, _15023_);
  and _37311_ (_15026_, _15022_, _09520_);
  and _37312_ (_15027_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _37313_ (_14025_, _15027_, _15026_);
  and _37314_ (_15028_, _15022_, _09523_);
  and _37315_ (_15029_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _37316_ (_14027_, _15029_, _15028_);
  and _37317_ (_15030_, _15022_, _09526_);
  and _37318_ (_15031_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _37319_ (_14028_, _15031_, _15030_);
  and _37320_ (_15032_, _15022_, _09529_);
  and _37321_ (_15033_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _37322_ (_14029_, _15033_, _15032_);
  and _37323_ (_15034_, _15022_, _09532_);
  and _37324_ (_15035_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _37325_ (_14030_, _15035_, _15034_);
  and _37326_ (_15036_, _15022_, _09535_);
  and _37327_ (_15037_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _37328_ (_14031_, _15037_, _15036_);
  and _37329_ (_15038_, _15022_, _09538_);
  and _37330_ (_15039_, _15024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _37331_ (_14032_, _15039_, _15038_);
  and _37332_ (_15040_, _14798_, _09755_);
  and _37333_ (_15041_, _15040_, _09513_);
  not _37334_ (_15042_, _15040_);
  and _37335_ (_15043_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or _37336_ (_14034_, _15043_, _15041_);
  and _37337_ (_15044_, _15040_, _09520_);
  and _37338_ (_15045_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or _37339_ (_14035_, _15045_, _15044_);
  and _37340_ (_15046_, _15040_, _09523_);
  and _37341_ (_15047_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or _37342_ (_14036_, _15047_, _15046_);
  and _37343_ (_15048_, _15040_, _09526_);
  and _37344_ (_15049_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or _37345_ (_14037_, _15049_, _15048_);
  and _37346_ (_15050_, _15040_, _09529_);
  and _37347_ (_15051_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or _37348_ (_14039_, _15051_, _15050_);
  and _37349_ (_15052_, _15040_, _09532_);
  and _37350_ (_15053_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or _37351_ (_14040_, _15053_, _15052_);
  and _37352_ (_15054_, _15040_, _09535_);
  and _37353_ (_15055_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or _37354_ (_14041_, _15055_, _15054_);
  and _37355_ (_15056_, _15040_, _09538_);
  and _37356_ (_15057_, _15042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or _37357_ (_14042_, _15057_, _15056_);
  and _37358_ (_15058_, _14798_, _09774_);
  and _37359_ (_15059_, _15058_, _09513_);
  not _37360_ (_15060_, _15058_);
  and _37361_ (_15061_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or _37362_ (_14043_, _15061_, _15059_);
  and _37363_ (_15062_, _15058_, _09520_);
  and _37364_ (_15063_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or _37365_ (_14044_, _15063_, _15062_);
  and _37366_ (_15064_, _15058_, _09523_);
  and _37367_ (_15065_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or _37368_ (_14046_, _15065_, _15064_);
  and _37369_ (_15066_, _15058_, _09526_);
  and _37370_ (_15067_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or _37371_ (_14047_, _15067_, _15066_);
  and _37372_ (_15068_, _15058_, _09529_);
  and _37373_ (_15069_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or _37374_ (_14048_, _15069_, _15068_);
  and _37375_ (_15070_, _15058_, _09532_);
  and _37376_ (_15071_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or _37377_ (_14049_, _15071_, _15070_);
  and _37378_ (_15072_, _15058_, _09535_);
  and _37379_ (_15073_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or _37380_ (_14051_, _15073_, _15072_);
  and _37381_ (_15074_, _15058_, _09538_);
  and _37382_ (_15075_, _15060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or _37383_ (_14052_, _15075_, _15074_);
  and _37384_ (_15076_, _14798_, _09793_);
  and _37385_ (_15077_, _15076_, _09513_);
  not _37386_ (_15078_, _15076_);
  and _37387_ (_15079_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _37388_ (_14053_, _15079_, _15077_);
  and _37389_ (_15080_, _15076_, _09520_);
  and _37390_ (_15081_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _37391_ (_14054_, _15081_, _15080_);
  and _37392_ (_15082_, _15076_, _09523_);
  and _37393_ (_15083_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _37394_ (_14055_, _15083_, _15082_);
  and _37395_ (_15084_, _15076_, _09526_);
  and _37396_ (_15085_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _37397_ (_14056_, _15085_, _15084_);
  and _37398_ (_15086_, _15076_, _09529_);
  and _37399_ (_15087_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _37400_ (_14058_, _15087_, _15086_);
  and _37401_ (_15088_, _15076_, _09532_);
  and _37402_ (_15089_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _37403_ (_14059_, _15089_, _15088_);
  and _37404_ (_15090_, _15076_, _09535_);
  and _37405_ (_15091_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _37406_ (_14060_, _15091_, _15090_);
  and _37407_ (_15092_, _15076_, _09538_);
  and _37408_ (_15093_, _15078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _37409_ (_14061_, _15093_, _15092_);
  and _37410_ (_15094_, _06008_, _02681_);
  and _37411_ (_15095_, _15094_, _09254_);
  and _37412_ (_15096_, _15095_, _09265_);
  not _37413_ (_15097_, _15096_);
  and _37414_ (_15098_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and _37415_ (_15099_, _15096_, _09334_);
  or _37416_ (_14063_, _15099_, _15098_);
  and _37417_ (_15100_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  and _37418_ (_15101_, _15096_, _09453_);
  or _37419_ (_14064_, _15101_, _15100_);
  and _37420_ (_15102_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  and _37421_ (_15103_, _15096_, _09463_);
  or _37422_ (_14065_, _15103_, _15102_);
  and _37423_ (_15104_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  and _37424_ (_15105_, _15096_, _09472_);
  or _37425_ (_14066_, _15105_, _15104_);
  and _37426_ (_15106_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  and _37427_ (_15107_, _15096_, _09482_);
  or _37428_ (_14067_, _15107_, _15106_);
  and _37429_ (_15108_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  and _37430_ (_15109_, _15096_, _09492_);
  or _37431_ (_14068_, _15109_, _15108_);
  and _37432_ (_15110_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  and _37433_ (_15111_, _15096_, _09502_);
  or _37434_ (_14070_, _15111_, _15110_);
  and _37435_ (_15112_, _15097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and _37436_ (_15113_, _15096_, _09510_);
  or _37437_ (_14071_, _15113_, _15112_);
  and _37438_ (_15114_, _15095_, _09515_);
  not _37439_ (_15115_, _15114_);
  and _37440_ (_15116_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and _37441_ (_15117_, _15114_, _09334_);
  or _37442_ (_14072_, _15117_, _15116_);
  and _37443_ (_15118_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and _37444_ (_15119_, _15114_, _09453_);
  or _37445_ (_14074_, _15119_, _15118_);
  and _37446_ (_15120_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _37447_ (_15121_, _15114_, _09463_);
  or _37448_ (_14075_, _15121_, _15120_);
  and _37449_ (_15122_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and _37450_ (_15123_, _15114_, _09472_);
  or _37451_ (_14076_, _15123_, _15122_);
  and _37452_ (_15124_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and _37453_ (_15125_, _15114_, _09482_);
  or _37454_ (_14078_, _15125_, _15124_);
  and _37455_ (_15126_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and _37456_ (_15127_, _15114_, _09492_);
  or _37457_ (_14079_, _15127_, _15126_);
  and _37458_ (_15128_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and _37459_ (_15129_, _15114_, _09502_);
  or _37460_ (_14080_, _15129_, _15128_);
  and _37461_ (_15130_, _15115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and _37462_ (_15131_, _15114_, _09510_);
  or _37463_ (_14081_, _15131_, _15130_);
  and _37464_ (_15132_, _15095_, _09542_);
  not _37465_ (_15133_, _15132_);
  and _37466_ (_15134_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and _37467_ (_15135_, _15132_, _09334_);
  or _37468_ (_14083_, _15135_, _15134_);
  and _37469_ (_15136_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _37470_ (_15137_, _15132_, _09453_);
  or _37471_ (_14084_, _15137_, _15136_);
  and _37472_ (_15138_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and _37473_ (_15139_, _15132_, _09463_);
  or _37474_ (_14085_, _15139_, _15138_);
  and _37475_ (_15140_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and _37476_ (_15141_, _15132_, _09472_);
  or _37477_ (_14086_, _15141_, _15140_);
  and _37478_ (_15142_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and _37479_ (_15143_, _15132_, _09482_);
  or _37480_ (_14087_, _15143_, _15142_);
  and _37481_ (_15144_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and _37482_ (_15145_, _15132_, _09492_);
  or _37483_ (_14088_, _15145_, _15144_);
  and _37484_ (_15146_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and _37485_ (_15147_, _15132_, _09502_);
  or _37486_ (_14090_, _15147_, _15146_);
  and _37487_ (_15148_, _15133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and _37488_ (_15149_, _15132_, _09510_);
  or _37489_ (_14091_, _15149_, _15148_);
  and _37490_ (_15150_, _15095_, _09562_);
  not _37491_ (_15151_, _15150_);
  and _37492_ (_15152_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and _37493_ (_15153_, _15150_, _09334_);
  or _37494_ (_14092_, _15153_, _15152_);
  and _37495_ (_15154_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  and _37496_ (_15155_, _15150_, _09453_);
  or _37497_ (_14093_, _15155_, _15154_);
  and _37498_ (_15156_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  and _37499_ (_15157_, _15150_, _09463_);
  or _37500_ (_14095_, _15157_, _15156_);
  and _37501_ (_15158_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  and _37502_ (_15159_, _15150_, _09472_);
  or _37503_ (_14096_, _15159_, _15158_);
  and _37504_ (_15160_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  and _37505_ (_15161_, _15150_, _09482_);
  or _37506_ (_14097_, _15161_, _15160_);
  and _37507_ (_15162_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  and _37508_ (_15163_, _15150_, _09492_);
  or _37509_ (_14098_, _15163_, _15162_);
  and _37510_ (_15164_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  and _37511_ (_15165_, _15150_, _09502_);
  or _37512_ (_14099_, _15165_, _15164_);
  and _37513_ (_15166_, _15151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  and _37514_ (_15167_, _15150_, _09510_);
  or _37515_ (_14100_, _15167_, _15166_);
  and _37516_ (_15168_, _15095_, _09582_);
  not _37517_ (_15169_, _15168_);
  and _37518_ (_15170_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and _37519_ (_15171_, _15168_, _09334_);
  or _37520_ (_14102_, _15171_, _15170_);
  and _37521_ (_15172_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  and _37522_ (_15173_, _15168_, _09453_);
  or _37523_ (_14103_, _15173_, _15172_);
  and _37524_ (_15174_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  and _37525_ (_15175_, _15168_, _09463_);
  or _37526_ (_14104_, _15175_, _15174_);
  and _37527_ (_15176_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  and _37528_ (_15177_, _15168_, _09472_);
  or _37529_ (_14105_, _15177_, _15176_);
  and _37530_ (_15178_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  and _37531_ (_15179_, _15168_, _09482_);
  or _37532_ (_14107_, _15179_, _15178_);
  and _37533_ (_15180_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  and _37534_ (_15181_, _15168_, _09492_);
  or _37535_ (_14108_, _15181_, _15180_);
  and _37536_ (_15182_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  and _37537_ (_15183_, _15168_, _09502_);
  or _37538_ (_14109_, _15183_, _15182_);
  and _37539_ (_15184_, _15169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  and _37540_ (_15185_, _15168_, _09510_);
  or _37541_ (_14110_, _15185_, _15184_);
  and _37542_ (_15186_, _15095_, _09601_);
  not _37543_ (_15187_, _15186_);
  and _37544_ (_15188_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and _37545_ (_15189_, _15186_, _09334_);
  or _37546_ (_14111_, _15189_, _15188_);
  and _37547_ (_15190_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and _37548_ (_15191_, _15186_, _09453_);
  or _37549_ (_14112_, _15191_, _15190_);
  and _37550_ (_15192_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and _37551_ (_15193_, _15186_, _09463_);
  or _37552_ (_14114_, _15193_, _15192_);
  and _37553_ (_15194_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and _37554_ (_15195_, _15186_, _09472_);
  or _37555_ (_14115_, _15195_, _15194_);
  and _37556_ (_15196_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _37557_ (_15197_, _15186_, _09482_);
  or _37558_ (_14116_, _15197_, _15196_);
  and _37559_ (_15198_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and _37560_ (_15199_, _15186_, _09492_);
  or _37561_ (_14117_, _15199_, _15198_);
  and _37562_ (_15200_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and _37563_ (_15201_, _15186_, _09502_);
  or _37564_ (_14119_, _15201_, _15200_);
  and _37565_ (_15202_, _15187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and _37566_ (_15203_, _15186_, _09510_);
  or _37567_ (_14120_, _15203_, _15202_);
  and _37568_ (_15204_, _15095_, _09620_);
  not _37569_ (_15205_, _15204_);
  and _37570_ (_15206_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and _37571_ (_15207_, _15204_, _09334_);
  or _37572_ (_14121_, _15207_, _15206_);
  and _37573_ (_15208_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and _37574_ (_15209_, _15204_, _09453_);
  or _37575_ (_14122_, _15209_, _15208_);
  and _37576_ (_15210_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _37577_ (_15211_, _15204_, _09463_);
  or _37578_ (_14123_, _15211_, _15210_);
  and _37579_ (_15212_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and _37580_ (_15213_, _15204_, _09472_);
  or _37581_ (_14124_, _15213_, _15212_);
  and _37582_ (_15214_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and _37583_ (_15215_, _15204_, _09482_);
  or _37584_ (_14126_, _15215_, _15214_);
  and _37585_ (_15216_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and _37586_ (_15217_, _15204_, _09492_);
  or _37587_ (_14127_, _15217_, _15216_);
  and _37588_ (_15218_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and _37589_ (_15219_, _15204_, _09502_);
  or _37590_ (_14128_, _15219_, _15218_);
  and _37591_ (_15220_, _15205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and _37592_ (_15221_, _15204_, _09510_);
  or _37593_ (_14129_, _15221_, _15220_);
  and _37594_ (_15222_, _15095_, _09639_);
  not _37595_ (_15223_, _15222_);
  and _37596_ (_15224_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and _37597_ (_15225_, _15222_, _09334_);
  or _37598_ (_14131_, _15225_, _15224_);
  and _37599_ (_15226_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  and _37600_ (_15227_, _15222_, _09453_);
  or _37601_ (_14132_, _15227_, _15226_);
  and _37602_ (_15228_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  and _37603_ (_15229_, _15222_, _09463_);
  or _37604_ (_14133_, _15229_, _15228_);
  and _37605_ (_15230_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  and _37606_ (_15231_, _15222_, _09472_);
  or _37607_ (_14134_, _15231_, _15230_);
  and _37608_ (_15232_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  and _37609_ (_15233_, _15222_, _09482_);
  or _37610_ (_14135_, _15233_, _15232_);
  and _37611_ (_15234_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  and _37612_ (_15235_, _15222_, _09492_);
  or _37613_ (_14136_, _15235_, _15234_);
  and _37614_ (_15236_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  and _37615_ (_15237_, _15222_, _09502_);
  or _37616_ (_14138_, _15237_, _15236_);
  and _37617_ (_15238_, _15223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and _37618_ (_15239_, _15222_, _09510_);
  or _37619_ (_14139_, _15239_, _15238_);
  and _37620_ (_15240_, _15095_, _09659_);
  not _37621_ (_15241_, _15240_);
  and _37622_ (_15242_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and _37623_ (_15243_, _15240_, _09334_);
  or _37624_ (_14140_, _15243_, _15242_);
  and _37625_ (_15244_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and _37626_ (_15245_, _15240_, _09453_);
  or _37627_ (_14141_, _15245_, _15244_);
  and _37628_ (_15246_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and _37629_ (_15247_, _15240_, _09463_);
  or _37630_ (_14143_, _15247_, _15246_);
  and _37631_ (_15248_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and _37632_ (_15249_, _15240_, _09472_);
  or _37633_ (_14144_, _15249_, _15248_);
  and _37634_ (_15250_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and _37635_ (_15251_, _15240_, _09482_);
  or _37636_ (_14145_, _15251_, _15250_);
  and _37637_ (_15252_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and _37638_ (_15253_, _15240_, _09492_);
  or _37639_ (_14146_, _15253_, _15252_);
  and _37640_ (_15254_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _37641_ (_15255_, _15240_, _09502_);
  or _37642_ (_14147_, _15255_, _15254_);
  and _37643_ (_15256_, _15241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and _37644_ (_15257_, _15240_, _09510_);
  or _37645_ (_14148_, _15257_, _15256_);
  and _37646_ (_15258_, _15095_, _09678_);
  not _37647_ (_15259_, _15258_);
  and _37648_ (_15260_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and _37649_ (_15261_, _15258_, _09334_);
  or _37650_ (_14150_, _15261_, _15260_);
  and _37651_ (_15262_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  and _37652_ (_15263_, _15258_, _09453_);
  or _37653_ (_14151_, _15263_, _15262_);
  and _37654_ (_15264_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  and _37655_ (_15265_, _15258_, _09463_);
  or _37656_ (_14152_, _15265_, _15264_);
  and _37657_ (_15266_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  and _37658_ (_15267_, _15258_, _09472_);
  or _37659_ (_14153_, _15267_, _15266_);
  and _37660_ (_15268_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  and _37661_ (_15269_, _15258_, _09482_);
  or _37662_ (_14155_, _15269_, _15268_);
  and _37663_ (_15270_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and _37664_ (_15271_, _15258_, _09492_);
  or _37665_ (_14156_, _15271_, _15270_);
  and _37666_ (_15272_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  and _37667_ (_15273_, _15258_, _09502_);
  or _37668_ (_14157_, _15273_, _15272_);
  and _37669_ (_15274_, _15259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  and _37670_ (_15275_, _15258_, _09510_);
  or _37671_ (_14158_, _15275_, _15274_);
  and _37672_ (_15276_, _15095_, _09697_);
  not _37673_ (_15277_, _15276_);
  and _37674_ (_15278_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and _37675_ (_15279_, _15276_, _09334_);
  or _37676_ (_14159_, _15279_, _15278_);
  and _37677_ (_15280_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  and _37678_ (_15281_, _15276_, _09453_);
  or _37679_ (_14160_, _15281_, _15280_);
  and _37680_ (_15282_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  and _37681_ (_15283_, _15276_, _09463_);
  or _37682_ (_14162_, _15283_, _15282_);
  and _37683_ (_15284_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  and _37684_ (_15285_, _15276_, _09472_);
  or _37685_ (_14163_, _15285_, _15284_);
  and _37686_ (_15286_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  and _37687_ (_15287_, _15276_, _09482_);
  or _37688_ (_14164_, _15287_, _15286_);
  and _37689_ (_15288_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  and _37690_ (_15289_, _15276_, _09492_);
  or _37691_ (_14165_, _15289_, _15288_);
  and _37692_ (_15290_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  and _37693_ (_15291_, _15276_, _09502_);
  or _37694_ (_14167_, _15291_, _15290_);
  and _37695_ (_15292_, _15277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and _37696_ (_15293_, _15276_, _09510_);
  or _37697_ (_14168_, _15293_, _15292_);
  and _37698_ (_15294_, _15095_, _09716_);
  not _37699_ (_15295_, _15294_);
  and _37700_ (_15296_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and _37701_ (_15297_, _15294_, _09334_);
  or _37702_ (_14169_, _15297_, _15296_);
  and _37703_ (_15298_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and _37704_ (_15299_, _15294_, _09453_);
  or _37705_ (_14170_, _15299_, _15298_);
  and _37706_ (_15300_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and _37707_ (_15301_, _15294_, _09463_);
  or _37708_ (_14171_, _15301_, _15300_);
  and _37709_ (_15302_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and _37710_ (_15303_, _15294_, _09472_);
  or _37711_ (_14172_, _15303_, _15302_);
  and _37712_ (_15304_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _37713_ (_15305_, _15294_, _09482_);
  or _37714_ (_14174_, _15305_, _15304_);
  and _37715_ (_15306_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and _37716_ (_15307_, _15294_, _09492_);
  or _37717_ (_14175_, _15307_, _15306_);
  and _37718_ (_15308_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and _37719_ (_15309_, _15294_, _09502_);
  or _37720_ (_14176_, _15309_, _15308_);
  and _37721_ (_15310_, _15295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and _37722_ (_15311_, _15294_, _09510_);
  or _37723_ (_14177_, _15311_, _15310_);
  and _37724_ (_15312_, _15095_, _09736_);
  not _37725_ (_15313_, _15312_);
  and _37726_ (_15314_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and _37727_ (_15315_, _15312_, _09334_);
  or _37728_ (_14179_, _15315_, _15314_);
  and _37729_ (_15316_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and _37730_ (_15317_, _15312_, _09453_);
  or _37731_ (_14180_, _15317_, _15316_);
  and _37732_ (_15318_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _37733_ (_15319_, _15312_, _09463_);
  or _37734_ (_14181_, _15319_, _15318_);
  and _37735_ (_15320_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and _37736_ (_15321_, _15312_, _09472_);
  or _37737_ (_14183_, _15321_, _15320_);
  and _37738_ (_15322_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and _37739_ (_15323_, _15312_, _09482_);
  or _37740_ (_14184_, _15323_, _15322_);
  and _37741_ (_15324_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and _37742_ (_15325_, _15312_, _09492_);
  or _37743_ (_14185_, _15325_, _15324_);
  and _37744_ (_15326_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and _37745_ (_15327_, _15312_, _09502_);
  or _37746_ (_14187_, _15327_, _15326_);
  and _37747_ (_15328_, _15313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and _37748_ (_15329_, _15312_, _09510_);
  or _37749_ (_14188_, _15329_, _15328_);
  and _37750_ (_15330_, _15095_, _09755_);
  not _37751_ (_15331_, _15330_);
  and _37752_ (_15332_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and _37753_ (_15333_, _15330_, _09334_);
  or _37754_ (_14189_, _15333_, _15332_);
  and _37755_ (_15334_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  and _37756_ (_15335_, _15330_, _09453_);
  or _37757_ (_14190_, _15335_, _15334_);
  and _37758_ (_15336_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  and _37759_ (_15337_, _15330_, _09463_);
  or _37760_ (_14191_, _15337_, _15336_);
  and _37761_ (_15338_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  and _37762_ (_15339_, _15330_, _09472_);
  or _37763_ (_14192_, _15339_, _15338_);
  and _37764_ (_15340_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  and _37765_ (_15341_, _15330_, _09482_);
  or _37766_ (_14193_, _15341_, _15340_);
  and _37767_ (_15342_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  and _37768_ (_15343_, _15330_, _09492_);
  or _37769_ (_14195_, _15343_, _15342_);
  and _37770_ (_15344_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  and _37771_ (_15345_, _15330_, _09502_);
  or _37772_ (_14196_, _15345_, _15344_);
  and _37773_ (_15346_, _15331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  and _37774_ (_15347_, _15330_, _09510_);
  or _37775_ (_14197_, _15347_, _15346_);
  and _37776_ (_15348_, _15095_, _09774_);
  not _37777_ (_15349_, _15348_);
  and _37778_ (_15350_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and _37779_ (_15351_, _15348_, _09334_);
  or _37780_ (_14199_, _15351_, _15350_);
  and _37781_ (_15352_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  and _37782_ (_15353_, _15348_, _09453_);
  or _37783_ (_14200_, _15353_, _15352_);
  and _37784_ (_15354_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  and _37785_ (_15355_, _15348_, _09463_);
  or _37786_ (_14201_, _15355_, _15354_);
  and _37787_ (_15356_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  and _37788_ (_15357_, _15348_, _09472_);
  or _37789_ (_14202_, _15357_, _15356_);
  and _37790_ (_15358_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  and _37791_ (_15359_, _15348_, _09482_);
  or _37792_ (_14203_, _15359_, _15358_);
  and _37793_ (_15360_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  and _37794_ (_15361_, _15348_, _09492_);
  or _37795_ (_14204_, _15361_, _15360_);
  and _37796_ (_15362_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  and _37797_ (_15363_, _15348_, _09502_);
  or _37798_ (_14205_, _15363_, _15362_);
  and _37799_ (_15364_, _15349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and _37800_ (_15365_, _15348_, _09510_);
  or _37801_ (_14207_, _15365_, _15364_);
  and _37802_ (_15366_, _15095_, _09793_);
  not _37803_ (_15367_, _15366_);
  and _37804_ (_15368_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and _37805_ (_15369_, _15366_, _09334_);
  or _37806_ (_14208_, _15369_, _15368_);
  and _37807_ (_15370_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and _37808_ (_15371_, _15366_, _09453_);
  or _37809_ (_14209_, _15371_, _15370_);
  and _37810_ (_15372_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and _37811_ (_15373_, _15366_, _09463_);
  or _37812_ (_14211_, _15373_, _15372_);
  and _37813_ (_15374_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and _37814_ (_15375_, _15366_, _09472_);
  or _37815_ (_14212_, _15375_, _15374_);
  and _37816_ (_15376_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and _37817_ (_15377_, _15366_, _09482_);
  or _37818_ (_14213_, _15377_, _15376_);
  and _37819_ (_15378_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and _37820_ (_15379_, _15366_, _09492_);
  or _37821_ (_14214_, _15379_, _15378_);
  and _37822_ (_15380_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _37823_ (_15381_, _15366_, _09502_);
  or _37824_ (_14215_, _15381_, _15380_);
  and _37825_ (_15382_, _15367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and _37826_ (_15383_, _15366_, _09510_);
  or _37827_ (_14216_, _15383_, _15382_);
  and _37828_ (_15384_, _09813_, _02681_);
  and _37829_ (_15385_, _15384_, _09265_);
  and _37830_ (_15386_, _15385_, _09513_);
  not _37831_ (_15387_, _15385_);
  and _37832_ (_15388_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  or _37833_ (_14217_, _15388_, _15386_);
  and _37834_ (_15389_, _15385_, _09520_);
  and _37835_ (_15390_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  or _37836_ (_14219_, _15390_, _15389_);
  and _37837_ (_15391_, _15385_, _09523_);
  and _37838_ (_15392_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  or _37839_ (_14220_, _15392_, _15391_);
  and _37840_ (_15393_, _15385_, _09526_);
  and _37841_ (_15394_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  or _37842_ (_14221_, _15394_, _15393_);
  and _37843_ (_15395_, _15385_, _09529_);
  and _37844_ (_15396_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  or _37845_ (_14223_, _15396_, _15395_);
  and _37846_ (_15397_, _15385_, _09532_);
  and _37847_ (_15398_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  or _37848_ (_14224_, _15398_, _15397_);
  and _37849_ (_15399_, _15385_, _09535_);
  and _37850_ (_15400_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  or _37851_ (_14225_, _15400_, _15399_);
  and _37852_ (_15401_, _15385_, _09538_);
  and _37853_ (_15402_, _15387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  or _37854_ (_14226_, _15402_, _15401_);
  and _37855_ (_15403_, _15384_, _09515_);
  and _37856_ (_15404_, _15403_, _09513_);
  not _37857_ (_15405_, _15403_);
  and _37858_ (_15406_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _37859_ (_14227_, _15406_, _15404_);
  and _37860_ (_15407_, _15403_, _09520_);
  and _37861_ (_15408_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _37862_ (_14228_, _15408_, _15407_);
  and _37863_ (_15409_, _15403_, _09523_);
  and _37864_ (_15410_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _37865_ (_14229_, _15410_, _15409_);
  and _37866_ (_15411_, _15403_, _09526_);
  and _37867_ (_15412_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or _37868_ (_14231_, _15412_, _15411_);
  and _37869_ (_15413_, _15403_, _09529_);
  and _37870_ (_15414_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or _37871_ (_14232_, _15414_, _15413_);
  and _37872_ (_15415_, _15403_, _09532_);
  and _37873_ (_15416_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _37874_ (_14233_, _15416_, _15415_);
  and _37875_ (_15417_, _15403_, _09535_);
  and _37876_ (_15418_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or _37877_ (_14235_, _15418_, _15417_);
  and _37878_ (_15419_, _15403_, _09538_);
  and _37879_ (_15420_, _15405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _37880_ (_14236_, _15420_, _15419_);
  and _37881_ (_15421_, _15384_, _09542_);
  and _37882_ (_15422_, _15421_, _09513_);
  not _37883_ (_15423_, _15421_);
  and _37884_ (_15424_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or _37885_ (_14237_, _15424_, _15422_);
  and _37886_ (_15425_, _15421_, _09520_);
  and _37887_ (_15426_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or _37888_ (_14238_, _15426_, _15425_);
  and _37889_ (_15427_, _15421_, _09523_);
  and _37890_ (_15428_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or _37891_ (_14239_, _15428_, _15427_);
  and _37892_ (_15429_, _15421_, _09526_);
  and _37893_ (_15430_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _37894_ (_14240_, _15430_, _15429_);
  and _37895_ (_15431_, _15421_, _09529_);
  and _37896_ (_15432_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _37897_ (_14241_, _15432_, _15431_);
  and _37898_ (_15433_, _15421_, _09532_);
  and _37899_ (_15434_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or _37900_ (_14243_, _15434_, _15433_);
  and _37901_ (_15435_, _15421_, _09535_);
  and _37902_ (_15436_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _37903_ (_14244_, _15436_, _15435_);
  and _37904_ (_15437_, _15421_, _09538_);
  and _37905_ (_15438_, _15423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _37906_ (_14245_, _15438_, _15437_);
  and _37907_ (_15439_, _15384_, _09562_);
  and _37908_ (_15440_, _15439_, _09513_);
  not _37909_ (_15441_, _15439_);
  and _37910_ (_15442_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  or _37911_ (_14247_, _15442_, _15440_);
  and _37912_ (_15443_, _15439_, _09520_);
  and _37913_ (_15444_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  or _37914_ (_14248_, _15444_, _15443_);
  and _37915_ (_15445_, _15439_, _09523_);
  and _37916_ (_15446_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  or _37917_ (_14249_, _15446_, _15445_);
  and _37918_ (_15447_, _15439_, _09526_);
  and _37919_ (_15448_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  or _37920_ (_14250_, _15448_, _15447_);
  and _37921_ (_15449_, _15439_, _09529_);
  and _37922_ (_15450_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  or _37923_ (_14251_, _15450_, _15449_);
  and _37924_ (_15451_, _15439_, _09532_);
  and _37925_ (_15452_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  or _37926_ (_14252_, _15452_, _15451_);
  and _37927_ (_15453_, _15439_, _09535_);
  and _37928_ (_15454_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  or _37929_ (_14253_, _15454_, _15453_);
  and _37930_ (_15455_, _15439_, _09538_);
  and _37931_ (_15456_, _15441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  or _37932_ (_14255_, _15456_, _15455_);
  and _37933_ (_15458_, _15384_, _09582_);
  and _37934_ (_15459_, _15458_, _09513_);
  not _37935_ (_15460_, _15458_);
  and _37936_ (_15461_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  or _37937_ (_14256_, _15461_, _15459_);
  and _37938_ (_15462_, _15458_, _09520_);
  and _37939_ (_15463_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  or _37940_ (_14257_, _15463_, _15462_);
  and _37941_ (_15464_, _15458_, _09523_);
  and _37942_ (_15465_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  or _37943_ (_14259_, _15465_, _15464_);
  and _37944_ (_15466_, _15458_, _09526_);
  and _37945_ (_15467_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  or _37946_ (_14260_, _15467_, _15466_);
  and _37947_ (_15468_, _15458_, _09529_);
  and _37948_ (_15469_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  or _37949_ (_14261_, _15469_, _15468_);
  and _37950_ (_15470_, _15458_, _09532_);
  and _37951_ (_15471_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or _37952_ (_14262_, _15471_, _15470_);
  and _37953_ (_15473_, _15458_, _09535_);
  and _37954_ (_15474_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  or _37955_ (_14263_, _15474_, _15473_);
  and _37956_ (_15475_, _15458_, _09538_);
  and _37957_ (_15476_, _15460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or _37958_ (_14264_, _15476_, _15475_);
  and _37959_ (_15477_, _15384_, _09601_);
  and _37960_ (_15478_, _15477_, _09513_);
  not _37961_ (_15479_, _15477_);
  and _37962_ (_15480_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or _37963_ (_14265_, _15480_, _15478_);
  and _37964_ (_15481_, _15477_, _09520_);
  and _37965_ (_15482_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or _37966_ (_14267_, _15482_, _15481_);
  and _37967_ (_15483_, _15477_, _09523_);
  and _37968_ (_15484_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _37969_ (_14268_, _15484_, _15483_);
  and _37970_ (_15485_, _15477_, _09526_);
  and _37971_ (_15486_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _37972_ (_14269_, _15486_, _15485_);
  and _37973_ (_15487_, _15477_, _09529_);
  and _37974_ (_15488_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or _37975_ (_14271_, _15488_, _15487_);
  and _37976_ (_15489_, _15477_, _09532_);
  and _37977_ (_15490_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _37978_ (_14272_, _15490_, _15489_);
  and _37979_ (_15491_, _15477_, _09535_);
  and _37980_ (_15492_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _37981_ (_14273_, _15492_, _15491_);
  and _37982_ (_15493_, _15477_, _09538_);
  and _37983_ (_15494_, _15479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _37984_ (_14274_, _15494_, _15493_);
  and _37985_ (_15495_, _15384_, _09620_);
  and _37986_ (_15496_, _15495_, _09513_);
  not _37987_ (_15497_, _15495_);
  and _37988_ (_15498_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _37989_ (_14275_, _15498_, _15496_);
  and _37990_ (_15499_, _15495_, _09520_);
  and _37991_ (_15500_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _37992_ (_14276_, _15500_, _15499_);
  and _37993_ (_15501_, _15495_, _09523_);
  and _37994_ (_15502_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or _37995_ (_14277_, _15502_, _15501_);
  and _37996_ (_15503_, _15495_, _09526_);
  and _37997_ (_15504_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or _37998_ (_14279_, _15504_, _15503_);
  and _37999_ (_15505_, _15495_, _09529_);
  and _38000_ (_15506_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _38001_ (_14280_, _15506_, _15505_);
  and _38002_ (_15507_, _15495_, _09532_);
  and _38003_ (_15508_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _38004_ (_14281_, _15508_, _15507_);
  and _38005_ (_15509_, _15495_, _09535_);
  and _38006_ (_15510_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or _38007_ (_14283_, _15510_, _15509_);
  and _38008_ (_15511_, _15495_, _09538_);
  and _38009_ (_15512_, _15497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _38010_ (_14284_, _15512_, _15511_);
  and _38011_ (_15513_, _15384_, _09639_);
  and _38012_ (_15514_, _15513_, _09513_);
  not _38013_ (_15515_, _15513_);
  and _38014_ (_15516_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  or _38015_ (_14285_, _15516_, _15514_);
  and _38016_ (_15517_, _15513_, _09520_);
  and _38017_ (_15518_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  or _38018_ (_14287_, _15518_, _15517_);
  and _38019_ (_15519_, _15513_, _09523_);
  and _38020_ (_15520_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  or _38021_ (_14288_, _15520_, _15519_);
  and _38022_ (_15521_, _15513_, _09526_);
  and _38023_ (_15522_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  or _38024_ (_14289_, _15522_, _15521_);
  and _38025_ (_15523_, _15513_, _09529_);
  and _38026_ (_15524_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  or _38027_ (_14290_, _15524_, _15523_);
  and _38028_ (_15525_, _15513_, _09532_);
  and _38029_ (_15526_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  or _38030_ (_14292_, _15526_, _15525_);
  and _38031_ (_15527_, _15513_, _09535_);
  and _38032_ (_15528_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  or _38033_ (_14293_, _15528_, _15527_);
  and _38034_ (_15529_, _15513_, _09538_);
  and _38035_ (_15530_, _15515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  or _38036_ (_14294_, _15530_, _15529_);
  and _38037_ (_15531_, _15384_, _09659_);
  and _38038_ (_15532_, _15531_, _09513_);
  not _38039_ (_15533_, _15531_);
  and _38040_ (_15534_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _38041_ (_14295_, _15534_, _15532_);
  and _38042_ (_15535_, _15531_, _09520_);
  and _38043_ (_15536_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _38044_ (_14296_, _15536_, _15535_);
  and _38045_ (_15537_, _15531_, _09523_);
  and _38046_ (_15538_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or _38047_ (_14297_, _15538_, _15537_);
  and _38048_ (_15539_, _15531_, _09526_);
  and _38049_ (_15540_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or _38050_ (_14299_, _15540_, _15539_);
  and _38051_ (_15541_, _15531_, _09529_);
  and _38052_ (_15542_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or _38053_ (_14300_, _15542_, _15541_);
  and _38054_ (_15543_, _15531_, _09532_);
  and _38055_ (_15544_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _38056_ (_14301_, _15544_, _15543_);
  and _38057_ (_15545_, _15531_, _09535_);
  and _38058_ (_15546_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or _38059_ (_14302_, _15546_, _15545_);
  and _38060_ (_15547_, _15531_, _09538_);
  and _38061_ (_15548_, _15533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _38062_ (_14304_, _15548_, _15547_);
  and _38063_ (_15549_, _15384_, _09678_);
  and _38064_ (_15550_, _15549_, _09513_);
  not _38065_ (_15551_, _15549_);
  and _38066_ (_15552_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  or _38067_ (_14305_, _15552_, _15550_);
  and _38068_ (_15553_, _15549_, _09520_);
  and _38069_ (_15554_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  or _38070_ (_14306_, _15554_, _15553_);
  and _38071_ (_15555_, _15549_, _09523_);
  and _38072_ (_15556_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  or _38073_ (_14307_, _15556_, _15555_);
  and _38074_ (_15557_, _15549_, _09526_);
  and _38075_ (_15558_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  or _38076_ (_14308_, _15558_, _15557_);
  and _38077_ (_15559_, _15549_, _09529_);
  and _38078_ (_15560_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  or _38079_ (_14309_, _15560_, _15559_);
  and _38080_ (_15561_, _15549_, _09532_);
  and _38081_ (_15562_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or _38082_ (_14311_, _15562_, _15561_);
  and _38083_ (_15563_, _15549_, _09535_);
  and _38084_ (_15564_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  or _38085_ (_14312_, _15564_, _15563_);
  and _38086_ (_15565_, _15549_, _09538_);
  and _38087_ (_15566_, _15551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  or _38088_ (_14313_, _15566_, _15565_);
  and _38089_ (_15567_, _15384_, _09697_);
  and _38090_ (_15568_, _15567_, _09513_);
  not _38091_ (_15569_, _15567_);
  and _38092_ (_15570_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  or _38093_ (_14314_, _15570_, _15568_);
  and _38094_ (_15571_, _15567_, _09520_);
  and _38095_ (_15572_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  or _38096_ (_14316_, _15572_, _15571_);
  and _38097_ (_15573_, _15567_, _09523_);
  and _38098_ (_15574_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  or _38099_ (_14317_, _15574_, _15573_);
  and _38100_ (_15575_, _15567_, _09526_);
  and _38101_ (_15576_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  or _38102_ (_14318_, _15576_, _15575_);
  and _38103_ (_15577_, _15567_, _09529_);
  and _38104_ (_15578_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  or _38105_ (_14319_, _15578_, _15577_);
  and _38106_ (_15579_, _15567_, _09532_);
  and _38107_ (_15580_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  or _38108_ (_14320_, _15580_, _15579_);
  and _38109_ (_15581_, _15567_, _09535_);
  and _38110_ (_15582_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  or _38111_ (_14321_, _15582_, _15581_);
  and _38112_ (_15583_, _15567_, _09538_);
  and _38113_ (_15584_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  or _38114_ (_14322_, _15584_, _15583_);
  and _38115_ (_15585_, _15384_, _09716_);
  and _38116_ (_15586_, _15585_, _09513_);
  not _38117_ (_15587_, _15585_);
  and _38118_ (_15588_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or _38119_ (_14324_, _15588_, _15586_);
  and _38120_ (_15589_, _15585_, _09520_);
  and _38121_ (_15590_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or _38122_ (_14325_, _15590_, _15589_);
  and _38123_ (_15591_, _15585_, _09523_);
  and _38124_ (_15592_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _38125_ (_14326_, _15592_, _15591_);
  and _38126_ (_15593_, _15585_, _09526_);
  and _38127_ (_15594_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _38128_ (_14328_, _15594_, _15593_);
  and _38129_ (_15595_, _15585_, _09529_);
  and _38130_ (_15596_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or _38131_ (_14329_, _15596_, _15595_);
  and _38132_ (_15597_, _15585_, _09532_);
  and _38133_ (_15598_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _38134_ (_14330_, _15598_, _15597_);
  and _38135_ (_15599_, _15585_, _09535_);
  and _38136_ (_15600_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or _38137_ (_14331_, _15600_, _15599_);
  and _38138_ (_15601_, _15585_, _09538_);
  and _38139_ (_15602_, _15587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or _38140_ (_14332_, _15602_, _15601_);
  and _38141_ (_15603_, _15384_, _09736_);
  and _38142_ (_15604_, _15603_, _09513_);
  not _38143_ (_15605_, _15603_);
  and _38144_ (_15606_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _38145_ (_14333_, _15606_, _15604_);
  and _38146_ (_15607_, _15603_, _09520_);
  and _38147_ (_15608_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _38148_ (_14335_, _15608_, _15607_);
  and _38149_ (_15609_, _15603_, _09523_);
  and _38150_ (_15610_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or _38151_ (_14336_, _15610_, _15609_);
  and _38152_ (_15611_, _15603_, _09526_);
  and _38153_ (_15612_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or _38154_ (_14337_, _15612_, _15611_);
  and _38155_ (_15613_, _15603_, _09529_);
  and _38156_ (_15614_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _38157_ (_14338_, _15614_, _15613_);
  and _38158_ (_15615_, _15603_, _09532_);
  and _38159_ (_15616_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or _38160_ (_14340_, _15616_, _15615_);
  and _38161_ (_15617_, _15603_, _09535_);
  and _38162_ (_15618_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _38163_ (_14341_, _15618_, _15617_);
  and _38164_ (_15619_, _15603_, _09538_);
  and _38165_ (_15620_, _15605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _38166_ (_14342_, _15620_, _15619_);
  and _38167_ (_15621_, _15384_, _09755_);
  and _38168_ (_15622_, _15621_, _09513_);
  not _38169_ (_15623_, _15621_);
  and _38170_ (_15624_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  or _38171_ (_14343_, _15624_, _15622_);
  and _38172_ (_15625_, _15621_, _09520_);
  and _38173_ (_15626_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  or _38174_ (_14344_, _15626_, _15625_);
  and _38175_ (_15627_, _15621_, _09523_);
  and _38176_ (_15628_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  or _38177_ (_14345_, _15628_, _15627_);
  and _38178_ (_15629_, _15621_, _09526_);
  and _38179_ (_15630_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  or _38180_ (_14347_, _15630_, _15629_);
  and _38181_ (_15631_, _15621_, _09529_);
  and _38182_ (_15632_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  or _38183_ (_14348_, _15632_, _15631_);
  and _38184_ (_15633_, _15621_, _09532_);
  and _38185_ (_15634_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or _38186_ (_14349_, _15634_, _15633_);
  and _38187_ (_15635_, _15621_, _09535_);
  and _38188_ (_15636_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  or _38189_ (_14350_, _15636_, _15635_);
  and _38190_ (_15637_, _15621_, _09538_);
  and _38191_ (_15638_, _15623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  or _38192_ (_14352_, _15638_, _15637_);
  and _38193_ (_15639_, _15384_, _09774_);
  and _38194_ (_15640_, _15639_, _09513_);
  not _38195_ (_15641_, _15639_);
  and _38196_ (_15642_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  or _38197_ (_14353_, _15642_, _15640_);
  and _38198_ (_15643_, _15639_, _09520_);
  and _38199_ (_15644_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  or _38200_ (_14354_, _15644_, _15643_);
  and _38201_ (_15645_, _15639_, _09523_);
  and _38202_ (_15646_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  or _38203_ (_14355_, _15646_, _15645_);
  and _38204_ (_15647_, _15639_, _09526_);
  and _38205_ (_15648_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  or _38206_ (_14356_, _15648_, _15647_);
  and _38207_ (_15649_, _15639_, _09529_);
  and _38208_ (_15650_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  or _38209_ (_14357_, _15650_, _15649_);
  and _38210_ (_15651_, _15639_, _09532_);
  and _38211_ (_15652_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  or _38212_ (_14359_, _15652_, _15651_);
  and _38213_ (_15653_, _15639_, _09535_);
  and _38214_ (_15654_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  or _38215_ (_14360_, _15654_, _15653_);
  and _38216_ (_15655_, _15639_, _09538_);
  and _38217_ (_15656_, _15641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  or _38218_ (_14361_, _15656_, _15655_);
  and _38219_ (_15657_, _15384_, _09793_);
  and _38220_ (_15658_, _15657_, _09513_);
  not _38221_ (_15659_, _15657_);
  and _38222_ (_15660_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or _38223_ (_14362_, _15660_, _15658_);
  and _38224_ (_15661_, _15657_, _09520_);
  and _38225_ (_15662_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _38226_ (_14364_, _15662_, _15661_);
  and _38227_ (_15663_, _15657_, _09523_);
  and _38228_ (_15664_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or _38229_ (_14365_, _15664_, _15663_);
  and _38230_ (_15665_, _15657_, _09526_);
  and _38231_ (_15666_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _38232_ (_14366_, _15666_, _15665_);
  and _38233_ (_15667_, _15657_, _09529_);
  and _38234_ (_15668_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _38235_ (_14367_, _15668_, _15667_);
  and _38236_ (_15669_, _15657_, _09532_);
  and _38237_ (_15670_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _38238_ (_14368_, _15670_, _15669_);
  and _38239_ (_15671_, _15657_, _09535_);
  and _38240_ (_15672_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or _38241_ (_14369_, _15672_, _15671_);
  and _38242_ (_15673_, _15657_, _09538_);
  and _38243_ (_15674_, _15659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _38244_ (_14370_, _15674_, _15673_);
  and _38245_ (_15675_, _10103_, _02681_);
  and _38246_ (_15676_, _15675_, _09265_);
  and _38247_ (_15677_, _15676_, _09513_);
  not _38248_ (_15678_, _15676_);
  and _38249_ (_15679_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _38250_ (_14372_, _15679_, _15677_);
  and _38251_ (_15680_, _15676_, _09520_);
  and _38252_ (_15681_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _38253_ (_14373_, _15681_, _15680_);
  and _38254_ (_15682_, _15676_, _09523_);
  and _38255_ (_15683_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _38256_ (_14375_, _15683_, _15682_);
  and _38257_ (_15684_, _15676_, _09526_);
  and _38258_ (_15685_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _38259_ (_14376_, _15685_, _15684_);
  and _38260_ (_15686_, _15676_, _09529_);
  and _38261_ (_15687_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _38262_ (_14377_, _15687_, _15686_);
  and _38263_ (_15688_, _15676_, _09532_);
  and _38264_ (_15689_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _38265_ (_14378_, _15689_, _15688_);
  and _38266_ (_15690_, _15676_, _09535_);
  and _38267_ (_15691_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _38268_ (_14379_, _15691_, _15690_);
  and _38269_ (_15692_, _15676_, _09538_);
  and _38270_ (_15693_, _15678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _38271_ (_14380_, _15693_, _15692_);
  and _38272_ (_15694_, _15675_, _09515_);
  and _38273_ (_15695_, _15694_, _09513_);
  not _38274_ (_15696_, _15694_);
  and _38275_ (_15697_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or _38276_ (_14381_, _15697_, _15695_);
  and _38277_ (_15698_, _15694_, _09520_);
  and _38278_ (_15699_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or _38279_ (_14383_, _15699_, _15698_);
  and _38280_ (_15700_, _15694_, _09523_);
  and _38281_ (_15701_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or _38282_ (_14384_, _15701_, _15700_);
  and _38283_ (_15702_, _15694_, _09526_);
  and _38284_ (_15703_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or _38285_ (_14385_, _15703_, _15702_);
  and _38286_ (_15704_, _15694_, _09529_);
  and _38287_ (_15705_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or _38288_ (_14387_, _15705_, _15704_);
  and _38289_ (_15706_, _15694_, _09532_);
  and _38290_ (_15707_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or _38291_ (_14388_, _15707_, _15706_);
  and _38292_ (_15708_, _15694_, _09535_);
  and _38293_ (_15709_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or _38294_ (_14389_, _15709_, _15708_);
  and _38295_ (_15710_, _15694_, _09538_);
  and _38296_ (_15711_, _15696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or _38297_ (_14390_, _15711_, _15710_);
  and _38298_ (_15712_, _15675_, _09542_);
  and _38299_ (_15713_, _15712_, _09513_);
  not _38300_ (_15714_, _15712_);
  and _38301_ (_15715_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or _38302_ (_14392_, _15715_, _15713_);
  and _38303_ (_15716_, _15712_, _09520_);
  and _38304_ (_15717_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or _38305_ (_14393_, _15717_, _15716_);
  and _38306_ (_15718_, _15712_, _09523_);
  and _38307_ (_15719_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or _38308_ (_14394_, _15719_, _15718_);
  and _38309_ (_15720_, _15712_, _09526_);
  and _38310_ (_15721_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or _38311_ (_14396_, _15721_, _15720_);
  and _38312_ (_15722_, _15712_, _09529_);
  and _38313_ (_15723_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or _38314_ (_14397_, _15723_, _15722_);
  and _38315_ (_15724_, _15712_, _09532_);
  and _38316_ (_15725_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or _38317_ (_14398_, _15725_, _15724_);
  and _38318_ (_15726_, _15712_, _09535_);
  and _38319_ (_15727_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or _38320_ (_14399_, _15727_, _15726_);
  and _38321_ (_15728_, _15712_, _09538_);
  and _38322_ (_15729_, _15714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or _38323_ (_14400_, _15729_, _15728_);
  and _38324_ (_15730_, _15675_, _09562_);
  and _38325_ (_15731_, _15730_, _09513_);
  not _38326_ (_15732_, _15730_);
  and _38327_ (_15733_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _38328_ (_14401_, _15733_, _15731_);
  and _38329_ (_15734_, _15730_, _09520_);
  and _38330_ (_15735_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _38331_ (_14402_, _15735_, _15734_);
  and _38332_ (_15736_, _15730_, _09523_);
  and _38333_ (_15737_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _38334_ (_14404_, _15737_, _15736_);
  and _38335_ (_15738_, _15730_, _09526_);
  and _38336_ (_15739_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _38337_ (_14405_, _15739_, _15738_);
  and _38338_ (_15740_, _15730_, _09529_);
  and _38339_ (_15741_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _38340_ (_14406_, _15741_, _15740_);
  and _38341_ (_15742_, _15730_, _09532_);
  and _38342_ (_15743_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _38343_ (_14408_, _15743_, _15742_);
  and _38344_ (_15744_, _15730_, _09535_);
  and _38345_ (_15745_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _38346_ (_14409_, _15745_, _15744_);
  and _38347_ (_15746_, _15730_, _09538_);
  and _38348_ (_15747_, _15732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _38349_ (_14410_, _15747_, _15746_);
  and _38350_ (_15748_, _15675_, _09582_);
  and _38351_ (_15749_, _15748_, _09513_);
  not _38352_ (_15750_, _15748_);
  and _38353_ (_15751_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _38354_ (_14411_, _15751_, _15749_);
  and _38355_ (_15752_, _15748_, _09520_);
  and _38356_ (_15753_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _38357_ (_14412_, _15753_, _15752_);
  and _38358_ (_15754_, _15748_, _09523_);
  and _38359_ (_15755_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _38360_ (_14413_, _15755_, _15754_);
  and _38361_ (_15756_, _15748_, _09526_);
  and _38362_ (_15757_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _38363_ (_14414_, _15757_, _15756_);
  and _38364_ (_15758_, _15748_, _09529_);
  and _38365_ (_15759_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _38366_ (_14416_, _15759_, _15758_);
  and _38367_ (_15760_, _15748_, _09532_);
  and _38368_ (_15761_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _38369_ (_14417_, _15761_, _15760_);
  and _38370_ (_15762_, _15748_, _09535_);
  and _38371_ (_15763_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _38372_ (_14418_, _15763_, _15762_);
  and _38373_ (_15764_, _15748_, _09538_);
  and _38374_ (_15765_, _15750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _38375_ (_14420_, _15765_, _15764_);
  and _38376_ (_15766_, _15675_, _09601_);
  and _38377_ (_15767_, _15766_, _09513_);
  not _38378_ (_15768_, _15766_);
  and _38379_ (_15769_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or _38380_ (_14421_, _15769_, _15767_);
  and _38381_ (_15770_, _15766_, _09520_);
  and _38382_ (_15771_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or _38383_ (_14422_, _15771_, _15770_);
  and _38384_ (_15772_, _15766_, _09523_);
  and _38385_ (_15773_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or _38386_ (_14423_, _15773_, _15772_);
  and _38387_ (_15774_, _15766_, _09526_);
  and _38388_ (_15775_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or _38389_ (_14424_, _15775_, _15774_);
  and _38390_ (_15776_, _15766_, _09529_);
  and _38391_ (_15777_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or _38392_ (_14425_, _15777_, _15776_);
  and _38393_ (_15778_, _15766_, _09532_);
  and _38394_ (_15779_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or _38395_ (_14426_, _15779_, _15778_);
  and _38396_ (_15780_, _15766_, _09535_);
  and _38397_ (_15781_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or _38398_ (_14428_, _15781_, _15780_);
  and _38399_ (_15782_, _15766_, _09538_);
  and _38400_ (_15783_, _15768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or _38401_ (_14429_, _15783_, _15782_);
  and _38402_ (_15784_, _15675_, _09620_);
  and _38403_ (_15785_, _15784_, _09513_);
  not _38404_ (_15786_, _15784_);
  and _38405_ (_15787_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or _38406_ (_14430_, _15787_, _15785_);
  and _38407_ (_15788_, _15784_, _09520_);
  and _38408_ (_15789_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or _38409_ (_14432_, _15789_, _15788_);
  and _38410_ (_15790_, _15784_, _09523_);
  and _38411_ (_15791_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or _38412_ (_14433_, _15791_, _15790_);
  and _38413_ (_15792_, _15784_, _09526_);
  and _38414_ (_15793_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or _38415_ (_14434_, _15793_, _15792_);
  and _38416_ (_15794_, _15784_, _09529_);
  and _38417_ (_15795_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or _38418_ (_14435_, _15795_, _15794_);
  and _38419_ (_15796_, _15784_, _09532_);
  and _38420_ (_15797_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or _38421_ (_14436_, _15797_, _15796_);
  and _38422_ (_15798_, _15784_, _09535_);
  and _38423_ (_15799_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or _38424_ (_14437_, _15799_, _15798_);
  and _38425_ (_15800_, _15784_, _09538_);
  and _38426_ (_15801_, _15786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or _38427_ (_14438_, _15801_, _15800_);
  and _38428_ (_15802_, _15675_, _09639_);
  and _38429_ (_15803_, _15802_, _09513_);
  not _38430_ (_15804_, _15802_);
  and _38431_ (_15805_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _38432_ (_14440_, _15805_, _15803_);
  and _38433_ (_15806_, _15802_, _09520_);
  and _38434_ (_15807_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _38435_ (_14441_, _15807_, _15806_);
  and _38436_ (_15808_, _15802_, _09523_);
  and _38437_ (_15809_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _38438_ (_14442_, _15809_, _15808_);
  and _38439_ (_15810_, _15802_, _09526_);
  and _38440_ (_15811_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _38441_ (_14444_, _15811_, _15810_);
  and _38442_ (_15812_, _15802_, _09529_);
  and _38443_ (_15813_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _38444_ (_14445_, _15813_, _15812_);
  and _38445_ (_15814_, _15802_, _09532_);
  and _38446_ (_15815_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _38447_ (_14446_, _15815_, _15814_);
  and _38448_ (_15816_, _15802_, _09535_);
  and _38449_ (_15817_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _38450_ (_14447_, _15817_, _15816_);
  and _38451_ (_15818_, _15802_, _09538_);
  and _38452_ (_15819_, _15804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _38453_ (_14448_, _15819_, _15818_);
  and _38454_ (_15820_, _15675_, _09659_);
  and _38455_ (_15821_, _15820_, _09513_);
  not _38456_ (_15822_, _15820_);
  and _38457_ (_15823_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or _38458_ (_14449_, _15823_, _15821_);
  and _38459_ (_15824_, _15820_, _09520_);
  and _38460_ (_15825_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or _38461_ (_14450_, _15825_, _15824_);
  and _38462_ (_15826_, _15820_, _09523_);
  and _38463_ (_15827_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or _38464_ (_14452_, _15827_, _15826_);
  and _38465_ (_15828_, _15820_, _09526_);
  and _38466_ (_15829_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or _38467_ (_14453_, _15829_, _15828_);
  and _38468_ (_15830_, _15820_, _09529_);
  and _38469_ (_15831_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or _38470_ (_14454_, _15831_, _15830_);
  and _38471_ (_15832_, _15820_, _09532_);
  and _38472_ (_15833_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or _38473_ (_14456_, _15833_, _15832_);
  and _38474_ (_15834_, _15820_, _09535_);
  and _38475_ (_15835_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or _38476_ (_14457_, _15835_, _15834_);
  and _38477_ (_15836_, _15820_, _09538_);
  and _38478_ (_15837_, _15822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or _38479_ (_14458_, _15837_, _15836_);
  and _38480_ (_15838_, _15675_, _09678_);
  and _38481_ (_15839_, _15838_, _09513_);
  not _38482_ (_15840_, _15838_);
  and _38483_ (_15841_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _38484_ (_14459_, _15841_, _15839_);
  and _38485_ (_15842_, _15838_, _09520_);
  and _38486_ (_15843_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _38487_ (_14460_, _15843_, _15842_);
  and _38488_ (_15844_, _15838_, _09523_);
  and _38489_ (_15845_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _38490_ (_14461_, _15845_, _15844_);
  and _38491_ (_15846_, _15838_, _09526_);
  and _38492_ (_15847_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _38493_ (_14462_, _15847_, _15846_);
  and _38494_ (_15848_, _15838_, _09529_);
  and _38495_ (_15849_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _38496_ (_14464_, _15849_, _15848_);
  and _38497_ (_15850_, _15838_, _09532_);
  and _38498_ (_15851_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _38499_ (_14465_, _15851_, _15850_);
  and _38500_ (_15852_, _15838_, _09535_);
  and _38501_ (_15853_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _38502_ (_14466_, _15853_, _15852_);
  and _38503_ (_15854_, _15838_, _09538_);
  and _38504_ (_15855_, _15840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _38505_ (_14468_, _15855_, _15854_);
  and _38506_ (_15856_, _15675_, _09697_);
  and _38507_ (_15857_, _15856_, _09513_);
  not _38508_ (_15858_, _15856_);
  and _38509_ (_15859_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _38510_ (_14469_, _15859_, _15857_);
  and _38511_ (_15860_, _15856_, _09520_);
  and _38512_ (_15861_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _38513_ (_14470_, _15861_, _15860_);
  and _38514_ (_15862_, _15856_, _09523_);
  and _38515_ (_15863_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _38516_ (_14471_, _15863_, _15862_);
  and _38517_ (_15864_, _15856_, _09526_);
  and _38518_ (_15865_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _38519_ (_14472_, _15865_, _15864_);
  and _38520_ (_15866_, _15856_, _09529_);
  and _38521_ (_15867_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _38522_ (_14473_, _15867_, _15866_);
  and _38523_ (_15868_, _15856_, _09532_);
  and _38524_ (_15869_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _38525_ (_14474_, _15869_, _15868_);
  and _38526_ (_15870_, _15856_, _09535_);
  and _38527_ (_15871_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _38528_ (_14476_, _15871_, _15870_);
  and _38529_ (_15872_, _15856_, _09538_);
  and _38530_ (_15873_, _15858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _38531_ (_14477_, _15873_, _15872_);
  and _38532_ (_15874_, _15675_, _09716_);
  and _38533_ (_15875_, _15874_, _09513_);
  not _38534_ (_15876_, _15874_);
  and _38535_ (_15877_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or _38536_ (_14478_, _15877_, _15875_);
  and _38537_ (_15878_, _15874_, _09520_);
  and _38538_ (_15879_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or _38539_ (_14480_, _15879_, _15878_);
  and _38540_ (_15880_, _15874_, _09523_);
  and _38541_ (_15881_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or _38542_ (_14481_, _15881_, _15880_);
  and _38543_ (_15882_, _15874_, _09526_);
  and _38544_ (_15883_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or _38545_ (_14482_, _15883_, _15882_);
  and _38546_ (_15884_, _15874_, _09529_);
  and _38547_ (_15885_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or _38548_ (_14483_, _15885_, _15884_);
  and _38549_ (_15886_, _15874_, _09532_);
  and _38550_ (_15887_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or _38551_ (_14484_, _15887_, _15886_);
  and _38552_ (_15888_, _15874_, _09535_);
  and _38553_ (_15889_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or _38554_ (_14485_, _15889_, _15888_);
  and _38555_ (_15890_, _15874_, _09538_);
  and _38556_ (_15891_, _15876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or _38557_ (_14486_, _15891_, _15890_);
  and _38558_ (_15892_, _15675_, _09736_);
  and _38559_ (_15893_, _15892_, _09513_);
  not _38560_ (_15894_, _15892_);
  and _38561_ (_15895_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or _38562_ (_14488_, _15895_, _15893_);
  and _38563_ (_15896_, _15892_, _09520_);
  and _38564_ (_15897_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or _38565_ (_14489_, _15897_, _15896_);
  and _38566_ (_15898_, _15892_, _09523_);
  and _38567_ (_15899_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or _38568_ (_14490_, _15899_, _15898_);
  and _38569_ (_15900_, _15892_, _09526_);
  and _38570_ (_15901_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or _38571_ (_14492_, _15901_, _15900_);
  and _38572_ (_15902_, _15892_, _09529_);
  and _38573_ (_15903_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or _38574_ (_14493_, _15903_, _15902_);
  and _38575_ (_15904_, _15892_, _09532_);
  and _38576_ (_15905_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or _38577_ (_14494_, _15905_, _15904_);
  and _38578_ (_15906_, _15892_, _09535_);
  and _38579_ (_15907_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or _38580_ (_14496_, _15907_, _15906_);
  and _38581_ (_15908_, _15892_, _09538_);
  and _38582_ (_15909_, _15894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or _38583_ (_14497_, _15909_, _15908_);
  and _38584_ (_15910_, _15675_, _09755_);
  and _38585_ (_15911_, _15910_, _09513_);
  not _38586_ (_15912_, _15910_);
  and _38587_ (_15913_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _38588_ (_14498_, _15913_, _15911_);
  and _38589_ (_15914_, _15910_, _09520_);
  and _38590_ (_15915_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _38591_ (_14499_, _15915_, _15914_);
  and _38592_ (_15916_, _15910_, _09523_);
  and _38593_ (_15917_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _38594_ (_14501_, _15917_, _15916_);
  and _38595_ (_15918_, _15910_, _09526_);
  and _38596_ (_15919_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _38597_ (_14502_, _15919_, _15918_);
  and _38598_ (_15920_, _15910_, _09529_);
  and _38599_ (_15921_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _38600_ (_14503_, _15921_, _15920_);
  and _38601_ (_15922_, _15910_, _09532_);
  and _38602_ (_15923_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _38603_ (_14504_, _15923_, _15922_);
  and _38604_ (_15924_, _15910_, _09535_);
  and _38605_ (_15925_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _38606_ (_14505_, _15925_, _15924_);
  and _38607_ (_15926_, _15910_, _09538_);
  and _38608_ (_15927_, _15912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _38609_ (_14506_, _15927_, _15926_);
  and _38610_ (_15928_, _15675_, _09774_);
  and _38611_ (_15929_, _15928_, _09513_);
  not _38612_ (_15930_, _15928_);
  and _38613_ (_15931_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _38614_ (_14508_, _15931_, _15929_);
  and _38615_ (_15932_, _15928_, _09520_);
  and _38616_ (_15933_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _38617_ (_14509_, _15933_, _15932_);
  and _38618_ (_15934_, _15928_, _09523_);
  and _38619_ (_15935_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _38620_ (_14510_, _15935_, _15934_);
  and _38621_ (_15936_, _15928_, _09526_);
  and _38622_ (_15937_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _38623_ (_14511_, _15937_, _15936_);
  and _38624_ (_15938_, _15928_, _09529_);
  and _38625_ (_15939_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _38626_ (_14513_, _15939_, _15938_);
  and _38627_ (_15940_, _15928_, _09532_);
  and _38628_ (_15941_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _38629_ (_14514_, _15941_, _15940_);
  and _38630_ (_15942_, _15928_, _09535_);
  and _38631_ (_15943_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _38632_ (_14515_, _15943_, _15942_);
  and _38633_ (_15944_, _15928_, _09538_);
  and _38634_ (_15945_, _15930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _38635_ (_14516_, _15945_, _15944_);
  and _38636_ (_15946_, _15675_, _09793_);
  and _38637_ (_15947_, _15946_, _09513_);
  not _38638_ (_15948_, _15946_);
  and _38639_ (_15949_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or _38640_ (_14517_, _15949_, _15947_);
  and _38641_ (_15950_, _15946_, _09520_);
  and _38642_ (_15951_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or _38643_ (_14518_, _15951_, _15950_);
  and _38644_ (_15952_, _15946_, _09523_);
  and _38645_ (_15953_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or _38646_ (_14520_, _15953_, _15952_);
  and _38647_ (_15954_, _15946_, _09526_);
  and _38648_ (_15955_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or _38649_ (_14521_, _15955_, _15954_);
  and _38650_ (_15956_, _15946_, _09529_);
  and _38651_ (_15957_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or _38652_ (_14522_, _15957_, _15956_);
  and _38653_ (_15958_, _15946_, _09532_);
  and _38654_ (_15959_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or _38655_ (_14523_, _15959_, _15958_);
  and _38656_ (_15960_, _15946_, _09535_);
  and _38657_ (_15961_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or _38658_ (_14525_, _15961_, _15960_);
  and _38659_ (_15962_, _15946_, _09538_);
  and _38660_ (_15963_, _15948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or _38661_ (_14526_, _15963_, _15962_);
  and _38662_ (_15964_, _10393_, _02681_);
  and _38663_ (_15965_, _15964_, _09265_);
  not _38664_ (_15966_, _15965_);
  and _38665_ (_15967_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _38666_ (_15968_, _15965_, _09513_);
  or _38667_ (_14527_, _15968_, _15967_);
  and _38668_ (_15969_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and _38669_ (_15970_, _15965_, _09520_);
  or _38670_ (_14528_, _15970_, _15969_);
  and _38671_ (_15971_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _38672_ (_15972_, _15965_, _09523_);
  or _38673_ (_14529_, _15972_, _15971_);
  and _38674_ (_15973_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _38675_ (_15974_, _15965_, _09526_);
  or _38676_ (_14530_, _15974_, _15973_);
  and _38677_ (_15975_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _38678_ (_15976_, _15965_, _09529_);
  or _38679_ (_14532_, _15976_, _15975_);
  and _38680_ (_15977_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _38681_ (_15978_, _15965_, _09532_);
  or _38682_ (_14533_, _15978_, _15977_);
  and _38683_ (_15979_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _38684_ (_15980_, _15965_, _09535_);
  or _38685_ (_14534_, _15980_, _15979_);
  and _38686_ (_15981_, _15966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and _38687_ (_15982_, _15965_, _09538_);
  or _38688_ (_14535_, _15982_, _15981_);
  and _38689_ (_15983_, _15964_, _09515_);
  not _38690_ (_15984_, _15983_);
  and _38691_ (_15985_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  and _38692_ (_15986_, _15983_, _09513_);
  or _38693_ (_14537_, _15986_, _15985_);
  and _38694_ (_15987_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  and _38695_ (_15988_, _15983_, _09520_);
  or _38696_ (_14538_, _15988_, _15987_);
  and _38697_ (_15989_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  and _38698_ (_15990_, _15983_, _09523_);
  or _38699_ (_14539_, _15990_, _15989_);
  and _38700_ (_15991_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  and _38701_ (_15992_, _15983_, _09526_);
  or _38702_ (_14540_, _15992_, _15991_);
  and _38703_ (_15993_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  and _38704_ (_15994_, _15983_, _09529_);
  or _38705_ (_14541_, _15994_, _15993_);
  and _38706_ (_15995_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  and _38707_ (_15996_, _15983_, _09532_);
  or _38708_ (_14542_, _15996_, _15995_);
  and _38709_ (_15997_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  and _38710_ (_15998_, _15983_, _09535_);
  or _38711_ (_14544_, _15998_, _15997_);
  and _38712_ (_15999_, _15984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  and _38713_ (_16000_, _15983_, _09538_);
  or _38714_ (_14545_, _16000_, _15999_);
  and _38715_ (_16001_, _15964_, _09542_);
  not _38716_ (_16002_, _16001_);
  and _38717_ (_16003_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  and _38718_ (_16004_, _16001_, _09513_);
  or _38719_ (_14546_, _16004_, _16003_);
  and _38720_ (_16005_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  and _38721_ (_16006_, _16001_, _09520_);
  or _38722_ (_14548_, _16006_, _16005_);
  and _38723_ (_16007_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  and _38724_ (_16008_, _16001_, _09523_);
  or _38725_ (_14549_, _16008_, _16007_);
  and _38726_ (_16009_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  and _38727_ (_16010_, _16001_, _09526_);
  or _38728_ (_14550_, _16010_, _16009_);
  and _38729_ (_16011_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and _38730_ (_16012_, _16001_, _09529_);
  or _38731_ (_14551_, _16012_, _16011_);
  and _38732_ (_16013_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  and _38733_ (_16014_, _16001_, _09532_);
  or _38734_ (_14552_, _16014_, _16013_);
  and _38735_ (_16015_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  and _38736_ (_16016_, _16001_, _09535_);
  or _38737_ (_14553_, _16016_, _16015_);
  and _38738_ (_16017_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and _38739_ (_16018_, _16001_, _09538_);
  or _38740_ (_14554_, _16018_, _16017_);
  and _38741_ (_16019_, _15964_, _09562_);
  not _38742_ (_16020_, _16019_);
  and _38743_ (_16021_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _38744_ (_16022_, _16019_, _09513_);
  or _38745_ (_14556_, _16022_, _16021_);
  and _38746_ (_16023_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _38747_ (_16024_, _16019_, _09520_);
  or _38748_ (_14557_, _16024_, _16023_);
  and _38749_ (_16025_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _38750_ (_16026_, _16019_, _09523_);
  or _38751_ (_14558_, _16026_, _16025_);
  and _38752_ (_16027_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _38753_ (_16028_, _16019_, _09526_);
  or _38754_ (_14560_, _16028_, _16027_);
  and _38755_ (_16029_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _38756_ (_16030_, _16019_, _09529_);
  or _38757_ (_14561_, _16030_, _16029_);
  and _38758_ (_16031_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _38759_ (_16032_, _16019_, _09532_);
  or _38760_ (_14562_, _16032_, _16031_);
  and _38761_ (_16033_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and _38762_ (_16034_, _16019_, _09535_);
  or _38763_ (_14563_, _16034_, _16033_);
  and _38764_ (_16035_, _16020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _38765_ (_16036_, _16019_, _09538_);
  or _38766_ (_14564_, _16036_, _16035_);
  and _38767_ (_16037_, _15964_, _09582_);
  not _38768_ (_16038_, _16037_);
  and _38769_ (_16039_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _38770_ (_16040_, _16037_, _09513_);
  or _38771_ (_14565_, _16040_, _16039_);
  and _38772_ (_16041_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _38773_ (_16042_, _16037_, _09520_);
  or _38774_ (_14566_, _16042_, _16041_);
  and _38775_ (_16043_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _38776_ (_16044_, _16037_, _09523_);
  or _38777_ (_14568_, _16044_, _16043_);
  and _38778_ (_16045_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _38779_ (_16046_, _16037_, _09526_);
  or _38780_ (_14569_, _16046_, _16045_);
  and _38781_ (_16047_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _38782_ (_16048_, _16037_, _09529_);
  or _38783_ (_14570_, _16048_, _16047_);
  and _38784_ (_16049_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and _38785_ (_16050_, _16037_, _09532_);
  or _38786_ (_14572_, _16050_, _16049_);
  and _38787_ (_16051_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _38788_ (_16052_, _16037_, _09535_);
  or _38789_ (_14573_, _16052_, _16051_);
  and _38790_ (_16053_, _16038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and _38791_ (_16054_, _16037_, _09538_);
  or _38792_ (_14574_, _16054_, _16053_);
  and _38793_ (_16055_, _15964_, _09601_);
  not _38794_ (_16056_, _16055_);
  and _38795_ (_16057_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  and _38796_ (_16058_, _16055_, _09513_);
  or _38797_ (_14575_, _16058_, _16057_);
  and _38798_ (_16059_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and _38799_ (_16060_, _16055_, _09520_);
  or _38800_ (_14576_, _16060_, _16059_);
  and _38801_ (_16061_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  and _38802_ (_16062_, _16055_, _09523_);
  or _38803_ (_14577_, _16062_, _16061_);
  and _38804_ (_16063_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and _38805_ (_16064_, _16055_, _09526_);
  or _38806_ (_14578_, _16064_, _16063_);
  and _38807_ (_16065_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and _38808_ (_16066_, _16055_, _09529_);
  or _38809_ (_14580_, _16066_, _16065_);
  and _38810_ (_16067_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and _38811_ (_16068_, _16055_, _09532_);
  or _38812_ (_14581_, _16068_, _16067_);
  and _38813_ (_16069_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and _38814_ (_16070_, _16055_, _09535_);
  or _38815_ (_14582_, _16070_, _16069_);
  and _38816_ (_16071_, _16056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and _38817_ (_16072_, _16055_, _09538_);
  or _38818_ (_14583_, _16072_, _16071_);
  and _38819_ (_16073_, _15964_, _09620_);
  not _38820_ (_16074_, _16073_);
  and _38821_ (_16075_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  and _38822_ (_16076_, _16073_, _09513_);
  or _38823_ (_14585_, _16076_, _16075_);
  and _38824_ (_16077_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  and _38825_ (_16078_, _16073_, _09520_);
  or _38826_ (_14586_, _16078_, _16077_);
  and _38827_ (_16079_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and _38828_ (_16080_, _16073_, _09523_);
  or _38829_ (_14587_, _16080_, _16079_);
  and _38830_ (_16081_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  and _38831_ (_16082_, _16073_, _09526_);
  or _38832_ (_14588_, _16082_, _16081_);
  and _38833_ (_16083_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  and _38834_ (_16084_, _16073_, _09529_);
  or _38835_ (_14589_, _16084_, _16083_);
  and _38836_ (_16085_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  and _38837_ (_16086_, _16073_, _09532_);
  or _38838_ (_14590_, _16086_, _16085_);
  and _38839_ (_16087_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  and _38840_ (_16088_, _16073_, _09535_);
  or _38841_ (_14592_, _16088_, _16087_);
  and _38842_ (_16089_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  and _38843_ (_16090_, _16073_, _09538_);
  or _38844_ (_14593_, _16090_, _16089_);
  and _38845_ (_16091_, _15964_, _09639_);
  not _38846_ (_16092_, _16091_);
  and _38847_ (_16093_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _38848_ (_16094_, _16091_, _09513_);
  or _38849_ (_14594_, _16094_, _16093_);
  and _38850_ (_16095_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _38851_ (_16096_, _16091_, _09520_);
  or _38852_ (_14596_, _16096_, _16095_);
  and _38853_ (_16097_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _38854_ (_16098_, _16091_, _09523_);
  or _38855_ (_14597_, _16098_, _16097_);
  and _38856_ (_16099_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _38857_ (_16100_, _16091_, _09526_);
  or _38858_ (_14598_, _16100_, _16099_);
  and _38859_ (_16101_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _38860_ (_16102_, _16091_, _09529_);
  or _38861_ (_14599_, _16102_, _16101_);
  and _38862_ (_16103_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _38863_ (_16104_, _16091_, _09532_);
  or _38864_ (_14601_, _16104_, _16103_);
  and _38865_ (_16105_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _38866_ (_16106_, _16091_, _09535_);
  or _38867_ (_14602_, _16106_, _16105_);
  and _38868_ (_16107_, _16092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and _38869_ (_16108_, _16091_, _09538_);
  or _38870_ (_14603_, _16108_, _16107_);
  and _38871_ (_16109_, _15964_, _09659_);
  not _38872_ (_16110_, _16109_);
  and _38873_ (_16112_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  and _38874_ (_16113_, _16109_, _09513_);
  or _38875_ (_14605_, _16113_, _16112_);
  and _38876_ (_16114_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  and _38877_ (_16115_, _16109_, _09520_);
  or _38878_ (_14606_, _16115_, _16114_);
  and _38879_ (_16116_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  and _38880_ (_16117_, _16109_, _09523_);
  or _38881_ (_14607_, _16117_, _16116_);
  and _38882_ (_16118_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  and _38883_ (_16120_, _16109_, _09526_);
  or _38884_ (_14608_, _16120_, _16118_);
  and _38885_ (_16121_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  and _38886_ (_16122_, _16109_, _09529_);
  or _38887_ (_14609_, _16122_, _16121_);
  and _38888_ (_16123_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  and _38889_ (_16124_, _16109_, _09532_);
  or _38890_ (_14610_, _16124_, _16123_);
  and _38891_ (_16125_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  and _38892_ (_16126_, _16109_, _09535_);
  or _38893_ (_14611_, _16126_, _16125_);
  and _38894_ (_16128_, _16110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  and _38895_ (_16129_, _16109_, _09538_);
  or _38896_ (_14613_, _16129_, _16128_);
  and _38897_ (_16130_, _15964_, _09678_);
  not _38898_ (_16131_, _16130_);
  and _38899_ (_16132_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _38900_ (_16133_, _16130_, _09513_);
  or _38901_ (_14614_, _16133_, _16132_);
  and _38902_ (_16134_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _38903_ (_16136_, _16130_, _09520_);
  or _38904_ (_14615_, _16136_, _16134_);
  and _38905_ (_16137_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _38906_ (_16138_, _16130_, _09523_);
  or _38907_ (_14617_, _16138_, _16137_);
  and _38908_ (_16139_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _38909_ (_16140_, _16130_, _09526_);
  or _38910_ (_14618_, _16140_, _16139_);
  and _38911_ (_16141_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _38912_ (_16142_, _16130_, _09529_);
  or _38913_ (_14619_, _16142_, _16141_);
  and _38914_ (_16144_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _38915_ (_16145_, _16130_, _09532_);
  or _38916_ (_14620_, _16145_, _16144_);
  and _38917_ (_16146_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and _38918_ (_16147_, _16130_, _09535_);
  or _38919_ (_14621_, _16147_, _16146_);
  and _38920_ (_16148_, _16131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _38921_ (_16149_, _16130_, _09538_);
  or _38922_ (_14622_, _16149_, _16148_);
  and _38923_ (_16151_, _15964_, _09697_);
  not _38924_ (_16152_, _16151_);
  and _38925_ (_16153_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _38926_ (_16154_, _16151_, _09513_);
  or _38927_ (_14623_, _16154_, _16153_);
  and _38928_ (_16155_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and _38929_ (_16156_, _16151_, _09520_);
  or _38930_ (_14625_, _16156_, _16155_);
  and _38931_ (_16157_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _38932_ (_16158_, _16151_, _09523_);
  or _38933_ (_14626_, _16158_, _16157_);
  and _38934_ (_16160_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _38935_ (_16161_, _16151_, _09526_);
  or _38936_ (_14627_, _16161_, _16160_);
  and _38937_ (_16162_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and _38938_ (_16163_, _16151_, _09529_);
  or _38939_ (_14629_, _16163_, _16162_);
  and _38940_ (_16164_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _38941_ (_16165_, _16151_, _09532_);
  or _38942_ (_14630_, _16165_, _16164_);
  and _38943_ (_16167_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _38944_ (_16168_, _16151_, _09535_);
  or _38945_ (_14631_, _16168_, _16167_);
  and _38946_ (_16169_, _16152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and _38947_ (_16170_, _16151_, _09538_);
  or _38948_ (_14632_, _16170_, _16169_);
  and _38949_ (_16171_, _15964_, _09716_);
  not _38950_ (_16172_, _16171_);
  and _38951_ (_16173_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  and _38952_ (_16174_, _16171_, _09513_);
  or _38953_ (_14633_, _16174_, _16173_);
  and _38954_ (_16176_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  and _38955_ (_16177_, _16171_, _09520_);
  or _38956_ (_14634_, _16177_, _16176_);
  and _38957_ (_16178_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  and _38958_ (_16179_, _16171_, _09523_);
  or _38959_ (_14635_, _16179_, _16178_);
  and _38960_ (_16180_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and _38961_ (_16181_, _16171_, _09526_);
  or _38962_ (_14637_, _16181_, _16180_);
  and _38963_ (_16183_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and _38964_ (_16184_, _16171_, _09529_);
  or _38965_ (_14638_, _16184_, _16183_);
  and _38966_ (_16185_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  and _38967_ (_16186_, _16171_, _09532_);
  or _38968_ (_14639_, _16186_, _16185_);
  and _38969_ (_16187_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  and _38970_ (_16188_, _16171_, _09535_);
  or _38971_ (_14641_, _16188_, _16187_);
  and _38972_ (_16189_, _16172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  and _38973_ (_16191_, _16171_, _09538_);
  or _38974_ (_14642_, _16191_, _16189_);
  and _38975_ (_16192_, _15964_, _09736_);
  not _38976_ (_16193_, _16192_);
  and _38977_ (_16194_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and _38978_ (_16195_, _16192_, _09513_);
  or _38979_ (_14643_, _16195_, _16194_);
  and _38980_ (_16196_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  and _38981_ (_16197_, _16192_, _09520_);
  or _38982_ (_14644_, _16197_, _16196_);
  and _38983_ (_16199_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  and _38984_ (_16200_, _16192_, _09523_);
  or _38985_ (_14645_, _16200_, _16199_);
  and _38986_ (_16201_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  and _38987_ (_16202_, _16192_, _09526_);
  or _38988_ (_14646_, _16202_, _16201_);
  and _38989_ (_16203_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  and _38990_ (_16204_, _16192_, _09529_);
  or _38991_ (_14647_, _16204_, _16203_);
  and _38992_ (_16205_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  and _38993_ (_16207_, _16192_, _09532_);
  or _38994_ (_14649_, _16207_, _16205_);
  and _38995_ (_16208_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  and _38996_ (_16209_, _16192_, _09535_);
  or _38997_ (_14650_, _16209_, _16208_);
  and _38998_ (_16210_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  and _38999_ (_16211_, _16192_, _09538_);
  or _39000_ (_14651_, _16211_, _16210_);
  and _39001_ (_16212_, _15964_, _09755_);
  not _39002_ (_16213_, _16212_);
  and _39003_ (_16215_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _39004_ (_16216_, _16212_, _09513_);
  or _39005_ (_14653_, _16216_, _16215_);
  and _39006_ (_16217_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _39007_ (_16218_, _16212_, _09520_);
  or _39008_ (_14654_, _16218_, _16217_);
  and _39009_ (_16219_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _39010_ (_16220_, _16212_, _09523_);
  or _39011_ (_14655_, _16220_, _16219_);
  and _39012_ (_16221_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _39013_ (_16222_, _16212_, _09526_);
  or _39014_ (_14656_, _16222_, _16221_);
  and _39015_ (_16223_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _39016_ (_16224_, _16212_, _09529_);
  or _39017_ (_14657_, _16224_, _16223_);
  and _39018_ (_16225_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _39019_ (_16226_, _16212_, _09532_);
  or _39020_ (_14658_, _16226_, _16225_);
  and _39021_ (_16227_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _39022_ (_16228_, _16212_, _09535_);
  or _39023_ (_14659_, _16228_, _16227_);
  and _39024_ (_16229_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _39025_ (_16230_, _16212_, _09538_);
  or _39026_ (_14661_, _16230_, _16229_);
  and _39027_ (_16231_, _15964_, _09774_);
  not _39028_ (_16232_, _16231_);
  and _39029_ (_16233_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and _39030_ (_16234_, _16231_, _09513_);
  or _39031_ (_14662_, _16234_, _16233_);
  and _39032_ (_16235_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _39033_ (_16236_, _16231_, _09520_);
  or _39034_ (_14663_, _16236_, _16235_);
  and _39035_ (_16237_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _39036_ (_16238_, _16231_, _09523_);
  or _39037_ (_14665_, _16238_, _16237_);
  and _39038_ (_16239_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _39039_ (_16240_, _16231_, _09526_);
  or _39040_ (_14666_, _16240_, _16239_);
  and _39041_ (_16241_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and _39042_ (_16242_, _16231_, _09529_);
  or _39043_ (_14667_, _16242_, _16241_);
  and _39044_ (_16243_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _39045_ (_16244_, _16231_, _09532_);
  or _39046_ (_14668_, _16244_, _16243_);
  and _39047_ (_16245_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _39048_ (_16246_, _16231_, _09535_);
  or _39049_ (_14669_, _16246_, _16245_);
  and _39050_ (_16247_, _16232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _39051_ (_16248_, _16231_, _09538_);
  or _39052_ (_14670_, _16248_, _16247_);
  and _39053_ (_16249_, _15964_, _09793_);
  not _39054_ (_16250_, _16249_);
  and _39055_ (_16251_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  and _39056_ (_16252_, _16249_, _09513_);
  or _39057_ (_14671_, _16252_, _16251_);
  and _39058_ (_16253_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  and _39059_ (_16254_, _16249_, _09520_);
  or _39060_ (_14673_, _16254_, _16253_);
  and _39061_ (_16255_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  and _39062_ (_16256_, _16249_, _09523_);
  or _39063_ (_14674_, _16256_, _16255_);
  and _39064_ (_16257_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  and _39065_ (_16258_, _16249_, _09526_);
  or _39066_ (_14675_, _16258_, _16257_);
  and _39067_ (_16259_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  and _39068_ (_16260_, _16249_, _09529_);
  or _39069_ (_14677_, _16260_, _16259_);
  and _39070_ (_16261_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  and _39071_ (_16262_, _16249_, _09532_);
  or _39072_ (_14678_, _16262_, _16261_);
  and _39073_ (_16263_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  and _39074_ (_16264_, _16249_, _09535_);
  or _39075_ (_14679_, _16264_, _16263_);
  and _39076_ (_16265_, _16250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  and _39077_ (_16266_, _16249_, _09538_);
  or _39078_ (_14680_, _16266_, _16265_);
  and _39079_ (_16267_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and _39080_ (_16268_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _39081_ (_16269_, _16268_, _16267_);
  and _39082_ (_16270_, _16269_, _05996_);
  and _39083_ (_16271_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and _39084_ (_16272_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _39085_ (_16273_, _16272_, _16271_);
  and _39086_ (_16274_, _16273_, _05997_);
  or _39087_ (_16275_, _16274_, _16270_);
  or _39088_ (_16276_, _16275_, _06021_);
  and _39089_ (_16277_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and _39090_ (_16278_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _39091_ (_16279_, _16278_, _16277_);
  and _39092_ (_16280_, _16279_, _05996_);
  and _39093_ (_16281_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and _39094_ (_16282_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _39095_ (_16283_, _16282_, _16281_);
  and _39096_ (_16284_, _16283_, _05997_);
  or _39097_ (_16285_, _16284_, _16280_);
  or _39098_ (_16286_, _16285_, _05920_);
  and _39099_ (_16287_, _16286_, _06033_);
  and _39100_ (_16288_, _16287_, _16276_);
  or _39101_ (_16289_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _39102_ (_16290_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and _39103_ (_16291_, _16290_, _16289_);
  and _39104_ (_16292_, _16291_, _05996_);
  or _39105_ (_16293_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _39106_ (_16294_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and _39107_ (_16295_, _16294_, _16293_);
  and _39108_ (_16296_, _16295_, _05997_);
  or _39109_ (_16297_, _16296_, _16292_);
  or _39110_ (_16298_, _16297_, _06021_);
  or _39111_ (_16299_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _39112_ (_16300_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and _39113_ (_16301_, _16300_, _16299_);
  and _39114_ (_16302_, _16301_, _05996_);
  or _39115_ (_16303_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _39116_ (_16304_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and _39117_ (_16305_, _16304_, _16303_);
  and _39118_ (_16306_, _16305_, _05997_);
  or _39119_ (_16307_, _16306_, _16302_);
  or _39120_ (_16308_, _16307_, _05920_);
  and _39121_ (_16309_, _16308_, _05933_);
  and _39122_ (_16310_, _16309_, _16298_);
  or _39123_ (_16311_, _16310_, _16288_);
  and _39124_ (_16312_, _16311_, _05776_);
  and _39125_ (_16313_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and _39126_ (_16314_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _39127_ (_16315_, _16314_, _16313_);
  and _39128_ (_16316_, _16315_, _05996_);
  and _39129_ (_16317_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and _39130_ (_16318_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _39131_ (_16319_, _16318_, _16317_);
  and _39132_ (_16320_, _16319_, _05997_);
  or _39133_ (_16321_, _16320_, _16316_);
  or _39134_ (_16322_, _16321_, _06021_);
  and _39135_ (_16323_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and _39136_ (_16324_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _39137_ (_16325_, _16324_, _16323_);
  and _39138_ (_16326_, _16325_, _05996_);
  and _39139_ (_16327_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and _39140_ (_16328_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _39141_ (_16329_, _16328_, _16327_);
  and _39142_ (_16330_, _16329_, _05997_);
  or _39143_ (_16331_, _16330_, _16326_);
  or _39144_ (_16332_, _16331_, _05920_);
  and _39145_ (_16333_, _16332_, _06033_);
  and _39146_ (_16334_, _16333_, _16322_);
  or _39147_ (_16335_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _39148_ (_16336_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and _39149_ (_16337_, _16336_, _05997_);
  and _39150_ (_16338_, _16337_, _16335_);
  or _39151_ (_16339_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _39152_ (_16340_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and _39153_ (_16341_, _16340_, _05996_);
  and _39154_ (_16342_, _16341_, _16339_);
  or _39155_ (_16343_, _16342_, _16338_);
  or _39156_ (_16344_, _16343_, _06021_);
  or _39157_ (_16345_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _39158_ (_16346_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and _39159_ (_16347_, _16346_, _05997_);
  and _39160_ (_16348_, _16347_, _16345_);
  or _39161_ (_16349_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _39162_ (_16350_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and _39163_ (_16351_, _16350_, _05996_);
  and _39164_ (_16352_, _16351_, _16349_);
  or _39165_ (_16353_, _16352_, _16348_);
  or _39166_ (_16354_, _16353_, _05920_);
  and _39167_ (_16355_, _16354_, _05933_);
  and _39168_ (_16356_, _16355_, _16344_);
  or _39169_ (_16357_, _16356_, _16334_);
  and _39170_ (_16358_, _16357_, _06071_);
  or _39171_ (_16359_, _16358_, _16312_);
  and _39172_ (_16360_, _16359_, _06070_);
  and _39173_ (_16361_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and _39174_ (_16362_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _39175_ (_16363_, _16362_, _16361_);
  and _39176_ (_16364_, _16363_, _05996_);
  and _39177_ (_16365_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _39178_ (_16366_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _39179_ (_16367_, _16366_, _16365_);
  and _39180_ (_16368_, _16367_, _05997_);
  or _39181_ (_16369_, _16368_, _16364_);
  and _39182_ (_16370_, _16369_, _05920_);
  and _39183_ (_16371_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and _39184_ (_16372_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _39185_ (_16373_, _16372_, _16371_);
  and _39186_ (_16374_, _16373_, _05996_);
  and _39187_ (_16375_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _39188_ (_16376_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _39189_ (_16377_, _16376_, _16375_);
  and _39190_ (_16378_, _16377_, _05997_);
  or _39191_ (_16379_, _16378_, _16374_);
  and _39192_ (_16380_, _16379_, _06021_);
  or _39193_ (_16381_, _16380_, _16370_);
  and _39194_ (_16382_, _16381_, _06033_);
  or _39195_ (_16383_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _39196_ (_16384_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _39197_ (_16385_, _16384_, _05997_);
  and _39198_ (_16386_, _16385_, _16383_);
  or _39199_ (_16387_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _39200_ (_16388_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _39201_ (_16389_, _16388_, _05996_);
  and _39202_ (_16390_, _16389_, _16387_);
  or _39203_ (_16391_, _16390_, _16386_);
  and _39204_ (_16392_, _16391_, _05920_);
  or _39205_ (_16393_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _39206_ (_16394_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _39207_ (_16395_, _16394_, _05997_);
  and _39208_ (_16396_, _16395_, _16393_);
  or _39209_ (_16397_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _39210_ (_16398_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and _39211_ (_16399_, _16398_, _05996_);
  and _39212_ (_16400_, _16399_, _16397_);
  or _39213_ (_16401_, _16400_, _16396_);
  and _39214_ (_16402_, _16401_, _06021_);
  or _39215_ (_16403_, _16402_, _16392_);
  and _39216_ (_16404_, _16403_, _05933_);
  or _39217_ (_16405_, _16404_, _16382_);
  and _39218_ (_16406_, _16405_, _06071_);
  and _39219_ (_16407_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and _39220_ (_16408_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _39221_ (_16409_, _16408_, _16407_);
  and _39222_ (_16410_, _16409_, _05996_);
  and _39223_ (_16411_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and _39224_ (_16412_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _39225_ (_16413_, _16412_, _16411_);
  and _39226_ (_16414_, _16413_, _05997_);
  or _39227_ (_16415_, _16414_, _16410_);
  and _39228_ (_16416_, _16415_, _05920_);
  and _39229_ (_16417_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and _39230_ (_16418_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _39231_ (_16419_, _16418_, _16417_);
  and _39232_ (_16420_, _16419_, _05996_);
  and _39233_ (_16421_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and _39234_ (_16422_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _39235_ (_16423_, _16422_, _16421_);
  and _39236_ (_16424_, _16423_, _05997_);
  or _39237_ (_16425_, _16424_, _16420_);
  and _39238_ (_16426_, _16425_, _06021_);
  or _39239_ (_16427_, _16426_, _16416_);
  and _39240_ (_16428_, _16427_, _06033_);
  or _39241_ (_16429_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _39242_ (_16430_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and _39243_ (_16431_, _16430_, _16429_);
  and _39244_ (_16432_, _16431_, _05996_);
  or _39245_ (_16433_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _39246_ (_16434_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and _39247_ (_16435_, _16434_, _16433_);
  and _39248_ (_16436_, _16435_, _05997_);
  or _39249_ (_16437_, _16436_, _16432_);
  and _39250_ (_16438_, _16437_, _05920_);
  or _39251_ (_16439_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _39252_ (_16440_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and _39253_ (_16441_, _16440_, _16439_);
  and _39254_ (_16442_, _16441_, _05996_);
  or _39255_ (_16443_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _39256_ (_16444_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and _39257_ (_16445_, _16444_, _16443_);
  and _39258_ (_16446_, _16445_, _05997_);
  or _39259_ (_16447_, _16446_, _16442_);
  and _39260_ (_16448_, _16447_, _06021_);
  or _39261_ (_16449_, _16448_, _16438_);
  and _39262_ (_16450_, _16449_, _05933_);
  or _39263_ (_16451_, _16450_, _16428_);
  and _39264_ (_16452_, _16451_, _05776_);
  or _39265_ (_16453_, _16452_, _16406_);
  and _39266_ (_16454_, _16453_, _05822_);
  or _39267_ (_16455_, _16454_, _16360_);
  or _39268_ (_16456_, _16455_, _05868_);
  and _39269_ (_16457_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and _39270_ (_16458_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _39271_ (_16459_, _16458_, _16457_);
  and _39272_ (_16460_, _16459_, _05996_);
  and _39273_ (_16461_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and _39274_ (_16462_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _39275_ (_16463_, _16462_, _16461_);
  and _39276_ (_16464_, _16463_, _05997_);
  or _39277_ (_16465_, _16464_, _16460_);
  or _39278_ (_16466_, _16465_, _06021_);
  and _39279_ (_16467_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and _39280_ (_16468_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _39281_ (_16469_, _16468_, _16467_);
  and _39282_ (_16470_, _16469_, _05996_);
  and _39283_ (_16471_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and _39284_ (_16472_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _39285_ (_16473_, _16472_, _16471_);
  and _39286_ (_16474_, _16473_, _05997_);
  or _39287_ (_16475_, _16474_, _16470_);
  or _39288_ (_16476_, _16475_, _05920_);
  and _39289_ (_16477_, _16476_, _06033_);
  and _39290_ (_16478_, _16477_, _16466_);
  or _39291_ (_16479_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _39292_ (_16480_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and _39293_ (_16481_, _16480_, _05997_);
  and _39294_ (_16482_, _16481_, _16479_);
  or _39295_ (_16483_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _39296_ (_16484_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and _39297_ (_16485_, _16484_, _05996_);
  and _39298_ (_16486_, _16485_, _16483_);
  or _39299_ (_16487_, _16486_, _16482_);
  or _39300_ (_16488_, _16487_, _06021_);
  or _39301_ (_16489_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _39302_ (_16490_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and _39303_ (_16491_, _16490_, _05997_);
  and _39304_ (_16492_, _16491_, _16489_);
  or _39305_ (_16493_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _39306_ (_16494_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and _39307_ (_16495_, _16494_, _05996_);
  and _39308_ (_16496_, _16495_, _16493_);
  or _39309_ (_16497_, _16496_, _16492_);
  or _39310_ (_16498_, _16497_, _05920_);
  and _39311_ (_16499_, _16498_, _05933_);
  and _39312_ (_16500_, _16499_, _16488_);
  or _39313_ (_16501_, _16500_, _16478_);
  and _39314_ (_16502_, _16501_, _06071_);
  and _39315_ (_16503_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and _39316_ (_16504_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _39317_ (_16505_, _16504_, _16503_);
  and _39318_ (_16506_, _16505_, _05996_);
  and _39319_ (_16507_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _39320_ (_16508_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _39321_ (_16509_, _16508_, _16507_);
  and _39322_ (_16510_, _16509_, _05997_);
  or _39323_ (_16511_, _16510_, _16506_);
  or _39324_ (_16512_, _16511_, _06021_);
  and _39325_ (_16513_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and _39326_ (_16514_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _39327_ (_16515_, _16514_, _16513_);
  and _39328_ (_16516_, _16515_, _05996_);
  and _39329_ (_16517_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _39330_ (_16518_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _39331_ (_16519_, _16518_, _16517_);
  and _39332_ (_16520_, _16519_, _05997_);
  or _39333_ (_16521_, _16520_, _16516_);
  or _39334_ (_16522_, _16521_, _05920_);
  and _39335_ (_16523_, _16522_, _06033_);
  and _39336_ (_16524_, _16523_, _16512_);
  or _39337_ (_16525_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _39338_ (_16526_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _39339_ (_16527_, _16526_, _16525_);
  and _39340_ (_16528_, _16527_, _05996_);
  or _39341_ (_16529_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _39342_ (_16530_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and _39343_ (_16531_, _16530_, _16529_);
  and _39344_ (_16532_, _16531_, _05997_);
  or _39345_ (_16533_, _16532_, _16528_);
  or _39346_ (_16534_, _16533_, _06021_);
  or _39347_ (_16535_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _39348_ (_16536_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and _39349_ (_16537_, _16536_, _16535_);
  and _39350_ (_16538_, _16537_, _05996_);
  or _39351_ (_16539_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _39352_ (_16540_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _39353_ (_16541_, _16540_, _16539_);
  and _39354_ (_16542_, _16541_, _05997_);
  or _39355_ (_16543_, _16542_, _16538_);
  or _39356_ (_16544_, _16543_, _05920_);
  and _39357_ (_16545_, _16544_, _05933_);
  and _39358_ (_16546_, _16545_, _16534_);
  or _39359_ (_16547_, _16546_, _16524_);
  and _39360_ (_16548_, _16547_, _05776_);
  or _39361_ (_16549_, _16548_, _16502_);
  and _39362_ (_16550_, _16549_, _06070_);
  or _39363_ (_16551_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _39364_ (_16552_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and _39365_ (_16553_, _16552_, _16551_);
  and _39366_ (_16554_, _16553_, _05996_);
  or _39367_ (_16555_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _39368_ (_16556_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and _39369_ (_16557_, _16556_, _16555_);
  and _39370_ (_16558_, _16557_, _05997_);
  or _39371_ (_16559_, _16558_, _16554_);
  and _39372_ (_16560_, _16559_, _06021_);
  or _39373_ (_16561_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _39374_ (_16562_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and _39375_ (_16563_, _16562_, _16561_);
  and _39376_ (_16564_, _16563_, _05996_);
  or _39377_ (_16565_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _39378_ (_16566_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and _39379_ (_16567_, _16566_, _16565_);
  and _39380_ (_16568_, _16567_, _05997_);
  or _39381_ (_16569_, _16568_, _16564_);
  and _39382_ (_16570_, _16569_, _05920_);
  or _39383_ (_16571_, _16570_, _16560_);
  and _39384_ (_16572_, _16571_, _05933_);
  and _39385_ (_16573_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and _39386_ (_16574_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _39387_ (_16575_, _16574_, _16573_);
  and _39388_ (_16576_, _16575_, _05996_);
  and _39389_ (_16577_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and _39390_ (_16578_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _39391_ (_16579_, _16578_, _16577_);
  and _39392_ (_16580_, _16579_, _05997_);
  or _39393_ (_16581_, _16580_, _16576_);
  and _39394_ (_16582_, _16581_, _06021_);
  and _39395_ (_16583_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and _39396_ (_16584_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _39397_ (_16585_, _16584_, _16583_);
  and _39398_ (_16586_, _16585_, _05996_);
  and _39399_ (_16587_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and _39400_ (_16588_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _39401_ (_16589_, _16588_, _16587_);
  and _39402_ (_16590_, _16589_, _05997_);
  or _39403_ (_16591_, _16590_, _16586_);
  and _39404_ (_16592_, _16591_, _05920_);
  or _39405_ (_16593_, _16592_, _16582_);
  and _39406_ (_16594_, _16593_, _06033_);
  or _39407_ (_16595_, _16594_, _16572_);
  and _39408_ (_16596_, _16595_, _05776_);
  or _39409_ (_16597_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _39410_ (_16598_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and _39411_ (_16599_, _16598_, _05997_);
  and _39412_ (_16600_, _16599_, _16597_);
  or _39413_ (_16601_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _39414_ (_16602_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and _39415_ (_16603_, _16602_, _05996_);
  and _39416_ (_16604_, _16603_, _16601_);
  or _39417_ (_16605_, _16604_, _16600_);
  and _39418_ (_16606_, _16605_, _06021_);
  or _39419_ (_16607_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _39420_ (_16608_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and _39421_ (_16609_, _16608_, _05997_);
  and _39422_ (_16610_, _16609_, _16607_);
  or _39423_ (_16611_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _39424_ (_16612_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and _39425_ (_16613_, _16612_, _05996_);
  and _39426_ (_16614_, _16613_, _16611_);
  or _39427_ (_16615_, _16614_, _16610_);
  and _39428_ (_16616_, _16615_, _05920_);
  or _39429_ (_16617_, _16616_, _16606_);
  and _39430_ (_16618_, _16617_, _05933_);
  and _39431_ (_16619_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and _39432_ (_16620_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _39433_ (_16621_, _16620_, _16619_);
  and _39434_ (_16622_, _16621_, _05996_);
  and _39435_ (_16623_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and _39436_ (_16624_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _39437_ (_16625_, _16624_, _16623_);
  and _39438_ (_16626_, _16625_, _05997_);
  or _39439_ (_16627_, _16626_, _16622_);
  and _39440_ (_16628_, _16627_, _06021_);
  and _39441_ (_16629_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and _39442_ (_16630_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _39443_ (_16631_, _16630_, _16629_);
  and _39444_ (_16632_, _16631_, _05996_);
  and _39445_ (_16633_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _39446_ (_16634_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _39447_ (_16635_, _16634_, _16633_);
  and _39448_ (_16636_, _16635_, _05997_);
  or _39449_ (_16637_, _16636_, _16632_);
  and _39450_ (_16638_, _16637_, _05920_);
  or _39451_ (_16639_, _16638_, _16628_);
  and _39452_ (_16640_, _16639_, _06033_);
  or _39453_ (_16641_, _16640_, _16618_);
  and _39454_ (_16642_, _16641_, _06071_);
  or _39455_ (_16643_, _16642_, _16596_);
  and _39456_ (_16644_, _16643_, _05822_);
  or _39457_ (_16645_, _16644_, _16550_);
  or _39458_ (_16646_, _16645_, _06616_);
  and _39459_ (_16647_, _16646_, _16456_);
  or _39460_ (_16648_, _16647_, _06020_);
  and _39461_ (_16649_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and _39462_ (_16650_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _39463_ (_16651_, _16650_, _16649_);
  and _39464_ (_16652_, _16651_, _05996_);
  and _39465_ (_16653_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and _39466_ (_16654_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _39467_ (_16655_, _16654_, _16653_);
  and _39468_ (_16656_, _16655_, _05997_);
  or _39469_ (_16657_, _16656_, _16652_);
  or _39470_ (_16658_, _16657_, _06021_);
  and _39471_ (_16659_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and _39472_ (_16660_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _39473_ (_16661_, _16660_, _16659_);
  and _39474_ (_16662_, _16661_, _05996_);
  and _39475_ (_16663_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and _39476_ (_16664_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _39477_ (_16665_, _16664_, _16663_);
  and _39478_ (_16666_, _16665_, _05997_);
  or _39479_ (_16667_, _16666_, _16662_);
  or _39480_ (_16668_, _16667_, _05920_);
  and _39481_ (_16669_, _16668_, _06033_);
  and _39482_ (_16670_, _16669_, _16658_);
  or _39483_ (_16671_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _39484_ (_16672_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and _39485_ (_16673_, _16672_, _16671_);
  and _39486_ (_16674_, _16673_, _05996_);
  or _39487_ (_16675_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _39488_ (_16676_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and _39489_ (_16677_, _16676_, _16675_);
  and _39490_ (_16678_, _16677_, _05997_);
  or _39491_ (_16679_, _16678_, _16674_);
  or _39492_ (_16680_, _16679_, _06021_);
  or _39493_ (_16681_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _39494_ (_16682_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and _39495_ (_16683_, _16682_, _16681_);
  and _39496_ (_16684_, _16683_, _05996_);
  or _39497_ (_16685_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _39498_ (_16686_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and _39499_ (_16687_, _16686_, _16685_);
  and _39500_ (_16688_, _16687_, _05997_);
  or _39501_ (_16689_, _16688_, _16684_);
  or _39502_ (_16690_, _16689_, _05920_);
  and _39503_ (_16691_, _16690_, _05933_);
  and _39504_ (_16692_, _16691_, _16680_);
  or _39505_ (_16693_, _16692_, _16670_);
  and _39506_ (_16694_, _16693_, _05776_);
  and _39507_ (_16695_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _39508_ (_16696_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _39509_ (_16697_, _16696_, _16695_);
  and _39510_ (_16698_, _16697_, _05996_);
  and _39511_ (_16699_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _39512_ (_16700_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _39513_ (_16701_, _16700_, _16699_);
  and _39514_ (_16702_, _16701_, _05997_);
  or _39515_ (_16703_, _16702_, _16698_);
  or _39516_ (_16704_, _16703_, _06021_);
  and _39517_ (_16705_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _39518_ (_16706_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or _39519_ (_16707_, _16706_, _16705_);
  and _39520_ (_16708_, _16707_, _05996_);
  and _39521_ (_16709_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _39522_ (_16710_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _39523_ (_16711_, _16710_, _16709_);
  and _39524_ (_16712_, _16711_, _05997_);
  or _39525_ (_16713_, _16712_, _16708_);
  or _39526_ (_16714_, _16713_, _05920_);
  and _39527_ (_16715_, _16714_, _06033_);
  and _39528_ (_16716_, _16715_, _16704_);
  or _39529_ (_16717_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or _39530_ (_16718_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _39531_ (_16719_, _16718_, _05997_);
  and _39532_ (_16720_, _16719_, _16717_);
  or _39533_ (_16721_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _39534_ (_16722_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _39535_ (_16723_, _16722_, _05996_);
  and _39536_ (_16724_, _16723_, _16721_);
  or _39537_ (_16725_, _16724_, _16720_);
  or _39538_ (_16726_, _16725_, _06021_);
  or _39539_ (_16727_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _39540_ (_16728_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _39541_ (_16729_, _16728_, _05997_);
  and _39542_ (_16730_, _16729_, _16727_);
  or _39543_ (_16731_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or _39544_ (_16732_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _39545_ (_16733_, _16732_, _05996_);
  and _39546_ (_16734_, _16733_, _16731_);
  or _39547_ (_16735_, _16734_, _16730_);
  or _39548_ (_16736_, _16735_, _05920_);
  and _39549_ (_16737_, _16736_, _05933_);
  and _39550_ (_16738_, _16737_, _16726_);
  or _39551_ (_16739_, _16738_, _16716_);
  and _39552_ (_16740_, _16739_, _06071_);
  or _39553_ (_16741_, _16740_, _16694_);
  and _39554_ (_16742_, _16741_, _06070_);
  and _39555_ (_16743_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _39556_ (_16744_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or _39557_ (_16745_, _16744_, _16743_);
  and _39558_ (_16746_, _16745_, _05996_);
  and _39559_ (_16747_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _39560_ (_16748_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _39561_ (_16749_, _16748_, _16747_);
  and _39562_ (_16750_, _16749_, _05997_);
  or _39563_ (_16751_, _16750_, _16746_);
  and _39564_ (_16752_, _16751_, _05920_);
  and _39565_ (_16753_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _39566_ (_16754_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or _39567_ (_16755_, _16754_, _16753_);
  and _39568_ (_16756_, _16755_, _05996_);
  and _39569_ (_16757_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _39570_ (_16758_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _39571_ (_16759_, _16758_, _16757_);
  and _39572_ (_16760_, _16759_, _05997_);
  or _39573_ (_16761_, _16760_, _16756_);
  and _39574_ (_16762_, _16761_, _06021_);
  or _39575_ (_16763_, _16762_, _16752_);
  and _39576_ (_16764_, _16763_, _06033_);
  or _39577_ (_16765_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _39578_ (_16766_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _39579_ (_16767_, _16766_, _05997_);
  and _39580_ (_16768_, _16767_, _16765_);
  or _39581_ (_16769_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or _39582_ (_16770_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _39583_ (_16771_, _16770_, _05996_);
  and _39584_ (_16772_, _16771_, _16769_);
  or _39585_ (_16773_, _16772_, _16768_);
  and _39586_ (_16774_, _16773_, _05920_);
  or _39587_ (_16775_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _39588_ (_16776_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _39589_ (_16777_, _16776_, _05997_);
  and _39590_ (_16778_, _16777_, _16775_);
  or _39591_ (_16779_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or _39592_ (_16780_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _39593_ (_16781_, _16780_, _05996_);
  and _39594_ (_16782_, _16781_, _16779_);
  or _39595_ (_16783_, _16782_, _16778_);
  and _39596_ (_16784_, _16783_, _06021_);
  or _39597_ (_16785_, _16784_, _16774_);
  and _39598_ (_16786_, _16785_, _05933_);
  or _39599_ (_16787_, _16786_, _16764_);
  and _39600_ (_16788_, _16787_, _06071_);
  and _39601_ (_16789_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and _39602_ (_16790_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _39603_ (_16791_, _16790_, _16789_);
  and _39604_ (_16792_, _16791_, _05996_);
  and _39605_ (_16793_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and _39606_ (_16794_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _39607_ (_16795_, _16794_, _16793_);
  and _39608_ (_16796_, _16795_, _05997_);
  or _39609_ (_16797_, _16796_, _16792_);
  and _39610_ (_16798_, _16797_, _05920_);
  and _39611_ (_16799_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _39612_ (_16800_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _39613_ (_16801_, _16800_, _16799_);
  and _39614_ (_16802_, _16801_, _05996_);
  and _39615_ (_16803_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and _39616_ (_16804_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _39617_ (_16805_, _16804_, _16803_);
  and _39618_ (_16806_, _16805_, _05997_);
  or _39619_ (_16807_, _16806_, _16802_);
  and _39620_ (_16808_, _16807_, _06021_);
  or _39621_ (_16809_, _16808_, _16798_);
  and _39622_ (_16810_, _16809_, _06033_);
  or _39623_ (_16811_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _39624_ (_16812_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and _39625_ (_16813_, _16812_, _16811_);
  and _39626_ (_16814_, _16813_, _05996_);
  or _39627_ (_16815_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _39628_ (_16816_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and _39629_ (_16817_, _16816_, _16815_);
  and _39630_ (_16818_, _16817_, _05997_);
  or _39631_ (_16819_, _16818_, _16814_);
  and _39632_ (_16820_, _16819_, _05920_);
  or _39633_ (_16821_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _39634_ (_16822_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and _39635_ (_16823_, _16822_, _16821_);
  and _39636_ (_16824_, _16823_, _05996_);
  or _39637_ (_16825_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _39638_ (_16826_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _39639_ (_16827_, _16826_, _16825_);
  and _39640_ (_16828_, _16827_, _05997_);
  or _39641_ (_16829_, _16828_, _16824_);
  and _39642_ (_16830_, _16829_, _06021_);
  or _39643_ (_16831_, _16830_, _16820_);
  and _39644_ (_16832_, _16831_, _05933_);
  or _39645_ (_16833_, _16832_, _16810_);
  and _39646_ (_16834_, _16833_, _05776_);
  or _39647_ (_16835_, _16834_, _16788_);
  and _39648_ (_16836_, _16835_, _05822_);
  or _39649_ (_16837_, _16836_, _16742_);
  or _39650_ (_16838_, _16837_, _05868_);
  and _39651_ (_16839_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and _39652_ (_16840_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _39653_ (_16841_, _16840_, _16839_);
  and _39654_ (_16842_, _16841_, _05996_);
  and _39655_ (_16843_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and _39656_ (_16844_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _39657_ (_16845_, _16844_, _16843_);
  and _39658_ (_16846_, _16845_, _05997_);
  or _39659_ (_16847_, _16846_, _16842_);
  or _39660_ (_16848_, _16847_, _06021_);
  and _39661_ (_16849_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and _39662_ (_16850_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _39663_ (_16851_, _16850_, _16849_);
  and _39664_ (_16852_, _16851_, _05996_);
  and _39665_ (_16853_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and _39666_ (_16854_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _39667_ (_16855_, _16854_, _16853_);
  and _39668_ (_16856_, _16855_, _05997_);
  or _39669_ (_16857_, _16856_, _16852_);
  or _39670_ (_16858_, _16857_, _05920_);
  and _39671_ (_16859_, _16858_, _06033_);
  and _39672_ (_16860_, _16859_, _16848_);
  or _39673_ (_16861_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _39674_ (_16862_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and _39675_ (_16863_, _16862_, _05997_);
  and _39676_ (_16864_, _16863_, _16861_);
  or _39677_ (_16865_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _39678_ (_16866_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and _39679_ (_16867_, _16866_, _05996_);
  and _39680_ (_16868_, _16867_, _16865_);
  or _39681_ (_16869_, _16868_, _16864_);
  or _39682_ (_16870_, _16869_, _06021_);
  or _39683_ (_16871_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _39684_ (_16872_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and _39685_ (_16873_, _16872_, _05997_);
  and _39686_ (_16874_, _16873_, _16871_);
  or _39687_ (_16875_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _39688_ (_16876_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and _39689_ (_16877_, _16876_, _05996_);
  and _39690_ (_16878_, _16877_, _16875_);
  or _39691_ (_16879_, _16878_, _16874_);
  or _39692_ (_16880_, _16879_, _05920_);
  and _39693_ (_16881_, _16880_, _05933_);
  and _39694_ (_16882_, _16881_, _16870_);
  or _39695_ (_16883_, _16882_, _16860_);
  and _39696_ (_16884_, _16883_, _06071_);
  and _39697_ (_16885_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _39698_ (_16886_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or _39699_ (_16887_, _16886_, _16885_);
  and _39700_ (_16888_, _16887_, _05996_);
  and _39701_ (_16889_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _39702_ (_16890_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _39703_ (_16891_, _16890_, _16889_);
  and _39704_ (_16892_, _16891_, _05997_);
  or _39705_ (_16893_, _16892_, _16888_);
  or _39706_ (_16894_, _16893_, _06021_);
  and _39707_ (_16895_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _39708_ (_16896_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or _39709_ (_16897_, _16896_, _16895_);
  and _39710_ (_16898_, _16897_, _05996_);
  and _39711_ (_16899_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _39712_ (_16900_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _39713_ (_16901_, _16900_, _16899_);
  and _39714_ (_16902_, _16901_, _05997_);
  or _39715_ (_16903_, _16902_, _16898_);
  or _39716_ (_16904_, _16903_, _05920_);
  and _39717_ (_16905_, _16904_, _06033_);
  and _39718_ (_16906_, _16905_, _16894_);
  or _39719_ (_16907_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or _39720_ (_16908_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _39721_ (_16909_, _16908_, _16907_);
  and _39722_ (_16910_, _16909_, _05996_);
  or _39723_ (_16911_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _39724_ (_16912_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _39725_ (_16913_, _16912_, _16911_);
  and _39726_ (_16914_, _16913_, _05997_);
  or _39727_ (_16915_, _16914_, _16910_);
  or _39728_ (_16916_, _16915_, _06021_);
  or _39729_ (_16917_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or _39730_ (_16918_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _39731_ (_16919_, _16918_, _16917_);
  and _39732_ (_16920_, _16919_, _05996_);
  or _39733_ (_16921_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _39734_ (_16922_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and _39735_ (_16923_, _16922_, _16921_);
  and _39736_ (_16924_, _16923_, _05997_);
  or _39737_ (_16925_, _16924_, _16920_);
  or _39738_ (_16926_, _16925_, _05920_);
  and _39739_ (_16927_, _16926_, _05933_);
  and _39740_ (_16928_, _16927_, _16916_);
  or _39741_ (_16929_, _16928_, _16906_);
  and _39742_ (_16930_, _16929_, _05776_);
  or _39743_ (_16931_, _16930_, _16884_);
  and _39744_ (_16932_, _16931_, _06070_);
  or _39745_ (_16933_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _39746_ (_16934_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _39747_ (_16935_, _16934_, _16933_);
  and _39748_ (_16936_, _16935_, _05996_);
  or _39749_ (_16937_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or _39750_ (_16938_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _39751_ (_16939_, _16938_, _16937_);
  and _39752_ (_16940_, _16939_, _05997_);
  or _39753_ (_16941_, _16940_, _16936_);
  and _39754_ (_16942_, _16941_, _06021_);
  or _39755_ (_16943_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _39756_ (_16944_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _39757_ (_16945_, _16944_, _16943_);
  and _39758_ (_16946_, _16945_, _05996_);
  or _39759_ (_16947_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or _39760_ (_16948_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _39761_ (_16949_, _16948_, _16947_);
  and _39762_ (_16950_, _16949_, _05997_);
  or _39763_ (_16951_, _16950_, _16946_);
  and _39764_ (_16952_, _16951_, _05920_);
  or _39765_ (_16953_, _16952_, _16942_);
  and _39766_ (_16954_, _16953_, _05933_);
  and _39767_ (_16955_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _39768_ (_16956_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or _39769_ (_16957_, _16956_, _16955_);
  and _39770_ (_16958_, _16957_, _05996_);
  and _39771_ (_16959_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _39772_ (_16960_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _39773_ (_16961_, _16960_, _16959_);
  and _39774_ (_16962_, _16961_, _05997_);
  or _39775_ (_16963_, _16962_, _16958_);
  and _39776_ (_16964_, _16963_, _06021_);
  and _39777_ (_16965_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _39778_ (_16966_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _39779_ (_16967_, _16966_, _16965_);
  and _39780_ (_16968_, _16967_, _05996_);
  and _39781_ (_16969_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _39782_ (_16970_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or _39783_ (_16971_, _16970_, _16969_);
  and _39784_ (_16972_, _16971_, _05997_);
  or _39785_ (_16973_, _16972_, _16968_);
  and _39786_ (_16974_, _16973_, _05920_);
  or _39787_ (_16975_, _16974_, _16964_);
  and _39788_ (_16976_, _16975_, _06033_);
  or _39789_ (_16977_, _16976_, _16954_);
  and _39790_ (_16978_, _16977_, _05776_);
  or _39791_ (_16979_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or _39792_ (_16980_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and _39793_ (_16981_, _16980_, _05997_);
  and _39794_ (_16982_, _16981_, _16979_);
  or _39795_ (_16983_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or _39796_ (_16984_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and _39797_ (_16985_, _16984_, _05996_);
  and _39798_ (_16986_, _16985_, _16983_);
  or _39799_ (_16987_, _16986_, _16982_);
  and _39800_ (_16988_, _16987_, _06021_);
  or _39801_ (_16989_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or _39802_ (_16990_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and _39803_ (_16991_, _16990_, _05997_);
  and _39804_ (_16992_, _16991_, _16989_);
  or _39805_ (_16993_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or _39806_ (_16994_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and _39807_ (_16995_, _16994_, _05996_);
  and _39808_ (_16996_, _16995_, _16993_);
  or _39809_ (_16997_, _16996_, _16992_);
  and _39810_ (_16998_, _16997_, _05920_);
  or _39811_ (_16999_, _16998_, _16988_);
  and _39812_ (_17000_, _16999_, _05933_);
  and _39813_ (_17001_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and _39814_ (_17002_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or _39815_ (_17003_, _17002_, _17001_);
  and _39816_ (_17004_, _17003_, _05996_);
  and _39817_ (_17005_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and _39818_ (_17006_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or _39819_ (_17007_, _17006_, _17005_);
  and _39820_ (_17008_, _17007_, _05997_);
  or _39821_ (_17009_, _17008_, _17004_);
  and _39822_ (_17010_, _17009_, _06021_);
  and _39823_ (_17011_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and _39824_ (_17012_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or _39825_ (_17013_, _17012_, _17011_);
  and _39826_ (_17014_, _17013_, _05996_);
  and _39827_ (_17015_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and _39828_ (_17016_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or _39829_ (_17017_, _17016_, _17015_);
  and _39830_ (_17018_, _17017_, _05997_);
  or _39831_ (_17019_, _17018_, _17014_);
  and _39832_ (_17020_, _17019_, _05920_);
  or _39833_ (_17021_, _17020_, _17010_);
  and _39834_ (_17022_, _17021_, _06033_);
  or _39835_ (_17023_, _17022_, _17000_);
  and _39836_ (_17024_, _17023_, _06071_);
  or _39837_ (_17025_, _17024_, _16978_);
  and _39838_ (_17026_, _17025_, _05822_);
  or _39839_ (_17027_, _17026_, _16932_);
  or _39840_ (_17028_, _17027_, _06616_);
  and _39841_ (_17029_, _17028_, _16838_);
  or _39842_ (_17030_, _17029_, _05584_);
  and _39843_ (_17031_, _17030_, _16648_);
  or _39844_ (_17032_, _17031_, _06019_);
  or _39845_ (_17033_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _39846_ (_17034_, _17033_, _25365_);
  and _39847_ (_14803_, _17034_, _17032_);
  and _39848_ (_17035_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and _39849_ (_17036_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _39850_ (_17037_, _17036_, _17035_);
  and _39851_ (_17038_, _17037_, _05997_);
  and _39852_ (_17039_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and _39853_ (_17040_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _39854_ (_17041_, _17040_, _17039_);
  and _39855_ (_17042_, _17041_, _05996_);
  or _39856_ (_17043_, _17042_, _17038_);
  or _39857_ (_17044_, _17043_, _06021_);
  and _39858_ (_17045_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and _39859_ (_17046_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _39860_ (_17047_, _17046_, _17045_);
  and _39861_ (_17048_, _17047_, _05997_);
  and _39862_ (_17049_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and _39863_ (_17050_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _39864_ (_17051_, _17050_, _17049_);
  and _39865_ (_17052_, _17051_, _05996_);
  or _39866_ (_17053_, _17052_, _17048_);
  or _39867_ (_17054_, _17053_, _05920_);
  and _39868_ (_17055_, _17054_, _06033_);
  and _39869_ (_17056_, _17055_, _17044_);
  or _39870_ (_17057_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _39871_ (_17058_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and _39872_ (_17059_, _17058_, _05996_);
  and _39873_ (_17060_, _17059_, _17057_);
  or _39874_ (_17061_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _39875_ (_17062_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and _39876_ (_17063_, _17062_, _05997_);
  and _39877_ (_17064_, _17063_, _17061_);
  or _39878_ (_17065_, _17064_, _17060_);
  or _39879_ (_17066_, _17065_, _06021_);
  or _39880_ (_17067_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _39881_ (_17068_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and _39882_ (_17069_, _17068_, _05996_);
  and _39883_ (_17070_, _17069_, _17067_);
  or _39884_ (_17071_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _39885_ (_17072_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and _39886_ (_17073_, _17072_, _05997_);
  and _39887_ (_17074_, _17073_, _17071_);
  or _39888_ (_17075_, _17074_, _17070_);
  or _39889_ (_17076_, _17075_, _05920_);
  and _39890_ (_17077_, _17076_, _05933_);
  and _39891_ (_17078_, _17077_, _17066_);
  or _39892_ (_17079_, _17078_, _17056_);
  or _39893_ (_17080_, _17079_, _05776_);
  and _39894_ (_17081_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and _39895_ (_17082_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _39896_ (_17083_, _17082_, _05996_);
  or _39897_ (_17084_, _17083_, _17081_);
  and _39898_ (_17085_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _39899_ (_17086_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _39900_ (_17087_, _17086_, _05997_);
  or _39901_ (_17088_, _17087_, _17085_);
  and _39902_ (_17089_, _17088_, _17084_);
  or _39903_ (_17090_, _17089_, _06021_);
  and _39904_ (_17091_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and _39905_ (_17092_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _39906_ (_17093_, _17092_, _05996_);
  or _39907_ (_17094_, _17093_, _17091_);
  and _39908_ (_17095_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and _39909_ (_17096_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _39910_ (_17097_, _17096_, _05997_);
  or _39911_ (_17098_, _17097_, _17095_);
  and _39912_ (_17099_, _17098_, _17094_);
  or _39913_ (_17100_, _17099_, _05920_);
  and _39914_ (_17101_, _17100_, _06033_);
  and _39915_ (_17102_, _17101_, _17090_);
  or _39916_ (_17103_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _39917_ (_17104_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and _39918_ (_17105_, _17104_, _17103_);
  or _39919_ (_17106_, _17105_, _05997_);
  or _39920_ (_17107_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _39921_ (_17108_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and _39922_ (_17109_, _17108_, _17107_);
  or _39923_ (_17110_, _17109_, _05996_);
  and _39924_ (_17111_, _17110_, _17106_);
  or _39925_ (_17112_, _17111_, _06021_);
  or _39926_ (_17113_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _39927_ (_17114_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and _39928_ (_17115_, _17114_, _17113_);
  or _39929_ (_17116_, _17115_, _05997_);
  or _39930_ (_17117_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _39931_ (_17118_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and _39932_ (_17119_, _17118_, _17117_);
  or _39933_ (_17120_, _17119_, _05996_);
  and _39934_ (_17121_, _17120_, _17116_);
  or _39935_ (_17122_, _17121_, _05920_);
  and _39936_ (_17123_, _17122_, _05933_);
  and _39937_ (_17124_, _17123_, _17112_);
  or _39938_ (_17125_, _17124_, _17102_);
  or _39939_ (_17126_, _17125_, _06071_);
  and _39940_ (_17127_, _17126_, _06070_);
  and _39941_ (_17128_, _17127_, _17080_);
  and _39942_ (_17129_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _39943_ (_17130_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _39944_ (_17131_, _17130_, _17129_);
  and _39945_ (_17132_, _17131_, _05996_);
  and _39946_ (_17133_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and _39947_ (_17134_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _39948_ (_17135_, _17134_, _17133_);
  and _39949_ (_17136_, _17135_, _05997_);
  or _39950_ (_17137_, _17136_, _17132_);
  and _39951_ (_17138_, _17137_, _05920_);
  and _39952_ (_17139_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and _39953_ (_17140_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _39954_ (_17141_, _17140_, _17139_);
  and _39955_ (_17142_, _17141_, _05996_);
  and _39956_ (_17143_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _39957_ (_17144_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _39958_ (_17145_, _17144_, _17143_);
  and _39959_ (_17146_, _17145_, _05997_);
  or _39960_ (_17147_, _17146_, _17142_);
  and _39961_ (_17148_, _17147_, _06021_);
  or _39962_ (_17149_, _17148_, _17138_);
  and _39963_ (_17150_, _17149_, _06033_);
  or _39964_ (_17151_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _39965_ (_17152_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _39966_ (_17153_, _17152_, _17151_);
  and _39967_ (_17154_, _17153_, _05996_);
  or _39968_ (_17155_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _39969_ (_17156_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _39970_ (_17157_, _17156_, _17155_);
  and _39971_ (_17158_, _17157_, _05997_);
  or _39972_ (_17159_, _17158_, _17154_);
  and _39973_ (_17160_, _17159_, _05920_);
  or _39974_ (_17161_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _39975_ (_17162_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _39976_ (_17163_, _17162_, _17161_);
  and _39977_ (_17164_, _17163_, _05996_);
  or _39978_ (_17165_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _39979_ (_17166_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _39980_ (_17167_, _17166_, _17165_);
  and _39981_ (_17168_, _17167_, _05997_);
  or _39982_ (_17169_, _17168_, _17164_);
  and _39983_ (_17170_, _17169_, _06021_);
  or _39984_ (_17171_, _17170_, _17160_);
  and _39985_ (_17172_, _17171_, _05933_);
  or _39986_ (_17173_, _17172_, _17150_);
  and _39987_ (_17174_, _17173_, _06071_);
  and _39988_ (_17175_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and _39989_ (_17176_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _39990_ (_17177_, _17176_, _17175_);
  and _39991_ (_17178_, _17177_, _05996_);
  and _39992_ (_17179_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and _39993_ (_17180_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _39994_ (_17181_, _17180_, _17179_);
  and _39995_ (_17182_, _17181_, _05997_);
  or _39996_ (_17183_, _17182_, _17178_);
  and _39997_ (_17184_, _17183_, _05920_);
  and _39998_ (_17185_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and _39999_ (_17186_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _40000_ (_17187_, _17186_, _17185_);
  and _40001_ (_17188_, _17187_, _05996_);
  and _40002_ (_17189_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and _40003_ (_17190_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _40004_ (_17191_, _17190_, _17189_);
  and _40005_ (_17192_, _17191_, _05997_);
  or _40006_ (_17193_, _17192_, _17188_);
  and _40007_ (_17194_, _17193_, _06021_);
  or _40008_ (_17195_, _17194_, _17184_);
  and _40009_ (_17196_, _17195_, _06033_);
  or _40010_ (_17197_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _40011_ (_17198_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and _40012_ (_17199_, _17198_, _17197_);
  and _40013_ (_17200_, _17199_, _05996_);
  or _40014_ (_17201_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _40015_ (_17202_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and _40016_ (_17203_, _17202_, _17201_);
  and _40017_ (_17204_, _17203_, _05997_);
  or _40018_ (_17205_, _17204_, _17200_);
  and _40019_ (_17206_, _17205_, _05920_);
  or _40020_ (_17207_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _40021_ (_17208_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and _40022_ (_17209_, _17208_, _17207_);
  and _40023_ (_17210_, _17209_, _05996_);
  or _40024_ (_17211_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _40025_ (_17212_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and _40026_ (_17213_, _17212_, _17211_);
  and _40027_ (_17214_, _17213_, _05997_);
  or _40028_ (_17215_, _17214_, _17210_);
  and _40029_ (_17216_, _17215_, _06021_);
  or _40030_ (_17217_, _17216_, _17206_);
  and _40031_ (_17218_, _17217_, _05933_);
  or _40032_ (_17219_, _17218_, _17196_);
  and _40033_ (_17220_, _17219_, _05776_);
  or _40034_ (_17221_, _17220_, _17174_);
  and _40035_ (_17222_, _17221_, _05822_);
  or _40036_ (_17223_, _17222_, _17128_);
  or _40037_ (_17224_, _17223_, _05868_);
  and _40038_ (_17225_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and _40039_ (_17226_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _40040_ (_17227_, _17226_, _17225_);
  and _40041_ (_17228_, _17227_, _05996_);
  and _40042_ (_17229_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and _40043_ (_17230_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _40044_ (_17231_, _17230_, _17229_);
  and _40045_ (_17232_, _17231_, _05997_);
  or _40046_ (_17233_, _17232_, _17228_);
  or _40047_ (_17234_, _17233_, _06021_);
  and _40048_ (_17235_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and _40049_ (_17236_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _40050_ (_17237_, _17236_, _17235_);
  and _40051_ (_17238_, _17237_, _05996_);
  and _40052_ (_17239_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and _40053_ (_17240_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _40054_ (_17241_, _17240_, _17239_);
  and _40055_ (_17242_, _17241_, _05997_);
  or _40056_ (_17243_, _17242_, _17238_);
  or _40057_ (_17244_, _17243_, _05920_);
  and _40058_ (_17245_, _17244_, _06033_);
  and _40059_ (_17246_, _17245_, _17234_);
  or _40060_ (_17247_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _40061_ (_17248_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and _40062_ (_17249_, _17248_, _05997_);
  and _40063_ (_17250_, _17249_, _17247_);
  or _40064_ (_17251_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _40065_ (_17252_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and _40066_ (_17253_, _17252_, _05996_);
  and _40067_ (_17254_, _17253_, _17251_);
  or _40068_ (_17255_, _17254_, _17250_);
  or _40069_ (_17256_, _17255_, _06021_);
  or _40070_ (_17257_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _40071_ (_17258_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and _40072_ (_17259_, _17258_, _05997_);
  and _40073_ (_17260_, _17259_, _17257_);
  or _40074_ (_17261_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _40075_ (_17262_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and _40076_ (_17263_, _17262_, _05996_);
  and _40077_ (_17264_, _17263_, _17261_);
  or _40078_ (_17265_, _17264_, _17260_);
  or _40079_ (_17266_, _17265_, _05920_);
  and _40080_ (_17267_, _17266_, _05933_);
  and _40081_ (_17268_, _17267_, _17256_);
  or _40082_ (_17269_, _17268_, _17246_);
  and _40083_ (_17270_, _17269_, _06071_);
  and _40084_ (_17271_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and _40085_ (_17272_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _40086_ (_17273_, _17272_, _17271_);
  and _40087_ (_17274_, _17273_, _05996_);
  and _40088_ (_17275_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and _40089_ (_17276_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _40090_ (_17277_, _17276_, _17275_);
  and _40091_ (_17278_, _17277_, _05997_);
  or _40092_ (_17279_, _17278_, _17274_);
  or _40093_ (_17280_, _17279_, _06021_);
  and _40094_ (_17281_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and _40095_ (_17282_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _40096_ (_17283_, _17282_, _17281_);
  and _40097_ (_17284_, _17283_, _05996_);
  and _40098_ (_17285_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and _40099_ (_17286_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _40100_ (_17287_, _17286_, _17285_);
  and _40101_ (_17288_, _17287_, _05997_);
  or _40102_ (_17289_, _17288_, _17284_);
  or _40103_ (_17290_, _17289_, _05920_);
  and _40104_ (_17291_, _17290_, _06033_);
  and _40105_ (_17292_, _17291_, _17280_);
  or _40106_ (_17293_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _40107_ (_17294_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and _40108_ (_17295_, _17294_, _17293_);
  and _40109_ (_17296_, _17295_, _05996_);
  or _40110_ (_17297_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _40111_ (_17298_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and _40112_ (_17299_, _17298_, _17297_);
  and _40113_ (_17300_, _17299_, _05997_);
  or _40114_ (_17301_, _17300_, _17296_);
  or _40115_ (_17302_, _17301_, _06021_);
  or _40116_ (_17303_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _40117_ (_17304_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and _40118_ (_17305_, _17304_, _17303_);
  and _40119_ (_17306_, _17305_, _05996_);
  or _40120_ (_17307_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _40121_ (_17308_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and _40122_ (_17309_, _17308_, _17307_);
  and _40123_ (_17310_, _17309_, _05997_);
  or _40124_ (_17311_, _17310_, _17306_);
  or _40125_ (_17312_, _17311_, _05920_);
  and _40126_ (_17313_, _17312_, _05933_);
  and _40127_ (_17314_, _17313_, _17302_);
  or _40128_ (_17315_, _17314_, _17292_);
  and _40129_ (_17316_, _17315_, _05776_);
  or _40130_ (_17317_, _17316_, _17270_);
  and _40131_ (_17318_, _17317_, _06070_);
  or _40132_ (_17319_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _40133_ (_17320_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and _40134_ (_17321_, _17320_, _17319_);
  and _40135_ (_17322_, _17321_, _05996_);
  or _40136_ (_17323_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _40137_ (_17324_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and _40138_ (_17325_, _17324_, _17323_);
  and _40139_ (_17326_, _17325_, _05997_);
  or _40140_ (_17327_, _17326_, _17322_);
  and _40141_ (_17328_, _17327_, _06021_);
  or _40142_ (_17329_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _40143_ (_17330_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and _40144_ (_17331_, _17330_, _17329_);
  and _40145_ (_17332_, _17331_, _05996_);
  or _40146_ (_17333_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _40147_ (_17334_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and _40148_ (_17335_, _17334_, _17333_);
  and _40149_ (_17336_, _17335_, _05997_);
  or _40150_ (_17337_, _17336_, _17332_);
  and _40151_ (_17338_, _17337_, _05920_);
  or _40152_ (_17339_, _17338_, _17328_);
  and _40153_ (_17340_, _17339_, _05933_);
  and _40154_ (_17341_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and _40155_ (_17342_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _40156_ (_17343_, _17342_, _17341_);
  and _40157_ (_17344_, _17343_, _05996_);
  and _40158_ (_17345_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and _40159_ (_17346_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _40160_ (_17347_, _17346_, _17345_);
  and _40161_ (_17348_, _17347_, _05997_);
  or _40162_ (_17349_, _17348_, _17344_);
  and _40163_ (_17350_, _17349_, _06021_);
  and _40164_ (_17351_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and _40165_ (_17352_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _40166_ (_17353_, _17352_, _17351_);
  and _40167_ (_17354_, _17353_, _05996_);
  and _40168_ (_17355_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and _40169_ (_17356_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _40170_ (_17357_, _17356_, _17355_);
  and _40171_ (_17358_, _17357_, _05997_);
  or _40172_ (_17359_, _17358_, _17354_);
  and _40173_ (_17360_, _17359_, _05920_);
  or _40174_ (_17361_, _17360_, _17350_);
  and _40175_ (_17362_, _17361_, _06033_);
  or _40176_ (_17363_, _17362_, _17340_);
  and _40177_ (_17364_, _17363_, _05776_);
  or _40178_ (_17365_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or _40179_ (_17366_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and _40180_ (_17367_, _17366_, _05997_);
  and _40181_ (_17368_, _17367_, _17365_);
  or _40182_ (_17369_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or _40183_ (_17370_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and _40184_ (_17371_, _17370_, _05996_);
  and _40185_ (_17372_, _17371_, _17369_);
  or _40186_ (_17373_, _17372_, _17368_);
  and _40187_ (_17374_, _17373_, _06021_);
  or _40188_ (_17375_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or _40189_ (_17376_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and _40190_ (_17377_, _17376_, _05997_);
  and _40191_ (_17378_, _17377_, _17375_);
  or _40192_ (_17379_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or _40193_ (_17380_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and _40194_ (_17381_, _17380_, _05996_);
  and _40195_ (_17382_, _17381_, _17379_);
  or _40196_ (_17383_, _17382_, _17378_);
  and _40197_ (_17384_, _17383_, _05920_);
  or _40198_ (_17385_, _17384_, _17374_);
  and _40199_ (_17386_, _17385_, _05933_);
  and _40200_ (_17387_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and _40201_ (_17388_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or _40202_ (_17389_, _17388_, _17387_);
  and _40203_ (_17390_, _17389_, _05996_);
  and _40204_ (_17391_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and _40205_ (_17392_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or _40206_ (_17393_, _17392_, _17391_);
  and _40207_ (_17394_, _17393_, _05997_);
  or _40208_ (_17395_, _17394_, _17390_);
  and _40209_ (_17396_, _17395_, _06021_);
  and _40210_ (_17397_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and _40211_ (_17398_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or _40212_ (_17399_, _17398_, _17397_);
  and _40213_ (_17400_, _17399_, _05996_);
  and _40214_ (_17401_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and _40215_ (_17402_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or _40216_ (_17403_, _17402_, _17401_);
  and _40217_ (_17404_, _17403_, _05997_);
  or _40218_ (_17405_, _17404_, _17400_);
  and _40219_ (_17406_, _17405_, _05920_);
  or _40220_ (_17407_, _17406_, _17396_);
  and _40221_ (_17408_, _17407_, _06033_);
  or _40222_ (_17409_, _17408_, _17386_);
  and _40223_ (_17410_, _17409_, _06071_);
  or _40224_ (_17411_, _17410_, _17364_);
  and _40225_ (_17412_, _17411_, _05822_);
  or _40226_ (_17413_, _17412_, _17318_);
  or _40227_ (_17414_, _17413_, _06616_);
  and _40228_ (_17415_, _17414_, _17224_);
  or _40229_ (_17416_, _17415_, _06020_);
  and _40230_ (_17417_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and _40231_ (_17418_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _40232_ (_17419_, _17418_, _17417_);
  and _40233_ (_17420_, _17419_, _05996_);
  and _40234_ (_17421_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and _40235_ (_17422_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _40236_ (_17423_, _17422_, _17421_);
  and _40237_ (_17424_, _17423_, _05997_);
  or _40238_ (_17425_, _17424_, _17420_);
  or _40239_ (_17426_, _17425_, _06021_);
  and _40240_ (_17427_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and _40241_ (_17428_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _40242_ (_17429_, _17428_, _17427_);
  and _40243_ (_17430_, _17429_, _05996_);
  and _40244_ (_17431_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and _40245_ (_17432_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _40246_ (_17433_, _17432_, _17431_);
  and _40247_ (_17434_, _17433_, _05997_);
  or _40248_ (_17435_, _17434_, _17430_);
  or _40249_ (_17436_, _17435_, _05920_);
  and _40250_ (_17437_, _17436_, _06033_);
  and _40251_ (_17438_, _17437_, _17426_);
  or _40252_ (_17439_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _40253_ (_17440_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and _40254_ (_17441_, _17440_, _17439_);
  and _40255_ (_17442_, _17441_, _05996_);
  or _40256_ (_17443_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _40257_ (_17444_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and _40258_ (_17445_, _17444_, _17443_);
  and _40259_ (_17446_, _17445_, _05997_);
  or _40260_ (_17447_, _17446_, _17442_);
  or _40261_ (_17448_, _17447_, _06021_);
  or _40262_ (_17449_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _40263_ (_17450_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and _40264_ (_17451_, _17450_, _17449_);
  and _40265_ (_17452_, _17451_, _05996_);
  or _40266_ (_17453_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _40267_ (_17454_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and _40268_ (_17455_, _17454_, _17453_);
  and _40269_ (_17456_, _17455_, _05997_);
  or _40270_ (_17457_, _17456_, _17452_);
  or _40271_ (_17458_, _17457_, _05920_);
  and _40272_ (_17459_, _17458_, _05933_);
  and _40273_ (_17460_, _17459_, _17448_);
  or _40274_ (_17461_, _17460_, _17438_);
  and _40275_ (_17462_, _17461_, _05776_);
  and _40276_ (_17463_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and _40277_ (_17464_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or _40278_ (_17465_, _17464_, _17463_);
  and _40279_ (_17466_, _17465_, _05996_);
  and _40280_ (_17467_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _40281_ (_17468_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or _40282_ (_17469_, _17468_, _17467_);
  and _40283_ (_17470_, _17469_, _05997_);
  or _40284_ (_17471_, _17470_, _17466_);
  or _40285_ (_17472_, _17471_, _06021_);
  and _40286_ (_17473_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _40287_ (_17474_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _40288_ (_17475_, _17474_, _17473_);
  and _40289_ (_17476_, _17475_, _05996_);
  and _40290_ (_17477_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _40291_ (_17478_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _40292_ (_17479_, _17478_, _17477_);
  and _40293_ (_17480_, _17479_, _05997_);
  or _40294_ (_17481_, _17480_, _17476_);
  or _40295_ (_17482_, _17481_, _05920_);
  and _40296_ (_17483_, _17482_, _06033_);
  and _40297_ (_17484_, _17483_, _17472_);
  or _40298_ (_17485_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or _40299_ (_17486_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _40300_ (_17487_, _17486_, _05997_);
  and _40301_ (_17488_, _17487_, _17485_);
  or _40302_ (_17489_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _40303_ (_17490_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _40304_ (_17491_, _17490_, _05996_);
  and _40305_ (_17492_, _17491_, _17489_);
  or _40306_ (_17493_, _17492_, _17488_);
  or _40307_ (_17494_, _17493_, _06021_);
  or _40308_ (_17495_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or _40309_ (_17496_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and _40310_ (_17497_, _17496_, _05997_);
  and _40311_ (_17498_, _17497_, _17495_);
  or _40312_ (_17499_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _40313_ (_17500_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _40314_ (_17501_, _17500_, _05996_);
  and _40315_ (_17502_, _17501_, _17499_);
  or _40316_ (_17503_, _17502_, _17498_);
  or _40317_ (_17504_, _17503_, _05920_);
  and _40318_ (_17505_, _17504_, _05933_);
  and _40319_ (_17506_, _17505_, _17494_);
  or _40320_ (_17507_, _17506_, _17484_);
  and _40321_ (_17508_, _17507_, _06071_);
  or _40322_ (_17509_, _17508_, _17462_);
  and _40323_ (_17510_, _17509_, _06070_);
  and _40324_ (_17511_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and _40325_ (_17512_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or _40326_ (_17513_, _17512_, _17511_);
  and _40327_ (_17514_, _17513_, _05996_);
  and _40328_ (_17515_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _40329_ (_17516_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or _40330_ (_17517_, _17516_, _17515_);
  and _40331_ (_17518_, _17517_, _05997_);
  or _40332_ (_17519_, _17518_, _17514_);
  and _40333_ (_17520_, _17519_, _05920_);
  and _40334_ (_17521_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and _40335_ (_17522_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or _40336_ (_17523_, _17522_, _17521_);
  and _40337_ (_17524_, _17523_, _05996_);
  and _40338_ (_17525_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and _40339_ (_17526_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or _40340_ (_17527_, _17526_, _17525_);
  and _40341_ (_17528_, _17527_, _05997_);
  or _40342_ (_17529_, _17528_, _17524_);
  and _40343_ (_17530_, _17529_, _06021_);
  or _40344_ (_17531_, _17530_, _17520_);
  and _40345_ (_17532_, _17531_, _06033_);
  or _40346_ (_17533_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or _40347_ (_17534_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and _40348_ (_17535_, _17534_, _05997_);
  and _40349_ (_17536_, _17535_, _17533_);
  or _40350_ (_17537_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or _40351_ (_17538_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and _40352_ (_17539_, _17538_, _05996_);
  and _40353_ (_17540_, _17539_, _17537_);
  or _40354_ (_17541_, _17540_, _17536_);
  and _40355_ (_17542_, _17541_, _05920_);
  or _40356_ (_17543_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or _40357_ (_17544_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and _40358_ (_17545_, _17544_, _05997_);
  and _40359_ (_17546_, _17545_, _17543_);
  or _40360_ (_17547_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or _40361_ (_17548_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and _40362_ (_17549_, _17548_, _05996_);
  and _40363_ (_17550_, _17549_, _17547_);
  or _40364_ (_17551_, _17550_, _17546_);
  and _40365_ (_17552_, _17551_, _06021_);
  or _40366_ (_17553_, _17552_, _17542_);
  and _40367_ (_17554_, _17553_, _05933_);
  or _40368_ (_17555_, _17554_, _17532_);
  and _40369_ (_17556_, _17555_, _06071_);
  and _40370_ (_17557_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _40371_ (_17558_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _40372_ (_17559_, _17558_, _17557_);
  and _40373_ (_17560_, _17559_, _05996_);
  and _40374_ (_17561_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and _40375_ (_17562_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _40376_ (_17563_, _17562_, _17561_);
  and _40377_ (_17564_, _17563_, _05997_);
  or _40378_ (_17565_, _17564_, _17560_);
  and _40379_ (_17566_, _17565_, _05920_);
  and _40380_ (_17567_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and _40381_ (_17568_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _40382_ (_17569_, _17568_, _17567_);
  and _40383_ (_17570_, _17569_, _05996_);
  and _40384_ (_17571_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and _40385_ (_17572_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _40386_ (_17573_, _17572_, _17571_);
  and _40387_ (_17574_, _17573_, _05997_);
  or _40388_ (_17575_, _17574_, _17570_);
  and _40389_ (_17576_, _17575_, _06021_);
  or _40390_ (_17577_, _17576_, _17566_);
  and _40391_ (_17578_, _17577_, _06033_);
  or _40392_ (_17579_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _40393_ (_17580_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and _40394_ (_17581_, _17580_, _17579_);
  and _40395_ (_17582_, _17581_, _05996_);
  or _40396_ (_17583_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _40397_ (_17584_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and _40398_ (_17585_, _17584_, _17583_);
  and _40399_ (_17586_, _17585_, _05997_);
  or _40400_ (_17587_, _17586_, _17582_);
  and _40401_ (_17588_, _17587_, _05920_);
  or _40402_ (_17589_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _40403_ (_17590_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _40404_ (_17591_, _17590_, _17589_);
  and _40405_ (_17592_, _17591_, _05996_);
  or _40406_ (_17593_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _40407_ (_17594_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and _40408_ (_17595_, _17594_, _17593_);
  and _40409_ (_17596_, _17595_, _05997_);
  or _40410_ (_17597_, _17596_, _17592_);
  and _40411_ (_17598_, _17597_, _06021_);
  or _40412_ (_17599_, _17598_, _17588_);
  and _40413_ (_17601_, _17599_, _05933_);
  or _40414_ (_17602_, _17601_, _17578_);
  and _40415_ (_17603_, _17602_, _05776_);
  or _40416_ (_17604_, _17603_, _17556_);
  and _40417_ (_17605_, _17604_, _05822_);
  or _40418_ (_17606_, _17605_, _17510_);
  or _40419_ (_17607_, _17606_, _05868_);
  and _40420_ (_17608_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and _40421_ (_17609_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _40422_ (_17610_, _17609_, _17608_);
  and _40423_ (_17611_, _17610_, _05996_);
  and _40424_ (_17612_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and _40425_ (_17613_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _40426_ (_17614_, _17613_, _17612_);
  and _40427_ (_17615_, _17614_, _05997_);
  or _40428_ (_17616_, _17615_, _17611_);
  or _40429_ (_17617_, _17616_, _06021_);
  and _40430_ (_17618_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and _40431_ (_17619_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _40432_ (_17620_, _17619_, _17618_);
  and _40433_ (_17621_, _17620_, _05996_);
  and _40434_ (_17622_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and _40435_ (_17623_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _40436_ (_17624_, _17623_, _17622_);
  and _40437_ (_17625_, _17624_, _05997_);
  or _40438_ (_17626_, _17625_, _17621_);
  or _40439_ (_17627_, _17626_, _05920_);
  and _40440_ (_17628_, _17627_, _06033_);
  and _40441_ (_17629_, _17628_, _17617_);
  or _40442_ (_17630_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _40443_ (_17631_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and _40444_ (_17632_, _17631_, _05997_);
  and _40445_ (_17633_, _17632_, _17630_);
  or _40446_ (_17634_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _40447_ (_17635_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and _40448_ (_17636_, _17635_, _05996_);
  and _40449_ (_17637_, _17636_, _17634_);
  or _40450_ (_17638_, _17637_, _17633_);
  or _40451_ (_17639_, _17638_, _06021_);
  or _40452_ (_17640_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _40453_ (_17641_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and _40454_ (_17642_, _17641_, _05997_);
  and _40455_ (_17643_, _17642_, _17640_);
  or _40456_ (_17644_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _40457_ (_17645_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and _40458_ (_17646_, _17645_, _05996_);
  and _40459_ (_17647_, _17646_, _17644_);
  or _40460_ (_17648_, _17647_, _17643_);
  or _40461_ (_17649_, _17648_, _05920_);
  and _40462_ (_17650_, _17649_, _05933_);
  and _40463_ (_17651_, _17650_, _17639_);
  or _40464_ (_17652_, _17651_, _17629_);
  and _40465_ (_17653_, _17652_, _06071_);
  and _40466_ (_17654_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and _40467_ (_17655_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or _40468_ (_17656_, _17655_, _17654_);
  and _40469_ (_17657_, _17656_, _05996_);
  and _40470_ (_17658_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _40471_ (_17659_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _40472_ (_17660_, _17659_, _17658_);
  and _40473_ (_17661_, _17660_, _05997_);
  or _40474_ (_17662_, _17661_, _17657_);
  or _40475_ (_17663_, _17662_, _06021_);
  and _40476_ (_17664_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _40477_ (_17665_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or _40478_ (_17666_, _17665_, _17664_);
  and _40479_ (_17667_, _17666_, _05996_);
  and _40480_ (_17668_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _40481_ (_17669_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _40482_ (_17670_, _17669_, _17668_);
  and _40483_ (_17671_, _17670_, _05997_);
  or _40484_ (_17672_, _17671_, _17667_);
  or _40485_ (_17673_, _17672_, _05920_);
  and _40486_ (_17674_, _17673_, _06033_);
  and _40487_ (_17675_, _17674_, _17663_);
  or _40488_ (_17676_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _40489_ (_17677_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _40490_ (_17678_, _17677_, _17676_);
  and _40491_ (_17679_, _17678_, _05996_);
  or _40492_ (_17680_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _40493_ (_17681_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and _40494_ (_17682_, _17681_, _17680_);
  and _40495_ (_17683_, _17682_, _05997_);
  or _40496_ (_17684_, _17683_, _17679_);
  or _40497_ (_17685_, _17684_, _06021_);
  or _40498_ (_17686_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or _40499_ (_17687_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _40500_ (_17688_, _17687_, _17686_);
  and _40501_ (_17689_, _17688_, _05996_);
  or _40502_ (_17690_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _40503_ (_17691_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _40504_ (_17692_, _17691_, _17690_);
  and _40505_ (_17693_, _17692_, _05997_);
  or _40506_ (_17694_, _17693_, _17689_);
  or _40507_ (_17695_, _17694_, _05920_);
  and _40508_ (_17696_, _17695_, _05933_);
  and _40509_ (_17697_, _17696_, _17685_);
  or _40510_ (_17698_, _17697_, _17675_);
  and _40511_ (_17699_, _17698_, _05776_);
  or _40512_ (_17700_, _17699_, _17653_);
  and _40513_ (_17701_, _17700_, _06070_);
  or _40514_ (_17702_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _40515_ (_17703_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and _40516_ (_17704_, _17703_, _17702_);
  and _40517_ (_17705_, _17704_, _05996_);
  or _40518_ (_17706_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _40519_ (_17707_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _40520_ (_17708_, _17707_, _17706_);
  and _40521_ (_17709_, _17708_, _05997_);
  or _40522_ (_17710_, _17709_, _17705_);
  and _40523_ (_17711_, _17710_, _06021_);
  or _40524_ (_17712_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _40525_ (_17713_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _40526_ (_17714_, _17713_, _17712_);
  and _40527_ (_17715_, _17714_, _05996_);
  or _40528_ (_17716_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or _40529_ (_17717_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _40530_ (_17718_, _17717_, _17716_);
  and _40531_ (_17719_, _17718_, _05997_);
  or _40532_ (_17720_, _17719_, _17715_);
  and _40533_ (_17721_, _17720_, _05920_);
  or _40534_ (_17722_, _17721_, _17711_);
  and _40535_ (_17723_, _17722_, _05933_);
  and _40536_ (_17724_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _40537_ (_17725_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or _40538_ (_17726_, _17725_, _17724_);
  and _40539_ (_17727_, _17726_, _05996_);
  and _40540_ (_17728_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _40541_ (_17729_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _40542_ (_17730_, _17729_, _17728_);
  and _40543_ (_17731_, _17730_, _05997_);
  or _40544_ (_17732_, _17731_, _17727_);
  and _40545_ (_17733_, _17732_, _06021_);
  and _40546_ (_17734_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _40547_ (_17735_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _40548_ (_17736_, _17735_, _17734_);
  and _40549_ (_17737_, _17736_, _05996_);
  and _40550_ (_17738_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _40551_ (_17739_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or _40552_ (_17740_, _17739_, _17738_);
  and _40553_ (_17741_, _17740_, _05997_);
  or _40554_ (_17742_, _17741_, _17737_);
  and _40555_ (_17743_, _17742_, _05920_);
  or _40556_ (_17744_, _17743_, _17733_);
  and _40557_ (_17745_, _17744_, _06033_);
  or _40558_ (_17746_, _17745_, _17723_);
  and _40559_ (_17747_, _17746_, _05776_);
  or _40560_ (_17748_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _40561_ (_17749_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and _40562_ (_17750_, _17749_, _05997_);
  and _40563_ (_17751_, _17750_, _17748_);
  or _40564_ (_17752_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _40565_ (_17753_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and _40566_ (_17754_, _17753_, _05996_);
  and _40567_ (_17755_, _17754_, _17752_);
  or _40568_ (_17756_, _17755_, _17751_);
  and _40569_ (_17757_, _17756_, _06021_);
  or _40570_ (_17758_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _40571_ (_17759_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and _40572_ (_17760_, _17759_, _05997_);
  and _40573_ (_17761_, _17760_, _17758_);
  or _40574_ (_17762_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _40575_ (_17763_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and _40576_ (_17764_, _17763_, _05996_);
  and _40577_ (_17765_, _17764_, _17762_);
  or _40578_ (_17766_, _17765_, _17761_);
  and _40579_ (_17767_, _17766_, _05920_);
  or _40580_ (_17768_, _17767_, _17757_);
  and _40581_ (_17769_, _17768_, _05933_);
  and _40582_ (_17770_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and _40583_ (_17771_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _40584_ (_17772_, _17771_, _17770_);
  and _40585_ (_17773_, _17772_, _05996_);
  and _40586_ (_17774_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and _40587_ (_17775_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _40588_ (_17776_, _17775_, _17774_);
  and _40589_ (_17777_, _17776_, _05997_);
  or _40590_ (_17778_, _17777_, _17773_);
  and _40591_ (_17779_, _17778_, _06021_);
  and _40592_ (_17780_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and _40593_ (_17781_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _40594_ (_17782_, _17781_, _17780_);
  and _40595_ (_17783_, _17782_, _05996_);
  and _40596_ (_17784_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _40597_ (_17785_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _40598_ (_17786_, _17785_, _17784_);
  and _40599_ (_17787_, _17786_, _05997_);
  or _40600_ (_17788_, _17787_, _17783_);
  and _40601_ (_17789_, _17788_, _05920_);
  or _40602_ (_17790_, _17789_, _17779_);
  and _40603_ (_17791_, _17790_, _06033_);
  or _40604_ (_17792_, _17791_, _17769_);
  and _40605_ (_17793_, _17792_, _06071_);
  or _40606_ (_17794_, _17793_, _17747_);
  and _40607_ (_17795_, _17794_, _05822_);
  or _40608_ (_17796_, _17795_, _17701_);
  or _40609_ (_17797_, _17796_, _06616_);
  and _40610_ (_17798_, _17797_, _17607_);
  or _40611_ (_17799_, _17798_, _05584_);
  and _40612_ (_17800_, _17799_, _17416_);
  or _40613_ (_17801_, _17800_, _06019_);
  or _40614_ (_17802_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _40615_ (_17803_, _17802_, _25365_);
  and _40616_ (_14804_, _17803_, _17801_);
  and _40617_ (_17804_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and _40618_ (_17805_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _40619_ (_17806_, _17805_, _17804_);
  and _40620_ (_17807_, _17806_, _05996_);
  and _40621_ (_17808_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and _40622_ (_17809_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _40623_ (_17810_, _17809_, _17808_);
  and _40624_ (_17811_, _17810_, _05997_);
  or _40625_ (_17812_, _17811_, _17807_);
  or _40626_ (_17813_, _17812_, _06021_);
  and _40627_ (_17814_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and _40628_ (_17815_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _40629_ (_17816_, _17815_, _17814_);
  and _40630_ (_17817_, _17816_, _05996_);
  and _40631_ (_17818_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and _40632_ (_17819_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _40633_ (_17820_, _17819_, _17818_);
  and _40634_ (_17821_, _17820_, _05997_);
  or _40635_ (_17822_, _17821_, _17817_);
  or _40636_ (_17823_, _17822_, _05920_);
  and _40637_ (_17824_, _17823_, _06033_);
  and _40638_ (_17825_, _17824_, _17813_);
  or _40639_ (_17826_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _40640_ (_17827_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and _40641_ (_17828_, _17827_, _17826_);
  and _40642_ (_17829_, _17828_, _05996_);
  or _40643_ (_17830_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _40644_ (_17831_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and _40645_ (_17832_, _17831_, _17830_);
  and _40646_ (_17833_, _17832_, _05997_);
  or _40647_ (_17834_, _17833_, _17829_);
  or _40648_ (_17835_, _17834_, _06021_);
  or _40649_ (_17836_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _40650_ (_17837_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and _40651_ (_17838_, _17837_, _17836_);
  and _40652_ (_17839_, _17838_, _05996_);
  or _40653_ (_17840_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _40654_ (_17841_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and _40655_ (_17842_, _17841_, _17840_);
  and _40656_ (_17843_, _17842_, _05997_);
  or _40657_ (_17844_, _17843_, _17839_);
  or _40658_ (_17845_, _17844_, _05920_);
  and _40659_ (_17846_, _17845_, _05933_);
  and _40660_ (_17847_, _17846_, _17835_);
  or _40661_ (_17848_, _17847_, _17825_);
  or _40662_ (_17849_, _17848_, _06071_);
  and _40663_ (_17850_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and _40664_ (_17851_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _40665_ (_17852_, _17851_, _17850_);
  and _40666_ (_17853_, _17852_, _05996_);
  and _40667_ (_17854_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and _40668_ (_17855_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _40669_ (_17856_, _17855_, _17854_);
  and _40670_ (_17857_, _17856_, _05997_);
  or _40671_ (_17858_, _17857_, _17853_);
  or _40672_ (_17859_, _17858_, _06021_);
  and _40673_ (_17860_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and _40674_ (_17861_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _40675_ (_17862_, _17861_, _17860_);
  and _40676_ (_17863_, _17862_, _05996_);
  and _40677_ (_17864_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and _40678_ (_17865_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _40679_ (_17866_, _17865_, _17864_);
  and _40680_ (_17867_, _17866_, _05997_);
  or _40681_ (_17868_, _17867_, _17863_);
  or _40682_ (_17869_, _17868_, _05920_);
  and _40683_ (_17870_, _17869_, _06033_);
  and _40684_ (_17871_, _17870_, _17859_);
  or _40685_ (_17872_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _40686_ (_17873_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and _40687_ (_17874_, _17873_, _05997_);
  and _40688_ (_17875_, _17874_, _17872_);
  or _40689_ (_17876_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _40690_ (_17877_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and _40691_ (_17878_, _17877_, _05996_);
  and _40692_ (_17879_, _17878_, _17876_);
  or _40693_ (_17880_, _17879_, _17875_);
  or _40694_ (_17881_, _17880_, _06021_);
  or _40695_ (_17882_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _40696_ (_17883_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and _40697_ (_17884_, _17883_, _05997_);
  and _40698_ (_17885_, _17884_, _17882_);
  or _40699_ (_17886_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _40700_ (_17887_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and _40701_ (_17888_, _17887_, _05996_);
  and _40702_ (_17889_, _17888_, _17886_);
  or _40703_ (_17890_, _17889_, _17885_);
  or _40704_ (_17891_, _17890_, _05920_);
  and _40705_ (_17892_, _17891_, _05933_);
  and _40706_ (_17893_, _17892_, _17881_);
  or _40707_ (_17894_, _17893_, _17871_);
  or _40708_ (_17895_, _17894_, _05776_);
  and _40709_ (_17896_, _17895_, _06070_);
  and _40710_ (_17897_, _17896_, _17849_);
  and _40711_ (_17898_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _40712_ (_17899_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or _40713_ (_17900_, _17899_, _17898_);
  and _40714_ (_17901_, _17900_, _05996_);
  and _40715_ (_17902_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _40716_ (_17903_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _40717_ (_17904_, _17903_, _17902_);
  and _40718_ (_17905_, _17904_, _05997_);
  or _40719_ (_17906_, _17905_, _17901_);
  and _40720_ (_17907_, _17906_, _05920_);
  and _40721_ (_17908_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _40722_ (_17909_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _40723_ (_17910_, _17909_, _17908_);
  and _40724_ (_17911_, _17910_, _05996_);
  and _40725_ (_17912_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and _40726_ (_17913_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _40727_ (_17914_, _17913_, _17912_);
  and _40728_ (_17915_, _17914_, _05997_);
  or _40729_ (_17916_, _17915_, _17911_);
  and _40730_ (_17917_, _17916_, _06021_);
  or _40731_ (_17918_, _17917_, _05933_);
  or _40732_ (_17919_, _17918_, _17907_);
  or _40733_ (_17920_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _40734_ (_17921_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and _40735_ (_17922_, _17921_, _05997_);
  and _40736_ (_17923_, _17922_, _17920_);
  or _40737_ (_17924_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _40738_ (_17925_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _40739_ (_17926_, _17925_, _05996_);
  and _40740_ (_17927_, _17926_, _17924_);
  or _40741_ (_17928_, _17927_, _17923_);
  and _40742_ (_17929_, _17928_, _05920_);
  or _40743_ (_17930_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _40744_ (_17931_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _40745_ (_17932_, _17931_, _05997_);
  and _40746_ (_17933_, _17932_, _17930_);
  or _40747_ (_17934_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _40748_ (_17935_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _40749_ (_17936_, _17935_, _05996_);
  and _40750_ (_17937_, _17936_, _17934_);
  or _40751_ (_17938_, _17937_, _17933_);
  and _40752_ (_17939_, _17938_, _06021_);
  or _40753_ (_17940_, _17939_, _06033_);
  or _40754_ (_17941_, _17940_, _17929_);
  and _40755_ (_17942_, _17941_, _17919_);
  or _40756_ (_17943_, _17942_, _05776_);
  and _40757_ (_17944_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and _40758_ (_17945_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _40759_ (_17946_, _17945_, _17944_);
  and _40760_ (_17947_, _17946_, _05996_);
  and _40761_ (_17948_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and _40762_ (_17949_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _40763_ (_17950_, _17949_, _17948_);
  and _40764_ (_17951_, _17950_, _05997_);
  or _40765_ (_17952_, _17951_, _17947_);
  and _40766_ (_17953_, _17952_, _05920_);
  and _40767_ (_17954_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and _40768_ (_17955_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _40769_ (_17956_, _17955_, _17954_);
  and _40770_ (_17957_, _17956_, _05996_);
  and _40771_ (_17958_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and _40772_ (_17959_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _40773_ (_17960_, _17959_, _17958_);
  and _40774_ (_17961_, _17960_, _05997_);
  or _40775_ (_17962_, _17961_, _17957_);
  and _40776_ (_17963_, _17962_, _06021_);
  or _40777_ (_17964_, _17963_, _05933_);
  or _40778_ (_17965_, _17964_, _17953_);
  or _40779_ (_17966_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _40780_ (_17967_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and _40781_ (_17968_, _17967_, _17966_);
  and _40782_ (_17969_, _17968_, _05996_);
  or _40783_ (_17970_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _40784_ (_17971_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and _40785_ (_17972_, _17971_, _17970_);
  and _40786_ (_17973_, _17972_, _05997_);
  or _40787_ (_17974_, _17973_, _17969_);
  and _40788_ (_17975_, _17974_, _05920_);
  or _40789_ (_17976_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _40790_ (_17977_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and _40791_ (_17978_, _17977_, _17976_);
  and _40792_ (_17979_, _17978_, _05996_);
  or _40793_ (_17980_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _40794_ (_17981_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and _40795_ (_17982_, _17981_, _17980_);
  and _40796_ (_17983_, _17982_, _05997_);
  or _40797_ (_17984_, _17983_, _17979_);
  and _40798_ (_17985_, _17984_, _06021_);
  or _40799_ (_17986_, _17985_, _06033_);
  or _40800_ (_17987_, _17986_, _17975_);
  and _40801_ (_17988_, _17987_, _17965_);
  or _40802_ (_17989_, _17988_, _06071_);
  and _40803_ (_17990_, _17989_, _05822_);
  and _40804_ (_17991_, _17990_, _17943_);
  or _40805_ (_17992_, _17991_, _17897_);
  or _40806_ (_17993_, _17992_, _05868_);
  and _40807_ (_17994_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and _40808_ (_17995_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or _40809_ (_17996_, _17995_, _17994_);
  and _40810_ (_17997_, _17996_, _05996_);
  and _40811_ (_17998_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and _40812_ (_17999_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or _40813_ (_18000_, _17999_, _17998_);
  and _40814_ (_18001_, _18000_, _05997_);
  or _40815_ (_18002_, _18001_, _17997_);
  and _40816_ (_18003_, _18002_, _05920_);
  and _40817_ (_18004_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and _40818_ (_18005_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or _40819_ (_18006_, _18005_, _18004_);
  and _40820_ (_18007_, _18006_, _05996_);
  and _40821_ (_18008_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  and _40822_ (_18009_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or _40823_ (_18010_, _18009_, _18008_);
  and _40824_ (_18011_, _18010_, _05997_);
  or _40825_ (_18012_, _18011_, _18007_);
  and _40826_ (_18013_, _18012_, _06021_);
  or _40827_ (_18014_, _18013_, _05933_);
  or _40828_ (_18015_, _18014_, _18003_);
  or _40829_ (_18016_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or _40830_ (_18017_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and _40831_ (_18018_, _18017_, _18016_);
  and _40832_ (_18019_, _18018_, _05996_);
  or _40833_ (_18020_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or _40834_ (_18021_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  and _40835_ (_18022_, _18021_, _18020_);
  and _40836_ (_18023_, _18022_, _05997_);
  or _40837_ (_18024_, _18023_, _18019_);
  and _40838_ (_18025_, _18024_, _05920_);
  or _40839_ (_18026_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or _40840_ (_18027_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and _40841_ (_18028_, _18027_, _18026_);
  and _40842_ (_18029_, _18028_, _05996_);
  or _40843_ (_18030_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or _40844_ (_18031_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and _40845_ (_18032_, _18031_, _18030_);
  and _40846_ (_18033_, _18032_, _05997_);
  or _40847_ (_18034_, _18033_, _18029_);
  and _40848_ (_18035_, _18034_, _06021_);
  or _40849_ (_18036_, _18035_, _06033_);
  or _40850_ (_18037_, _18036_, _18025_);
  and _40851_ (_18038_, _18037_, _18015_);
  or _40852_ (_18039_, _18038_, _05776_);
  and _40853_ (_18040_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and _40854_ (_18041_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _40855_ (_18042_, _18041_, _18040_);
  and _40856_ (_18043_, _18042_, _05996_);
  and _40857_ (_18044_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and _40858_ (_18045_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _40859_ (_18046_, _18045_, _18044_);
  and _40860_ (_18047_, _18046_, _05997_);
  or _40861_ (_18048_, _18047_, _18043_);
  and _40862_ (_18049_, _18048_, _05920_);
  and _40863_ (_18050_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and _40864_ (_18051_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _40865_ (_18052_, _18051_, _18050_);
  and _40866_ (_18053_, _18052_, _05996_);
  and _40867_ (_18054_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and _40868_ (_18055_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _40869_ (_18056_, _18055_, _18054_);
  and _40870_ (_18057_, _18056_, _05997_);
  or _40871_ (_18058_, _18057_, _18053_);
  and _40872_ (_18059_, _18058_, _06021_);
  or _40873_ (_18060_, _18059_, _05933_);
  or _40874_ (_18061_, _18060_, _18049_);
  or _40875_ (_18062_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _40876_ (_18063_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and _40877_ (_18064_, _18063_, _18062_);
  and _40878_ (_18065_, _18064_, _05996_);
  or _40879_ (_18066_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _40880_ (_18067_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and _40881_ (_18068_, _18067_, _18066_);
  and _40882_ (_18069_, _18068_, _05997_);
  or _40883_ (_18070_, _18069_, _18065_);
  and _40884_ (_18071_, _18070_, _05920_);
  or _40885_ (_18072_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _40886_ (_18073_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and _40887_ (_18074_, _18073_, _18072_);
  and _40888_ (_18075_, _18074_, _05996_);
  or _40889_ (_18076_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _40890_ (_18077_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and _40891_ (_18078_, _18077_, _18076_);
  and _40892_ (_18079_, _18078_, _05997_);
  or _40893_ (_18080_, _18079_, _18075_);
  and _40894_ (_18081_, _18080_, _06021_);
  or _40895_ (_18082_, _18081_, _06033_);
  or _40896_ (_18083_, _18082_, _18071_);
  and _40897_ (_18084_, _18083_, _18061_);
  or _40898_ (_18085_, _18084_, _06071_);
  and _40899_ (_18086_, _18085_, _05822_);
  and _40900_ (_18087_, _18086_, _18039_);
  and _40901_ (_18088_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and _40902_ (_18089_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _40903_ (_18090_, _18089_, _18088_);
  and _40904_ (_18091_, _18090_, _05997_);
  and _40905_ (_18092_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and _40906_ (_18093_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _40907_ (_18094_, _18093_, _18092_);
  and _40908_ (_18095_, _18094_, _05996_);
  or _40909_ (_18096_, _18095_, _18091_);
  or _40910_ (_18097_, _18096_, _06021_);
  and _40911_ (_18098_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and _40912_ (_18099_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _40913_ (_18100_, _18099_, _18098_);
  and _40914_ (_18101_, _18100_, _05997_);
  and _40915_ (_18102_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and _40916_ (_18103_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _40917_ (_18104_, _18103_, _18102_);
  and _40918_ (_18105_, _18104_, _05996_);
  or _40919_ (_18106_, _18105_, _18101_);
  or _40920_ (_18107_, _18106_, _05920_);
  and _40921_ (_18108_, _18107_, _06033_);
  and _40922_ (_18109_, _18108_, _18097_);
  or _40923_ (_18110_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _40924_ (_18111_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and _40925_ (_18112_, _18111_, _05996_);
  and _40926_ (_18113_, _18112_, _18110_);
  or _40927_ (_18114_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _40928_ (_18115_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and _40929_ (_18116_, _18115_, _05997_);
  and _40930_ (_18117_, _18116_, _18114_);
  or _40931_ (_18118_, _18117_, _18113_);
  or _40932_ (_18119_, _18118_, _06021_);
  or _40933_ (_18120_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _40934_ (_18121_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and _40935_ (_18122_, _18121_, _05996_);
  and _40936_ (_18123_, _18122_, _18120_);
  or _40937_ (_18124_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _40938_ (_18125_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and _40939_ (_18126_, _18125_, _05997_);
  and _40940_ (_18127_, _18126_, _18124_);
  or _40941_ (_18128_, _18127_, _18123_);
  or _40942_ (_18129_, _18128_, _05920_);
  and _40943_ (_18130_, _18129_, _05933_);
  and _40944_ (_18131_, _18130_, _18119_);
  or _40945_ (_18132_, _18131_, _18109_);
  and _40946_ (_18133_, _18132_, _06071_);
  and _40947_ (_18134_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _40948_ (_18135_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _40949_ (_18136_, _18135_, _05996_);
  or _40950_ (_18137_, _18136_, _18134_);
  and _40951_ (_18138_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and _40952_ (_18139_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _40953_ (_18140_, _18139_, _05997_);
  or _40954_ (_18141_, _18140_, _18138_);
  and _40955_ (_18142_, _18141_, _18137_);
  or _40956_ (_18143_, _18142_, _06021_);
  and _40957_ (_18144_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and _40958_ (_18145_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _40959_ (_18146_, _18145_, _05996_);
  or _40960_ (_18147_, _18146_, _18144_);
  and _40961_ (_18148_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and _40962_ (_18149_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _40963_ (_18150_, _18149_, _05997_);
  or _40964_ (_18151_, _18150_, _18148_);
  and _40965_ (_18152_, _18151_, _18147_);
  or _40966_ (_18153_, _18152_, _05920_);
  and _40967_ (_18154_, _18153_, _06033_);
  and _40968_ (_18155_, _18154_, _18143_);
  or _40969_ (_18156_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _40970_ (_18157_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and _40971_ (_18158_, _18157_, _18156_);
  or _40972_ (_18159_, _18158_, _05997_);
  or _40973_ (_18160_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _40974_ (_18161_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _40975_ (_18162_, _18161_, _18160_);
  or _40976_ (_18163_, _18162_, _05996_);
  and _40977_ (_18164_, _18163_, _18159_);
  or _40978_ (_18165_, _18164_, _06021_);
  or _40979_ (_18166_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _40980_ (_18167_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and _40981_ (_18168_, _18167_, _18166_);
  or _40982_ (_18169_, _18168_, _05997_);
  or _40983_ (_18170_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _40984_ (_18171_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _40985_ (_18172_, _18171_, _18170_);
  or _40986_ (_18173_, _18172_, _05996_);
  and _40987_ (_18174_, _18173_, _18169_);
  or _40988_ (_18175_, _18174_, _05920_);
  and _40989_ (_18176_, _18175_, _05933_);
  and _40990_ (_18177_, _18176_, _18165_);
  or _40991_ (_18178_, _18177_, _18155_);
  and _40992_ (_18179_, _18178_, _05776_);
  or _40993_ (_18180_, _18179_, _18133_);
  and _40994_ (_18181_, _18180_, _06070_);
  or _40995_ (_18182_, _18181_, _18087_);
  or _40996_ (_18183_, _18182_, _06616_);
  and _40997_ (_18184_, _18183_, _17993_);
  or _40998_ (_18185_, _18184_, _06020_);
  and _40999_ (_18186_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and _41000_ (_18187_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _41001_ (_18188_, _18187_, _18186_);
  and _41002_ (_18189_, _18188_, _05996_);
  and _41003_ (_18190_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and _41004_ (_18191_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _41005_ (_18192_, _18191_, _18190_);
  and _41006_ (_18193_, _18192_, _05997_);
  or _41007_ (_18194_, _18193_, _18189_);
  or _41008_ (_18195_, _18194_, _06021_);
  and _41009_ (_18196_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and _41010_ (_18197_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _41011_ (_18198_, _18197_, _18196_);
  and _41012_ (_18199_, _18198_, _05996_);
  and _41013_ (_18200_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and _41014_ (_18201_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _41015_ (_18202_, _18201_, _18200_);
  and _41016_ (_18203_, _18202_, _05997_);
  or _41017_ (_18204_, _18203_, _18199_);
  or _41018_ (_18205_, _18204_, _05920_);
  and _41019_ (_18206_, _18205_, _06033_);
  and _41020_ (_18207_, _18206_, _18195_);
  or _41021_ (_18208_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _41022_ (_18209_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and _41023_ (_18210_, _18209_, _18208_);
  and _41024_ (_18211_, _18210_, _05996_);
  or _41025_ (_18212_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _41026_ (_18213_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and _41027_ (_18214_, _18213_, _18212_);
  and _41028_ (_18215_, _18214_, _05997_);
  or _41029_ (_18216_, _18215_, _18211_);
  or _41030_ (_18217_, _18216_, _06021_);
  or _41031_ (_18218_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _41032_ (_18219_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and _41033_ (_18220_, _18219_, _18218_);
  and _41034_ (_18221_, _18220_, _05996_);
  or _41035_ (_18222_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _41036_ (_18223_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and _41037_ (_18224_, _18223_, _18222_);
  and _41038_ (_18225_, _18224_, _05997_);
  or _41039_ (_18226_, _18225_, _18221_);
  or _41040_ (_18227_, _18226_, _05920_);
  and _41041_ (_18228_, _18227_, _05933_);
  and _41042_ (_18229_, _18228_, _18217_);
  or _41043_ (_18230_, _18229_, _18207_);
  and _41044_ (_18231_, _18230_, _05776_);
  and _41045_ (_18232_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and _41046_ (_18233_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _41047_ (_18234_, _18233_, _18232_);
  and _41048_ (_18235_, _18234_, _05996_);
  and _41049_ (_18236_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _41050_ (_18237_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _41051_ (_18238_, _18237_, _18236_);
  and _41052_ (_18239_, _18238_, _05997_);
  or _41053_ (_18240_, _18239_, _18235_);
  or _41054_ (_18241_, _18240_, _06021_);
  and _41055_ (_18242_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and _41056_ (_18243_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or _41057_ (_18244_, _18243_, _18242_);
  and _41058_ (_18245_, _18244_, _05996_);
  and _41059_ (_18246_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _41060_ (_18247_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _41061_ (_18248_, _18247_, _18246_);
  and _41062_ (_18249_, _18248_, _05997_);
  or _41063_ (_18250_, _18249_, _18245_);
  or _41064_ (_18251_, _18250_, _05920_);
  and _41065_ (_18252_, _18251_, _06033_);
  and _41066_ (_18253_, _18252_, _18241_);
  or _41067_ (_18254_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or _41068_ (_18255_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _41069_ (_18256_, _18255_, _05997_);
  and _41070_ (_18257_, _18256_, _18254_);
  or _41071_ (_18258_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _41072_ (_18259_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _41073_ (_18260_, _18259_, _05996_);
  and _41074_ (_18261_, _18260_, _18258_);
  or _41075_ (_18262_, _18261_, _18257_);
  or _41076_ (_18263_, _18262_, _06021_);
  or _41077_ (_18264_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _41078_ (_18265_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _41079_ (_18266_, _18265_, _05997_);
  and _41080_ (_18267_, _18266_, _18264_);
  or _41081_ (_18268_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or _41082_ (_18269_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and _41083_ (_18270_, _18269_, _05996_);
  and _41084_ (_18271_, _18270_, _18268_);
  or _41085_ (_18272_, _18271_, _18267_);
  or _41086_ (_18273_, _18272_, _05920_);
  and _41087_ (_18274_, _18273_, _05933_);
  and _41088_ (_18275_, _18274_, _18263_);
  or _41089_ (_18276_, _18275_, _18253_);
  and _41090_ (_18277_, _18276_, _06071_);
  or _41091_ (_18278_, _18277_, _18231_);
  and _41092_ (_18279_, _18278_, _06070_);
  and _41093_ (_18280_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and _41094_ (_18281_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or _41095_ (_18282_, _18281_, _18280_);
  and _41096_ (_18283_, _18282_, _05996_);
  and _41097_ (_18284_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and _41098_ (_18285_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or _41099_ (_18286_, _18285_, _18284_);
  and _41100_ (_18287_, _18286_, _05997_);
  or _41101_ (_18288_, _18287_, _18283_);
  and _41102_ (_18289_, _18288_, _05920_);
  and _41103_ (_18290_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and _41104_ (_18291_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or _41105_ (_18292_, _18291_, _18290_);
  and _41106_ (_18293_, _18292_, _05996_);
  and _41107_ (_18294_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _41108_ (_18295_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or _41109_ (_18296_, _18295_, _18294_);
  and _41110_ (_18297_, _18296_, _05997_);
  or _41111_ (_18298_, _18297_, _18293_);
  and _41112_ (_18299_, _18298_, _06021_);
  or _41113_ (_18300_, _18299_, _18289_);
  and _41114_ (_18301_, _18300_, _06033_);
  or _41115_ (_18302_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or _41116_ (_18303_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and _41117_ (_18304_, _18303_, _05997_);
  and _41118_ (_18305_, _18304_, _18302_);
  or _41119_ (_18306_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or _41120_ (_18307_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and _41121_ (_18308_, _18307_, _05996_);
  and _41122_ (_18309_, _18308_, _18306_);
  or _41123_ (_18310_, _18309_, _18305_);
  and _41124_ (_18311_, _18310_, _05920_);
  or _41125_ (_18312_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or _41126_ (_18313_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and _41127_ (_18314_, _18313_, _05997_);
  and _41128_ (_18315_, _18314_, _18312_);
  or _41129_ (_18316_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or _41130_ (_18317_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _41131_ (_18318_, _18317_, _05996_);
  and _41132_ (_18319_, _18318_, _18316_);
  or _41133_ (_18320_, _18319_, _18315_);
  and _41134_ (_18321_, _18320_, _06021_);
  or _41135_ (_18322_, _18321_, _18311_);
  and _41136_ (_18323_, _18322_, _05933_);
  or _41137_ (_18324_, _18323_, _18301_);
  and _41138_ (_18325_, _18324_, _06071_);
  and _41139_ (_18326_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _41140_ (_18327_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _41141_ (_18328_, _18327_, _18326_);
  and _41142_ (_18329_, _18328_, _05996_);
  and _41143_ (_18330_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _41144_ (_18331_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _41145_ (_18332_, _18331_, _18330_);
  and _41146_ (_18333_, _18332_, _05997_);
  or _41147_ (_18334_, _18333_, _18329_);
  and _41148_ (_18335_, _18334_, _05920_);
  and _41149_ (_18336_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and _41150_ (_18337_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _41151_ (_18338_, _18337_, _18336_);
  and _41152_ (_18339_, _18338_, _05996_);
  and _41153_ (_18340_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and _41154_ (_18341_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _41155_ (_18342_, _18341_, _18340_);
  and _41156_ (_18343_, _18342_, _05997_);
  or _41157_ (_18344_, _18343_, _18339_);
  and _41158_ (_18345_, _18344_, _06021_);
  or _41159_ (_18346_, _18345_, _18335_);
  and _41160_ (_18347_, _18346_, _06033_);
  or _41161_ (_18348_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _41162_ (_18349_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and _41163_ (_18350_, _18349_, _18348_);
  and _41164_ (_18351_, _18350_, _05996_);
  or _41165_ (_18352_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _41166_ (_18353_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and _41167_ (_18354_, _18353_, _18352_);
  and _41168_ (_18355_, _18354_, _05997_);
  or _41169_ (_18356_, _18355_, _18351_);
  and _41170_ (_18357_, _18356_, _05920_);
  or _41171_ (_18358_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _41172_ (_18359_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and _41173_ (_18360_, _18359_, _18358_);
  and _41174_ (_18361_, _18360_, _05996_);
  or _41175_ (_18362_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _41176_ (_18363_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _41177_ (_18364_, _18363_, _18362_);
  and _41178_ (_18365_, _18364_, _05997_);
  or _41179_ (_18366_, _18365_, _18361_);
  and _41180_ (_18367_, _18366_, _06021_);
  or _41181_ (_18368_, _18367_, _18357_);
  and _41182_ (_18369_, _18368_, _05933_);
  or _41183_ (_18370_, _18369_, _18347_);
  and _41184_ (_18371_, _18370_, _05776_);
  or _41185_ (_18372_, _18371_, _18325_);
  and _41186_ (_18373_, _18372_, _05822_);
  or _41187_ (_18374_, _18373_, _18279_);
  or _41188_ (_18375_, _18374_, _05868_);
  and _41189_ (_18376_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and _41190_ (_18377_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _41191_ (_18378_, _18377_, _18376_);
  and _41192_ (_18379_, _18378_, _05996_);
  and _41193_ (_18380_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and _41194_ (_18381_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _41195_ (_18382_, _18381_, _18380_);
  and _41196_ (_18383_, _18382_, _05997_);
  or _41197_ (_18384_, _18383_, _18379_);
  or _41198_ (_18385_, _18384_, _06021_);
  and _41199_ (_18386_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and _41200_ (_18387_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _41201_ (_18388_, _18387_, _18386_);
  and _41202_ (_18389_, _18388_, _05996_);
  and _41203_ (_18390_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and _41204_ (_18391_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _41205_ (_18392_, _18391_, _18390_);
  and _41206_ (_18393_, _18392_, _05997_);
  or _41207_ (_18394_, _18393_, _18389_);
  or _41208_ (_18395_, _18394_, _05920_);
  and _41209_ (_18396_, _18395_, _06033_);
  and _41210_ (_18397_, _18396_, _18385_);
  or _41211_ (_18398_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _41212_ (_18399_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and _41213_ (_18400_, _18399_, _05997_);
  and _41214_ (_18401_, _18400_, _18398_);
  or _41215_ (_18402_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _41216_ (_18403_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and _41217_ (_18404_, _18403_, _05996_);
  and _41218_ (_18405_, _18404_, _18402_);
  or _41219_ (_18406_, _18405_, _18401_);
  or _41220_ (_18407_, _18406_, _06021_);
  or _41221_ (_18408_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _41222_ (_18409_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and _41223_ (_18410_, _18409_, _05997_);
  and _41224_ (_18411_, _18410_, _18408_);
  or _41225_ (_18412_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _41226_ (_18413_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and _41227_ (_18414_, _18413_, _05996_);
  and _41228_ (_18415_, _18414_, _18412_);
  or _41229_ (_18416_, _18415_, _18411_);
  or _41230_ (_18417_, _18416_, _05920_);
  and _41231_ (_18418_, _18417_, _05933_);
  and _41232_ (_18419_, _18418_, _18407_);
  or _41233_ (_18420_, _18419_, _18397_);
  and _41234_ (_18421_, _18420_, _06071_);
  and _41235_ (_18422_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _41236_ (_18423_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _41237_ (_18424_, _18423_, _18422_);
  and _41238_ (_18425_, _18424_, _05996_);
  and _41239_ (_18426_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _41240_ (_18427_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or _41241_ (_18428_, _18427_, _18426_);
  and _41242_ (_18429_, _18428_, _05997_);
  or _41243_ (_18430_, _18429_, _18425_);
  or _41244_ (_18431_, _18430_, _06021_);
  and _41245_ (_18432_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _41246_ (_18433_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _41247_ (_18434_, _18433_, _18432_);
  and _41248_ (_18435_, _18434_, _05996_);
  and _41249_ (_18436_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _41250_ (_18437_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or _41251_ (_18438_, _18437_, _18436_);
  and _41252_ (_18439_, _18438_, _05997_);
  or _41253_ (_18440_, _18439_, _18435_);
  or _41254_ (_18441_, _18440_, _05920_);
  and _41255_ (_18442_, _18441_, _06033_);
  and _41256_ (_18443_, _18442_, _18431_);
  or _41257_ (_18444_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _41258_ (_18445_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _41259_ (_18446_, _18445_, _18444_);
  and _41260_ (_18447_, _18446_, _05996_);
  or _41261_ (_18448_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _41262_ (_18449_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _41263_ (_18450_, _18449_, _18448_);
  and _41264_ (_18451_, _18450_, _05997_);
  or _41265_ (_18452_, _18451_, _18447_);
  or _41266_ (_18453_, _18452_, _06021_);
  or _41267_ (_18454_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or _41268_ (_18455_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _41269_ (_18456_, _18455_, _18454_);
  and _41270_ (_18457_, _18456_, _05996_);
  or _41271_ (_18458_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _41272_ (_18459_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _41273_ (_18460_, _18459_, _18458_);
  and _41274_ (_18461_, _18460_, _05997_);
  or _41275_ (_18462_, _18461_, _18457_);
  or _41276_ (_18463_, _18462_, _05920_);
  and _41277_ (_18464_, _18463_, _05933_);
  and _41278_ (_18465_, _18464_, _18453_);
  or _41279_ (_18466_, _18465_, _18443_);
  and _41280_ (_18467_, _18466_, _05776_);
  or _41281_ (_18468_, _18467_, _18421_);
  and _41282_ (_18469_, _18468_, _06070_);
  or _41283_ (_18470_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or _41284_ (_18471_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _41285_ (_18472_, _18471_, _18470_);
  and _41286_ (_18473_, _18472_, _05996_);
  or _41287_ (_18474_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or _41288_ (_18475_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _41289_ (_18476_, _18475_, _18474_);
  and _41290_ (_18477_, _18476_, _05997_);
  or _41291_ (_18478_, _18477_, _18473_);
  and _41292_ (_18479_, _18478_, _06021_);
  or _41293_ (_18480_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or _41294_ (_18481_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _41295_ (_18482_, _18481_, _18480_);
  and _41296_ (_18483_, _18482_, _05996_);
  or _41297_ (_18484_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _41298_ (_18485_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and _41299_ (_18486_, _18485_, _18484_);
  and _41300_ (_18487_, _18486_, _05997_);
  or _41301_ (_18488_, _18487_, _18483_);
  and _41302_ (_18489_, _18488_, _05920_);
  or _41303_ (_18490_, _18489_, _18479_);
  and _41304_ (_18491_, _18490_, _05933_);
  and _41305_ (_18492_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _41306_ (_18493_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _41307_ (_18494_, _18493_, _18492_);
  and _41308_ (_18495_, _18494_, _05996_);
  and _41309_ (_18496_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and _41310_ (_18497_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or _41311_ (_18498_, _18497_, _18496_);
  and _41312_ (_18499_, _18498_, _05997_);
  or _41313_ (_18500_, _18499_, _18495_);
  and _41314_ (_18501_, _18500_, _06021_);
  and _41315_ (_18502_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _41316_ (_18503_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _41317_ (_18504_, _18503_, _18502_);
  and _41318_ (_18505_, _18504_, _05996_);
  and _41319_ (_18506_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and _41320_ (_18507_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or _41321_ (_18508_, _18507_, _18506_);
  and _41322_ (_18509_, _18508_, _05997_);
  or _41323_ (_18510_, _18509_, _18505_);
  and _41324_ (_18511_, _18510_, _05920_);
  or _41325_ (_18512_, _18511_, _18501_);
  and _41326_ (_18513_, _18512_, _06033_);
  or _41327_ (_18514_, _18513_, _18491_);
  and _41328_ (_18515_, _18514_, _05776_);
  or _41329_ (_18516_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _41330_ (_18517_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and _41331_ (_18518_, _18517_, _05997_);
  and _41332_ (_18519_, _18518_, _18516_);
  or _41333_ (_18520_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _41334_ (_18521_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _41335_ (_18522_, _18521_, _05996_);
  and _41336_ (_18523_, _18522_, _18520_);
  or _41337_ (_18524_, _18523_, _18519_);
  and _41338_ (_18525_, _18524_, _06021_);
  or _41339_ (_18526_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _41340_ (_18527_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and _41341_ (_18528_, _18527_, _05997_);
  and _41342_ (_18529_, _18528_, _18526_);
  or _41343_ (_18530_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _41344_ (_18531_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and _41345_ (_18532_, _18531_, _05996_);
  and _41346_ (_18533_, _18532_, _18530_);
  or _41347_ (_18534_, _18533_, _18529_);
  and _41348_ (_18535_, _18534_, _05920_);
  or _41349_ (_18536_, _18535_, _18525_);
  and _41350_ (_18537_, _18536_, _05933_);
  and _41351_ (_18538_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and _41352_ (_18539_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _41353_ (_18540_, _18539_, _18538_);
  and _41354_ (_18541_, _18540_, _05996_);
  and _41355_ (_18542_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _41356_ (_18543_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _41357_ (_18544_, _18543_, _18542_);
  and _41358_ (_18545_, _18544_, _05997_);
  or _41359_ (_18546_, _18545_, _18541_);
  and _41360_ (_18547_, _18546_, _06021_);
  and _41361_ (_18548_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _41362_ (_18549_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _41363_ (_18550_, _18549_, _18548_);
  and _41364_ (_18551_, _18550_, _05996_);
  and _41365_ (_18552_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and _41366_ (_18553_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _41367_ (_18554_, _18553_, _18552_);
  and _41368_ (_18555_, _18554_, _05997_);
  or _41369_ (_18556_, _18555_, _18551_);
  and _41370_ (_18557_, _18556_, _05920_);
  or _41371_ (_18558_, _18557_, _18547_);
  and _41372_ (_18559_, _18558_, _06033_);
  or _41373_ (_18560_, _18559_, _18537_);
  and _41374_ (_18561_, _18560_, _06071_);
  or _41375_ (_18562_, _18561_, _18515_);
  and _41376_ (_18563_, _18562_, _05822_);
  or _41377_ (_18564_, _18563_, _18469_);
  or _41378_ (_18565_, _18564_, _06616_);
  and _41379_ (_18566_, _18565_, _18375_);
  or _41380_ (_18567_, _18566_, _05584_);
  and _41381_ (_18568_, _18567_, _18185_);
  or _41382_ (_18569_, _18568_, _06019_);
  or _41383_ (_18570_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _41384_ (_18571_, _18570_, _25365_);
  and _41385_ (_14805_, _18571_, _18569_);
  and _41386_ (_18572_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _41387_ (_18573_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _41388_ (_18574_, _18573_, _18572_);
  and _41389_ (_18575_, _18574_, _05996_);
  and _41390_ (_18576_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and _41391_ (_18577_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _41392_ (_18578_, _18577_, _18576_);
  and _41393_ (_18579_, _18578_, _05997_);
  or _41394_ (_18580_, _18579_, _18575_);
  or _41395_ (_18581_, _18580_, _06021_);
  and _41396_ (_18582_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and _41397_ (_18583_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _41398_ (_18584_, _18583_, _18582_);
  and _41399_ (_18585_, _18584_, _05996_);
  and _41400_ (_18586_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and _41401_ (_18587_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _41402_ (_18588_, _18587_, _18586_);
  and _41403_ (_18589_, _18588_, _05997_);
  or _41404_ (_18590_, _18589_, _18585_);
  or _41405_ (_18591_, _18590_, _05920_);
  and _41406_ (_18592_, _18591_, _06033_);
  and _41407_ (_18593_, _18592_, _18581_);
  or _41408_ (_18594_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _41409_ (_18595_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and _41410_ (_18596_, _18595_, _18594_);
  and _41411_ (_18597_, _18596_, _05996_);
  or _41412_ (_18598_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _41413_ (_18599_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and _41414_ (_18600_, _18599_, _18598_);
  and _41415_ (_18601_, _18600_, _05997_);
  or _41416_ (_18602_, _18601_, _18597_);
  or _41417_ (_18603_, _18602_, _06021_);
  or _41418_ (_18604_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _41419_ (_18605_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and _41420_ (_18606_, _18605_, _18604_);
  and _41421_ (_18607_, _18606_, _05996_);
  or _41422_ (_18608_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _41423_ (_18609_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and _41424_ (_18610_, _18609_, _18608_);
  and _41425_ (_18611_, _18610_, _05997_);
  or _41426_ (_18612_, _18611_, _18607_);
  or _41427_ (_18613_, _18612_, _05920_);
  and _41428_ (_18614_, _18613_, _05933_);
  and _41429_ (_18615_, _18614_, _18603_);
  or _41430_ (_18616_, _18615_, _18593_);
  and _41431_ (_18617_, _18616_, _05776_);
  and _41432_ (_18618_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and _41433_ (_18619_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _41434_ (_18620_, _18619_, _18618_);
  and _41435_ (_18621_, _18620_, _05996_);
  and _41436_ (_18622_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and _41437_ (_18623_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _41438_ (_18624_, _18623_, _18622_);
  and _41439_ (_18625_, _18624_, _05997_);
  or _41440_ (_18626_, _18625_, _18621_);
  or _41441_ (_18627_, _18626_, _06021_);
  and _41442_ (_18628_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and _41443_ (_18629_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _41444_ (_18630_, _18629_, _18628_);
  and _41445_ (_18631_, _18630_, _05996_);
  and _41446_ (_18632_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and _41447_ (_18633_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _41448_ (_18634_, _18633_, _18632_);
  and _41449_ (_18635_, _18634_, _05997_);
  or _41450_ (_18636_, _18635_, _18631_);
  or _41451_ (_18637_, _18636_, _05920_);
  and _41452_ (_18638_, _18637_, _06033_);
  and _41453_ (_18639_, _18638_, _18627_);
  or _41454_ (_18640_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _41455_ (_18641_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and _41456_ (_18642_, _18641_, _05997_);
  and _41457_ (_18643_, _18642_, _18640_);
  or _41458_ (_18644_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _41459_ (_18645_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and _41460_ (_18646_, _18645_, _05996_);
  and _41461_ (_18647_, _18646_, _18644_);
  or _41462_ (_18648_, _18647_, _18643_);
  or _41463_ (_18649_, _18648_, _06021_);
  or _41464_ (_18650_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _41465_ (_18651_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and _41466_ (_18652_, _18651_, _05997_);
  and _41467_ (_18653_, _18652_, _18650_);
  or _41468_ (_18654_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _41469_ (_18655_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and _41470_ (_18656_, _18655_, _05996_);
  and _41471_ (_18657_, _18656_, _18654_);
  or _41472_ (_18658_, _18657_, _18653_);
  or _41473_ (_18659_, _18658_, _05920_);
  and _41474_ (_18660_, _18659_, _05933_);
  and _41475_ (_18661_, _18660_, _18649_);
  or _41476_ (_18662_, _18661_, _18639_);
  and _41477_ (_18663_, _18662_, _06071_);
  or _41478_ (_18664_, _18663_, _18617_);
  and _41479_ (_18665_, _18664_, _06070_);
  and _41480_ (_18666_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and _41481_ (_18667_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _41482_ (_18668_, _18667_, _18666_);
  and _41483_ (_18669_, _18668_, _05996_);
  and _41484_ (_18670_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and _41485_ (_18671_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _41486_ (_18672_, _18671_, _18670_);
  and _41487_ (_18673_, _18672_, _05997_);
  or _41488_ (_18674_, _18673_, _18669_);
  and _41489_ (_18675_, _18674_, _05920_);
  and _41490_ (_18676_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and _41491_ (_18677_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _41492_ (_18678_, _18677_, _18676_);
  and _41493_ (_18679_, _18678_, _05996_);
  and _41494_ (_18680_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _41495_ (_18681_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _41496_ (_18682_, _18681_, _18680_);
  and _41497_ (_18683_, _18682_, _05997_);
  or _41498_ (_18684_, _18683_, _18679_);
  and _41499_ (_18685_, _18684_, _06021_);
  or _41500_ (_18686_, _18685_, _18675_);
  and _41501_ (_18687_, _18686_, _06033_);
  or _41502_ (_18688_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _41503_ (_18689_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _41504_ (_18690_, _18689_, _05997_);
  and _41505_ (_18691_, _18690_, _18688_);
  or _41506_ (_18692_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _41507_ (_18693_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _41508_ (_18694_, _18693_, _05996_);
  and _41509_ (_18695_, _18694_, _18692_);
  or _41510_ (_18696_, _18695_, _18691_);
  and _41511_ (_18697_, _18696_, _05920_);
  or _41512_ (_18698_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _41513_ (_18699_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _41514_ (_18700_, _18699_, _05997_);
  and _41515_ (_18701_, _18700_, _18698_);
  or _41516_ (_18702_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _41517_ (_18703_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _41518_ (_18704_, _18703_, _05996_);
  and _41519_ (_18705_, _18704_, _18702_);
  or _41520_ (_18706_, _18705_, _18701_);
  and _41521_ (_18707_, _18706_, _06021_);
  or _41522_ (_18708_, _18707_, _18697_);
  and _41523_ (_18709_, _18708_, _05933_);
  or _41524_ (_18710_, _18709_, _18687_);
  and _41525_ (_18711_, _18710_, _06071_);
  and _41526_ (_18712_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and _41527_ (_18713_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _41528_ (_18714_, _18713_, _18712_);
  and _41529_ (_18715_, _18714_, _05996_);
  and _41530_ (_18716_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and _41531_ (_18717_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _41532_ (_18718_, _18717_, _18716_);
  and _41533_ (_18719_, _18718_, _05997_);
  or _41534_ (_18720_, _18719_, _18715_);
  and _41535_ (_18721_, _18720_, _05920_);
  and _41536_ (_18722_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and _41537_ (_18723_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _41538_ (_18724_, _18723_, _18722_);
  and _41539_ (_18725_, _18724_, _05996_);
  and _41540_ (_18726_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and _41541_ (_18727_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _41542_ (_18728_, _18727_, _18726_);
  and _41543_ (_18729_, _18728_, _05997_);
  or _41544_ (_18730_, _18729_, _18725_);
  and _41545_ (_18731_, _18730_, _06021_);
  or _41546_ (_18732_, _18731_, _18721_);
  and _41547_ (_18733_, _18732_, _06033_);
  or _41548_ (_18734_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _41549_ (_18735_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and _41550_ (_18736_, _18735_, _18734_);
  and _41551_ (_18737_, _18736_, _05996_);
  or _41552_ (_18738_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _41553_ (_18739_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and _41554_ (_18740_, _18739_, _18738_);
  and _41555_ (_18741_, _18740_, _05997_);
  or _41556_ (_18742_, _18741_, _18737_);
  and _41557_ (_18743_, _18742_, _05920_);
  or _41558_ (_18744_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _41559_ (_18745_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and _41560_ (_18746_, _18745_, _18744_);
  and _41561_ (_18747_, _18746_, _05996_);
  or _41562_ (_18748_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _41563_ (_18749_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and _41564_ (_18750_, _18749_, _18748_);
  and _41565_ (_18751_, _18750_, _05997_);
  or _41566_ (_18752_, _18751_, _18747_);
  and _41567_ (_18753_, _18752_, _06021_);
  or _41568_ (_18754_, _18753_, _18743_);
  and _41569_ (_18755_, _18754_, _05933_);
  or _41570_ (_18756_, _18755_, _18733_);
  and _41571_ (_18757_, _18756_, _05776_);
  or _41572_ (_18758_, _18757_, _18711_);
  and _41573_ (_18759_, _18758_, _05822_);
  or _41574_ (_18760_, _18759_, _18665_);
  or _41575_ (_18761_, _18760_, _05868_);
  and _41576_ (_18762_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and _41577_ (_18763_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _41578_ (_18764_, _18763_, _18762_);
  and _41579_ (_18765_, _18764_, _05996_);
  and _41580_ (_18766_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and _41581_ (_18767_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _41582_ (_18768_, _18767_, _18766_);
  and _41583_ (_18769_, _18768_, _05997_);
  or _41584_ (_18770_, _18769_, _18765_);
  or _41585_ (_18771_, _18770_, _06021_);
  and _41586_ (_18772_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and _41587_ (_18773_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _41588_ (_18774_, _18773_, _18772_);
  and _41589_ (_18775_, _18774_, _05996_);
  and _41590_ (_18776_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and _41591_ (_18777_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _41592_ (_18778_, _18777_, _18776_);
  and _41593_ (_18779_, _18778_, _05997_);
  or _41594_ (_18780_, _18779_, _18775_);
  or _41595_ (_18781_, _18780_, _05920_);
  and _41596_ (_18782_, _18781_, _06033_);
  and _41597_ (_18783_, _18782_, _18771_);
  or _41598_ (_18784_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _41599_ (_18785_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and _41600_ (_18786_, _18785_, _05997_);
  and _41601_ (_18787_, _18786_, _18784_);
  or _41602_ (_18788_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _41603_ (_18789_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and _41604_ (_18790_, _18789_, _05996_);
  and _41605_ (_18791_, _18790_, _18788_);
  or _41606_ (_18792_, _18791_, _18787_);
  or _41607_ (_18793_, _18792_, _06021_);
  or _41608_ (_18794_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _41609_ (_18795_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and _41610_ (_18796_, _18795_, _05997_);
  and _41611_ (_18797_, _18796_, _18794_);
  or _41612_ (_18798_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _41613_ (_18799_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and _41614_ (_18800_, _18799_, _05996_);
  and _41615_ (_18801_, _18800_, _18798_);
  or _41616_ (_18802_, _18801_, _18797_);
  or _41617_ (_18803_, _18802_, _05920_);
  and _41618_ (_18804_, _18803_, _05933_);
  and _41619_ (_18805_, _18804_, _18793_);
  or _41620_ (_18806_, _18805_, _18783_);
  and _41621_ (_18807_, _18806_, _06071_);
  and _41622_ (_18808_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _41623_ (_18809_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _41624_ (_18810_, _18809_, _18808_);
  and _41625_ (_18811_, _18810_, _05996_);
  and _41626_ (_18812_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and _41627_ (_18813_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _41628_ (_18814_, _18813_, _18812_);
  and _41629_ (_18815_, _18814_, _05997_);
  or _41630_ (_18816_, _18815_, _18811_);
  or _41631_ (_18817_, _18816_, _06021_);
  and _41632_ (_18818_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and _41633_ (_18819_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _41634_ (_18820_, _18819_, _18818_);
  and _41635_ (_18821_, _18820_, _05996_);
  and _41636_ (_18822_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _41637_ (_18823_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _41638_ (_18824_, _18823_, _18822_);
  and _41639_ (_18825_, _18824_, _05997_);
  or _41640_ (_18826_, _18825_, _18821_);
  or _41641_ (_18827_, _18826_, _05920_);
  and _41642_ (_18828_, _18827_, _06033_);
  and _41643_ (_18829_, _18828_, _18817_);
  or _41644_ (_18830_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _41645_ (_18831_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _41646_ (_18832_, _18831_, _18830_);
  and _41647_ (_18833_, _18832_, _05996_);
  or _41648_ (_18834_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _41649_ (_18835_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and _41650_ (_18836_, _18835_, _18834_);
  and _41651_ (_18837_, _18836_, _05997_);
  or _41652_ (_18838_, _18837_, _18833_);
  or _41653_ (_18839_, _18838_, _06021_);
  or _41654_ (_18840_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _41655_ (_18841_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and _41656_ (_18842_, _18841_, _18840_);
  and _41657_ (_18843_, _18842_, _05996_);
  or _41658_ (_18844_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _41659_ (_18845_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and _41660_ (_18846_, _18845_, _18844_);
  and _41661_ (_18847_, _18846_, _05997_);
  or _41662_ (_18848_, _18847_, _18843_);
  or _41663_ (_18849_, _18848_, _05920_);
  and _41664_ (_18850_, _18849_, _05933_);
  and _41665_ (_18851_, _18850_, _18839_);
  or _41666_ (_18852_, _18851_, _18829_);
  and _41667_ (_18853_, _18852_, _05776_);
  or _41668_ (_18854_, _18853_, _18807_);
  and _41669_ (_18855_, _18854_, _06070_);
  or _41670_ (_18856_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _41671_ (_18857_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and _41672_ (_18858_, _18857_, _18856_);
  and _41673_ (_18859_, _18858_, _05996_);
  or _41674_ (_18860_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _41675_ (_18861_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and _41676_ (_18862_, _18861_, _18860_);
  and _41677_ (_18863_, _18862_, _05997_);
  or _41678_ (_18864_, _18863_, _18859_);
  and _41679_ (_18865_, _18864_, _06021_);
  or _41680_ (_18866_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _41681_ (_18867_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and _41682_ (_18868_, _18867_, _18866_);
  and _41683_ (_18869_, _18868_, _05996_);
  or _41684_ (_18870_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _41685_ (_18871_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and _41686_ (_18872_, _18871_, _18870_);
  and _41687_ (_18873_, _18872_, _05997_);
  or _41688_ (_18874_, _18873_, _18869_);
  and _41689_ (_18875_, _18874_, _05920_);
  or _41690_ (_18876_, _18875_, _18865_);
  and _41691_ (_18877_, _18876_, _05933_);
  and _41692_ (_18878_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and _41693_ (_18879_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _41694_ (_18880_, _18879_, _18878_);
  and _41695_ (_18881_, _18880_, _05996_);
  and _41696_ (_18882_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and _41697_ (_18883_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _41698_ (_18884_, _18883_, _18882_);
  and _41699_ (_18885_, _18884_, _05997_);
  or _41700_ (_18886_, _18885_, _18881_);
  and _41701_ (_18887_, _18886_, _06021_);
  and _41702_ (_18888_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and _41703_ (_18889_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _41704_ (_18890_, _18889_, _18888_);
  and _41705_ (_18891_, _18890_, _05996_);
  and _41706_ (_18892_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and _41707_ (_18893_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _41708_ (_18894_, _18893_, _18892_);
  and _41709_ (_18895_, _18894_, _05997_);
  or _41710_ (_18896_, _18895_, _18891_);
  and _41711_ (_18897_, _18896_, _05920_);
  or _41712_ (_18898_, _18897_, _18887_);
  and _41713_ (_18899_, _18898_, _06033_);
  or _41714_ (_18900_, _18899_, _18877_);
  and _41715_ (_18901_, _18900_, _05776_);
  or _41716_ (_18902_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or _41717_ (_18903_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and _41718_ (_18904_, _18903_, _05997_);
  and _41719_ (_18905_, _18904_, _18902_);
  or _41720_ (_18906_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or _41721_ (_18907_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and _41722_ (_18908_, _18907_, _05996_);
  and _41723_ (_18909_, _18908_, _18906_);
  or _41724_ (_18910_, _18909_, _18905_);
  and _41725_ (_18911_, _18910_, _06021_);
  or _41726_ (_18912_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or _41727_ (_18913_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and _41728_ (_18914_, _18913_, _05997_);
  and _41729_ (_18915_, _18914_, _18912_);
  or _41730_ (_18916_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or _41731_ (_18917_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and _41732_ (_18918_, _18917_, _05996_);
  and _41733_ (_18919_, _18918_, _18916_);
  or _41734_ (_18920_, _18919_, _18915_);
  and _41735_ (_18921_, _18920_, _05920_);
  or _41736_ (_18922_, _18921_, _18911_);
  and _41737_ (_18923_, _18922_, _05933_);
  and _41738_ (_18924_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and _41739_ (_18925_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or _41740_ (_18926_, _18925_, _18924_);
  and _41741_ (_18927_, _18926_, _05996_);
  and _41742_ (_18928_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and _41743_ (_18929_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or _41744_ (_18930_, _18929_, _18928_);
  and _41745_ (_18931_, _18930_, _05997_);
  or _41746_ (_18932_, _18931_, _18927_);
  and _41747_ (_18933_, _18932_, _06021_);
  and _41748_ (_18934_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and _41749_ (_18935_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or _41750_ (_18936_, _18935_, _18934_);
  and _41751_ (_18937_, _18936_, _05996_);
  and _41752_ (_18938_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and _41753_ (_18939_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or _41754_ (_18940_, _18939_, _18938_);
  and _41755_ (_18941_, _18940_, _05997_);
  or _41756_ (_18942_, _18941_, _18937_);
  and _41757_ (_18943_, _18942_, _05920_);
  or _41758_ (_18944_, _18943_, _18933_);
  and _41759_ (_18945_, _18944_, _06033_);
  or _41760_ (_18946_, _18945_, _18923_);
  and _41761_ (_18947_, _18946_, _06071_);
  or _41762_ (_18948_, _18947_, _18901_);
  and _41763_ (_18949_, _18948_, _05822_);
  or _41764_ (_18950_, _18949_, _18855_);
  or _41765_ (_18951_, _18950_, _06616_);
  and _41766_ (_18952_, _18951_, _18761_);
  or _41767_ (_18953_, _18952_, _06020_);
  and _41768_ (_18954_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _41769_ (_18955_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or _41770_ (_18956_, _18955_, _18954_);
  and _41771_ (_18957_, _18956_, _05996_);
  and _41772_ (_18958_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _41773_ (_18959_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _41774_ (_18960_, _18959_, _18958_);
  and _41775_ (_18961_, _18960_, _05997_);
  or _41776_ (_18962_, _18961_, _18957_);
  and _41777_ (_18963_, _18962_, _05920_);
  and _41778_ (_18964_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _41779_ (_18965_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or _41780_ (_18966_, _18965_, _18964_);
  and _41781_ (_18967_, _18966_, _05996_);
  and _41782_ (_18968_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _41783_ (_18969_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _41784_ (_18970_, _18969_, _18968_);
  and _41785_ (_18971_, _18970_, _05997_);
  or _41786_ (_18972_, _18971_, _18967_);
  and _41787_ (_18973_, _18972_, _06021_);
  or _41788_ (_18974_, _18973_, _18963_);
  and _41789_ (_18975_, _18974_, _06033_);
  or _41790_ (_18976_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or _41791_ (_18977_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _41792_ (_18978_, _18977_, _05997_);
  and _41793_ (_18979_, _18978_, _18976_);
  or _41794_ (_18980_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _41795_ (_18981_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _41796_ (_18982_, _18981_, _05996_);
  and _41797_ (_18983_, _18982_, _18980_);
  or _41798_ (_18984_, _18983_, _18979_);
  and _41799_ (_18985_, _18984_, _05920_);
  or _41800_ (_18986_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or _41801_ (_18987_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _41802_ (_18988_, _18987_, _05997_);
  and _41803_ (_18989_, _18988_, _18986_);
  or _41804_ (_18990_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _41805_ (_18991_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and _41806_ (_18992_, _18991_, _05996_);
  and _41807_ (_18993_, _18992_, _18990_);
  or _41808_ (_18994_, _18993_, _18989_);
  and _41809_ (_18995_, _18994_, _06021_);
  or _41810_ (_18996_, _18995_, _18985_);
  and _41811_ (_18997_, _18996_, _05933_);
  or _41812_ (_18998_, _18997_, _18975_);
  and _41813_ (_18999_, _18998_, _06071_);
  and _41814_ (_19000_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and _41815_ (_19001_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _41816_ (_19002_, _19001_, _19000_);
  and _41817_ (_19003_, _19002_, _05996_);
  and _41818_ (_19004_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and _41819_ (_19005_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _41820_ (_19006_, _19005_, _19004_);
  and _41821_ (_19007_, _19006_, _05997_);
  or _41822_ (_19008_, _19007_, _19003_);
  and _41823_ (_19009_, _19008_, _05920_);
  and _41824_ (_19010_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and _41825_ (_19011_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _41826_ (_19012_, _19011_, _19010_);
  and _41827_ (_19013_, _19012_, _05996_);
  and _41828_ (_19014_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and _41829_ (_19015_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _41830_ (_19016_, _19015_, _19014_);
  and _41831_ (_19017_, _19016_, _05997_);
  or _41832_ (_19018_, _19017_, _19013_);
  and _41833_ (_19019_, _19018_, _06021_);
  or _41834_ (_19020_, _19019_, _19009_);
  and _41835_ (_19021_, _19020_, _06033_);
  or _41836_ (_19022_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _41837_ (_19023_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _41838_ (_19024_, _19023_, _19022_);
  and _41839_ (_19025_, _19024_, _05996_);
  or _41840_ (_19026_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _41841_ (_19027_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and _41842_ (_19028_, _19027_, _19026_);
  and _41843_ (_19029_, _19028_, _05997_);
  or _41844_ (_19030_, _19029_, _19025_);
  and _41845_ (_19031_, _19030_, _05920_);
  or _41846_ (_19032_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _41847_ (_19033_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and _41848_ (_19034_, _19033_, _19032_);
  and _41849_ (_19035_, _19034_, _05996_);
  or _41850_ (_19036_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _41851_ (_19037_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and _41852_ (_19038_, _19037_, _19036_);
  and _41853_ (_19039_, _19038_, _05997_);
  or _41854_ (_19040_, _19039_, _19035_);
  and _41855_ (_19041_, _19040_, _06021_);
  or _41856_ (_19042_, _19041_, _19031_);
  and _41857_ (_19043_, _19042_, _05933_);
  or _41858_ (_19044_, _19043_, _19021_);
  and _41859_ (_19045_, _19044_, _05776_);
  or _41860_ (_19046_, _19045_, _18999_);
  and _41861_ (_19047_, _19046_, _05822_);
  and _41862_ (_19048_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and _41863_ (_19049_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _41864_ (_19050_, _19049_, _19048_);
  and _41865_ (_19051_, _19050_, _05996_);
  and _41866_ (_19052_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and _41867_ (_19053_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _41868_ (_19054_, _19053_, _19052_);
  and _41869_ (_19055_, _19054_, _05997_);
  or _41870_ (_19056_, _19055_, _19051_);
  or _41871_ (_19057_, _19056_, _06021_);
  and _41872_ (_19058_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and _41873_ (_19059_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _41874_ (_19060_, _19059_, _19058_);
  and _41875_ (_19061_, _19060_, _05996_);
  and _41876_ (_19062_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and _41877_ (_19063_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _41878_ (_19064_, _19063_, _19062_);
  and _41879_ (_19065_, _19064_, _05997_);
  or _41880_ (_19066_, _19065_, _19061_);
  or _41881_ (_19067_, _19066_, _05920_);
  and _41882_ (_19068_, _19067_, _06033_);
  and _41883_ (_19069_, _19068_, _19057_);
  or _41884_ (_19070_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _41885_ (_19071_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and _41886_ (_19072_, _19071_, _19070_);
  and _41887_ (_19073_, _19072_, _05996_);
  or _41888_ (_19074_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _41889_ (_19075_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and _41890_ (_19076_, _19075_, _19074_);
  and _41891_ (_19077_, _19076_, _05997_);
  or _41892_ (_19078_, _19077_, _19073_);
  or _41893_ (_19079_, _19078_, _06021_);
  or _41894_ (_19080_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _41895_ (_19081_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and _41896_ (_19082_, _19081_, _19080_);
  and _41897_ (_19083_, _19082_, _05996_);
  or _41898_ (_19084_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _41899_ (_19085_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and _41900_ (_19086_, _19085_, _19084_);
  and _41901_ (_19087_, _19086_, _05997_);
  or _41902_ (_19088_, _19087_, _19083_);
  or _41903_ (_19089_, _19088_, _05920_);
  and _41904_ (_19090_, _19089_, _05933_);
  and _41905_ (_19091_, _19090_, _19079_);
  or _41906_ (_19092_, _19091_, _19069_);
  and _41907_ (_19093_, _19092_, _05776_);
  and _41908_ (_19094_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _41909_ (_19095_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _41910_ (_19096_, _19095_, _19094_);
  and _41911_ (_19097_, _19096_, _05996_);
  and _41912_ (_19098_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and _41913_ (_19099_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or _41914_ (_19100_, _19099_, _19098_);
  and _41915_ (_19101_, _19100_, _05997_);
  or _41916_ (_19102_, _19101_, _19097_);
  or _41917_ (_19103_, _19102_, _06021_);
  and _41918_ (_19104_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and _41919_ (_19105_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _41920_ (_19106_, _19105_, _19104_);
  and _41921_ (_19107_, _19106_, _05996_);
  and _41922_ (_19108_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _41923_ (_19109_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _41924_ (_19110_, _19109_, _19108_);
  and _41925_ (_19111_, _19110_, _05997_);
  or _41926_ (_19112_, _19111_, _19107_);
  or _41927_ (_19113_, _19112_, _05920_);
  and _41928_ (_19114_, _19113_, _06033_);
  and _41929_ (_19115_, _19114_, _19103_);
  or _41930_ (_19116_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or _41931_ (_19117_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _41932_ (_19118_, _19117_, _05997_);
  and _41933_ (_19119_, _19118_, _19116_);
  or _41934_ (_19120_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _41935_ (_19121_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _41936_ (_19122_, _19121_, _05996_);
  and _41937_ (_19123_, _19122_, _19120_);
  or _41938_ (_19124_, _19123_, _19119_);
  or _41939_ (_19125_, _19124_, _06021_);
  or _41940_ (_19126_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _41941_ (_19127_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and _41942_ (_19128_, _19127_, _05997_);
  and _41943_ (_19129_, _19128_, _19126_);
  or _41944_ (_19130_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or _41945_ (_19131_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _41946_ (_19132_, _19131_, _05996_);
  and _41947_ (_19133_, _19132_, _19130_);
  or _41948_ (_19134_, _19133_, _19129_);
  or _41949_ (_19135_, _19134_, _05920_);
  and _41950_ (_19136_, _19135_, _05933_);
  and _41951_ (_19137_, _19136_, _19125_);
  or _41952_ (_19138_, _19137_, _19115_);
  and _41953_ (_19139_, _19138_, _06071_);
  or _41954_ (_19140_, _19139_, _19093_);
  and _41955_ (_19141_, _19140_, _06070_);
  or _41956_ (_19142_, _19141_, _19047_);
  or _41957_ (_19143_, _19142_, _05868_);
  and _41958_ (_19144_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and _41959_ (_19145_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _41960_ (_19146_, _19145_, _19144_);
  and _41961_ (_19147_, _19146_, _05997_);
  and _41962_ (_19148_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and _41963_ (_19149_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _41964_ (_19150_, _19149_, _19148_);
  and _41965_ (_19151_, _19150_, _05996_);
  or _41966_ (_19152_, _19151_, _19147_);
  or _41967_ (_19153_, _19152_, _06021_);
  and _41968_ (_19154_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and _41969_ (_19155_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _41970_ (_19156_, _19155_, _19154_);
  and _41971_ (_19157_, _19156_, _05997_);
  and _41972_ (_19158_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and _41973_ (_19159_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _41974_ (_19160_, _19159_, _19158_);
  and _41975_ (_19161_, _19160_, _05996_);
  or _41976_ (_19162_, _19161_, _19157_);
  or _41977_ (_19163_, _19162_, _05920_);
  and _41978_ (_19164_, _19163_, _06033_);
  and _41979_ (_19165_, _19164_, _19153_);
  or _41980_ (_19166_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _41981_ (_19167_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and _41982_ (_19168_, _19167_, _05996_);
  and _41983_ (_19169_, _19168_, _19166_);
  or _41984_ (_19170_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _41985_ (_19171_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and _41986_ (_19172_, _19171_, _05997_);
  and _41987_ (_19173_, _19172_, _19170_);
  or _41988_ (_19174_, _19173_, _19169_);
  or _41989_ (_19175_, _19174_, _06021_);
  or _41990_ (_19176_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _41991_ (_19177_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and _41992_ (_19178_, _19177_, _05996_);
  and _41993_ (_19179_, _19178_, _19176_);
  or _41994_ (_19180_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _41995_ (_19181_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and _41996_ (_19182_, _19181_, _05997_);
  and _41997_ (_19183_, _19182_, _19180_);
  or _41998_ (_19184_, _19183_, _19179_);
  or _41999_ (_19185_, _19184_, _05920_);
  and _42000_ (_19186_, _19185_, _05933_);
  and _42001_ (_19187_, _19186_, _19175_);
  or _42002_ (_19188_, _19187_, _19165_);
  and _42003_ (_19189_, _19188_, _06071_);
  and _42004_ (_19190_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _42005_ (_19191_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or _42006_ (_19192_, _19191_, _05996_);
  or _42007_ (_19193_, _19192_, _19190_);
  and _42008_ (_19194_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _42009_ (_19195_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _42010_ (_19196_, _19195_, _05997_);
  or _42011_ (_19197_, _19196_, _19194_);
  and _42012_ (_19198_, _19197_, _19193_);
  or _42013_ (_19199_, _19198_, _06021_);
  and _42014_ (_19200_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _42015_ (_19201_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _42016_ (_19202_, _19201_, _05996_);
  or _42017_ (_19203_, _19202_, _19200_);
  and _42018_ (_19204_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _42019_ (_19205_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or _42020_ (_19206_, _19205_, _05997_);
  or _42021_ (_19207_, _19206_, _19204_);
  and _42022_ (_19208_, _19207_, _19203_);
  or _42023_ (_19209_, _19208_, _05920_);
  and _42024_ (_19210_, _19209_, _06033_);
  and _42025_ (_19211_, _19210_, _19199_);
  or _42026_ (_19212_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _42027_ (_19213_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _42028_ (_19214_, _19213_, _19212_);
  or _42029_ (_19215_, _19214_, _05997_);
  or _42030_ (_19216_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or _42031_ (_19217_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _42032_ (_19218_, _19217_, _19216_);
  or _42033_ (_19219_, _19218_, _05996_);
  and _42034_ (_19220_, _19219_, _19215_);
  or _42035_ (_19221_, _19220_, _06021_);
  or _42036_ (_19222_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _42037_ (_19223_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _42038_ (_19224_, _19223_, _19222_);
  or _42039_ (_19225_, _19224_, _05997_);
  or _42040_ (_19226_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _42041_ (_19227_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _42042_ (_19228_, _19227_, _19226_);
  or _42043_ (_19229_, _19228_, _05996_);
  and _42044_ (_19230_, _19229_, _19225_);
  or _42045_ (_19231_, _19230_, _05920_);
  and _42046_ (_19232_, _19231_, _05933_);
  and _42047_ (_19233_, _19232_, _19221_);
  or _42048_ (_19234_, _19233_, _19211_);
  and _42049_ (_19235_, _19234_, _05776_);
  or _42050_ (_19236_, _19235_, _19189_);
  and _42051_ (_19237_, _19236_, _06070_);
  and _42052_ (_19238_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _42053_ (_19239_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or _42054_ (_19240_, _19239_, _19238_);
  and _42055_ (_19241_, _19240_, _05996_);
  and _42056_ (_19242_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _42057_ (_19243_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _42058_ (_19244_, _19243_, _19242_);
  and _42059_ (_19245_, _19244_, _05997_);
  or _42060_ (_19246_, _19245_, _19241_);
  and _42061_ (_19247_, _19246_, _05920_);
  and _42062_ (_19248_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _42063_ (_19249_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _42064_ (_19250_, _19249_, _19248_);
  and _42065_ (_19251_, _19250_, _05996_);
  and _42066_ (_19252_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _42067_ (_19253_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or _42068_ (_19254_, _19253_, _19252_);
  and _42069_ (_19255_, _19254_, _05997_);
  or _42070_ (_19256_, _19255_, _19251_);
  and _42071_ (_19257_, _19256_, _06021_);
  or _42072_ (_19258_, _19257_, _19247_);
  and _42073_ (_19259_, _19258_, _06033_);
  or _42074_ (_19260_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or _42075_ (_19261_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and _42076_ (_19262_, _19261_, _19260_);
  and _42077_ (_19263_, _19262_, _05996_);
  or _42078_ (_19264_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _42079_ (_19265_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _42080_ (_19266_, _19265_, _19264_);
  and _42081_ (_19267_, _19266_, _05997_);
  or _42082_ (_19268_, _19267_, _19263_);
  and _42083_ (_19269_, _19268_, _05920_);
  or _42084_ (_19270_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or _42085_ (_19271_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and _42086_ (_19272_, _19271_, _19270_);
  and _42087_ (_19273_, _19272_, _05996_);
  or _42088_ (_19274_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _42089_ (_19275_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _42090_ (_19276_, _19275_, _19274_);
  and _42091_ (_19277_, _19276_, _05997_);
  or _42092_ (_19278_, _19277_, _19273_);
  and _42093_ (_19279_, _19278_, _06021_);
  or _42094_ (_19280_, _19279_, _19269_);
  and _42095_ (_19281_, _19280_, _05933_);
  or _42096_ (_19282_, _19281_, _19259_);
  and _42097_ (_19283_, _19282_, _05776_);
  and _42098_ (_19284_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  and _42099_ (_19285_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or _42100_ (_19286_, _19285_, _19284_);
  and _42101_ (_19287_, _19286_, _05996_);
  and _42102_ (_19288_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  and _42103_ (_19289_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or _42104_ (_19290_, _19289_, _19288_);
  and _42105_ (_19291_, _19290_, _05997_);
  or _42106_ (_19292_, _19291_, _19287_);
  and _42107_ (_19293_, _19292_, _05920_);
  and _42108_ (_19294_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  and _42109_ (_19295_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or _42110_ (_19296_, _19295_, _19294_);
  and _42111_ (_19297_, _19296_, _05996_);
  and _42112_ (_19298_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  and _42113_ (_19299_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or _42114_ (_19300_, _19299_, _19298_);
  and _42115_ (_19301_, _19300_, _05997_);
  or _42116_ (_19302_, _19301_, _19297_);
  and _42117_ (_19303_, _19302_, _06021_);
  or _42118_ (_19304_, _19303_, _19293_);
  and _42119_ (_19305_, _19304_, _06033_);
  or _42120_ (_19306_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or _42121_ (_19307_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  and _42122_ (_19308_, _19307_, _19306_);
  and _42123_ (_19309_, _19308_, _05996_);
  or _42124_ (_19310_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or _42125_ (_19311_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  and _42126_ (_19312_, _19311_, _19310_);
  and _42127_ (_19313_, _19312_, _05997_);
  or _42128_ (_19314_, _19313_, _19309_);
  and _42129_ (_19315_, _19314_, _05920_);
  or _42130_ (_19316_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or _42131_ (_19317_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  and _42132_ (_19318_, _19317_, _19316_);
  and _42133_ (_19319_, _19318_, _05996_);
  or _42134_ (_19320_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or _42135_ (_19321_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  and _42136_ (_19322_, _19321_, _19320_);
  and _42137_ (_19323_, _19322_, _05997_);
  or _42138_ (_19324_, _19323_, _19319_);
  and _42139_ (_19325_, _19324_, _06021_);
  or _42140_ (_19326_, _19325_, _19315_);
  and _42141_ (_19327_, _19326_, _05933_);
  or _42142_ (_19328_, _19327_, _19305_);
  and _42143_ (_19329_, _19328_, _06071_);
  or _42144_ (_19330_, _19329_, _19283_);
  and _42145_ (_19331_, _19330_, _05822_);
  or _42146_ (_19332_, _19331_, _19237_);
  or _42147_ (_19333_, _19332_, _06616_);
  and _42148_ (_19334_, _19333_, _19143_);
  or _42149_ (_19335_, _19334_, _05584_);
  and _42150_ (_19336_, _19335_, _18953_);
  or _42151_ (_19337_, _19336_, _06019_);
  or _42152_ (_19338_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _42153_ (_19339_, _19338_, _25365_);
  and _42154_ (_14806_, _19339_, _19337_);
  and _42155_ (_19340_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and _42156_ (_19341_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _42157_ (_19342_, _19341_, _19340_);
  and _42158_ (_19343_, _19342_, _05996_);
  and _42159_ (_19344_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and _42160_ (_19345_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _42161_ (_19346_, _19345_, _19344_);
  and _42162_ (_19347_, _19346_, _05997_);
  or _42163_ (_19348_, _19347_, _19343_);
  or _42164_ (_19349_, _19348_, _06021_);
  and _42165_ (_19350_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and _42166_ (_19351_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _42167_ (_19352_, _19351_, _19350_);
  and _42168_ (_19353_, _19352_, _05996_);
  and _42169_ (_19354_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and _42170_ (_19355_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _42171_ (_19356_, _19355_, _19354_);
  and _42172_ (_19357_, _19356_, _05997_);
  or _42173_ (_19358_, _19357_, _19353_);
  or _42174_ (_19359_, _19358_, _05920_);
  and _42175_ (_19360_, _19359_, _06033_);
  and _42176_ (_19361_, _19360_, _19349_);
  or _42177_ (_19362_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _42178_ (_19363_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and _42179_ (_19364_, _19363_, _19362_);
  and _42180_ (_19365_, _19364_, _05996_);
  or _42181_ (_19366_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _42182_ (_19367_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and _42183_ (_19368_, _19367_, _19366_);
  and _42184_ (_19369_, _19368_, _05997_);
  or _42185_ (_19370_, _19369_, _19365_);
  or _42186_ (_19371_, _19370_, _06021_);
  or _42187_ (_19372_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _42188_ (_19373_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and _42189_ (_19374_, _19373_, _19372_);
  and _42190_ (_19375_, _19374_, _05996_);
  or _42191_ (_19376_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _42192_ (_19377_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and _42193_ (_19378_, _19377_, _19376_);
  and _42194_ (_19379_, _19378_, _05997_);
  or _42195_ (_19380_, _19379_, _19375_);
  or _42196_ (_19381_, _19380_, _05920_);
  and _42197_ (_19382_, _19381_, _05933_);
  and _42198_ (_19383_, _19382_, _19371_);
  or _42199_ (_19384_, _19383_, _19361_);
  and _42200_ (_19385_, _19384_, _05776_);
  and _42201_ (_19386_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and _42202_ (_19387_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _42203_ (_19388_, _19387_, _19386_);
  and _42204_ (_19389_, _19388_, _05996_);
  and _42205_ (_19390_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and _42206_ (_19391_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _42207_ (_19392_, _19391_, _19390_);
  and _42208_ (_19393_, _19392_, _05997_);
  or _42209_ (_19394_, _19393_, _19389_);
  or _42210_ (_19395_, _19394_, _06021_);
  and _42211_ (_19396_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and _42212_ (_19397_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _42213_ (_19398_, _19397_, _19396_);
  and _42214_ (_19399_, _19398_, _05996_);
  and _42215_ (_19400_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and _42216_ (_19401_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _42217_ (_19402_, _19401_, _19400_);
  and _42218_ (_19403_, _19402_, _05997_);
  or _42219_ (_19404_, _19403_, _19399_);
  or _42220_ (_19405_, _19404_, _05920_);
  and _42221_ (_19406_, _19405_, _06033_);
  and _42222_ (_19407_, _19406_, _19395_);
  or _42223_ (_19408_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _42224_ (_19409_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and _42225_ (_19410_, _19409_, _05997_);
  and _42226_ (_19411_, _19410_, _19408_);
  or _42227_ (_19412_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _42228_ (_19413_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and _42229_ (_19414_, _19413_, _05996_);
  and _42230_ (_19415_, _19414_, _19412_);
  or _42231_ (_19416_, _19415_, _19411_);
  or _42232_ (_19417_, _19416_, _06021_);
  or _42233_ (_19418_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _42234_ (_19419_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and _42235_ (_19420_, _19419_, _05997_);
  and _42236_ (_19421_, _19420_, _19418_);
  or _42237_ (_19422_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _42238_ (_19423_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and _42239_ (_19424_, _19423_, _05996_);
  and _42240_ (_19425_, _19424_, _19422_);
  or _42241_ (_19426_, _19425_, _19421_);
  or _42242_ (_19427_, _19426_, _05920_);
  and _42243_ (_19428_, _19427_, _05933_);
  and _42244_ (_19429_, _19428_, _19417_);
  or _42245_ (_19430_, _19429_, _19407_);
  and _42246_ (_19431_, _19430_, _06071_);
  or _42247_ (_19432_, _19431_, _19385_);
  and _42248_ (_19433_, _19432_, _06070_);
  and _42249_ (_19434_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _42250_ (_19435_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _42251_ (_19436_, _19435_, _19434_);
  and _42252_ (_19437_, _19436_, _05996_);
  and _42253_ (_19438_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _42254_ (_19439_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _42255_ (_19440_, _19439_, _19438_);
  and _42256_ (_19441_, _19440_, _05997_);
  or _42257_ (_19442_, _19441_, _19437_);
  and _42258_ (_19443_, _19442_, _05920_);
  and _42259_ (_19444_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _42260_ (_19445_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _42261_ (_19446_, _19445_, _19444_);
  and _42262_ (_19447_, _19446_, _05996_);
  and _42263_ (_19448_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _42264_ (_19449_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _42265_ (_19450_, _19449_, _19448_);
  and _42266_ (_19451_, _19450_, _05997_);
  or _42267_ (_19452_, _19451_, _19447_);
  and _42268_ (_19453_, _19452_, _06021_);
  or _42269_ (_19454_, _19453_, _19443_);
  and _42270_ (_19455_, _19454_, _06033_);
  or _42271_ (_19456_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _42272_ (_19457_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _42273_ (_19458_, _19457_, _05997_);
  and _42274_ (_19459_, _19458_, _19456_);
  or _42275_ (_19460_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _42276_ (_19461_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _42277_ (_19462_, _19461_, _05996_);
  and _42278_ (_19463_, _19462_, _19460_);
  or _42279_ (_19464_, _19463_, _19459_);
  and _42280_ (_19465_, _19464_, _05920_);
  or _42281_ (_19466_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _42282_ (_19467_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _42283_ (_19468_, _19467_, _05997_);
  and _42284_ (_19469_, _19468_, _19466_);
  or _42285_ (_19470_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _42286_ (_19471_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _42287_ (_19472_, _19471_, _05996_);
  and _42288_ (_19473_, _19472_, _19470_);
  or _42289_ (_19474_, _19473_, _19469_);
  and _42290_ (_19475_, _19474_, _06021_);
  or _42291_ (_19476_, _19475_, _19465_);
  and _42292_ (_19477_, _19476_, _05933_);
  or _42293_ (_19478_, _19477_, _19455_);
  and _42294_ (_19479_, _19478_, _06071_);
  and _42295_ (_19480_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and _42296_ (_19481_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _42297_ (_19482_, _19481_, _19480_);
  and _42298_ (_19483_, _19482_, _05996_);
  and _42299_ (_19484_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and _42300_ (_19485_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _42301_ (_19486_, _19485_, _19484_);
  and _42302_ (_19487_, _19486_, _05997_);
  or _42303_ (_19488_, _19487_, _19483_);
  and _42304_ (_19489_, _19488_, _05920_);
  and _42305_ (_19490_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and _42306_ (_19491_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _42307_ (_19492_, _19491_, _19490_);
  and _42308_ (_19493_, _19492_, _05996_);
  and _42309_ (_19494_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and _42310_ (_19495_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _42311_ (_19496_, _19495_, _19494_);
  and _42312_ (_19497_, _19496_, _05997_);
  or _42313_ (_19498_, _19497_, _19493_);
  and _42314_ (_19499_, _19498_, _06021_);
  or _42315_ (_19500_, _19499_, _19489_);
  and _42316_ (_19501_, _19500_, _06033_);
  or _42317_ (_19502_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _42318_ (_19503_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and _42319_ (_19504_, _19503_, _19502_);
  and _42320_ (_19505_, _19504_, _05996_);
  or _42321_ (_19506_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _42322_ (_19507_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and _42323_ (_19508_, _19507_, _19506_);
  and _42324_ (_19509_, _19508_, _05997_);
  or _42325_ (_19510_, _19509_, _19505_);
  and _42326_ (_19511_, _19510_, _05920_);
  or _42327_ (_19512_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _42328_ (_19513_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and _42329_ (_19514_, _19513_, _19512_);
  and _42330_ (_19515_, _19514_, _05996_);
  or _42331_ (_19516_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _42332_ (_19517_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and _42333_ (_19518_, _19517_, _19516_);
  and _42334_ (_19519_, _19518_, _05997_);
  or _42335_ (_19520_, _19519_, _19515_);
  and _42336_ (_19521_, _19520_, _06021_);
  or _42337_ (_19522_, _19521_, _19511_);
  and _42338_ (_19523_, _19522_, _05933_);
  or _42339_ (_19524_, _19523_, _19501_);
  and _42340_ (_19525_, _19524_, _05776_);
  or _42341_ (_19526_, _19525_, _19479_);
  and _42342_ (_19527_, _19526_, _05822_);
  or _42343_ (_19528_, _19527_, _19433_);
  or _42344_ (_19529_, _19528_, _05868_);
  and _42345_ (_19530_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and _42346_ (_19531_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _42347_ (_19532_, _19531_, _19530_);
  and _42348_ (_19533_, _19532_, _05996_);
  and _42349_ (_19534_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and _42350_ (_19535_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _42351_ (_19536_, _19535_, _19534_);
  and _42352_ (_19537_, _19536_, _05997_);
  or _42353_ (_19538_, _19537_, _19533_);
  or _42354_ (_19539_, _19538_, _06021_);
  and _42355_ (_19540_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and _42356_ (_19541_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _42357_ (_19542_, _19541_, _19540_);
  and _42358_ (_19543_, _19542_, _05996_);
  and _42359_ (_19544_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and _42360_ (_19545_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _42361_ (_19546_, _19545_, _19544_);
  and _42362_ (_19547_, _19546_, _05997_);
  or _42363_ (_19548_, _19547_, _19543_);
  or _42364_ (_19549_, _19548_, _05920_);
  and _42365_ (_19550_, _19549_, _06033_);
  and _42366_ (_19551_, _19550_, _19539_);
  or _42367_ (_19552_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _42368_ (_19553_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and _42369_ (_19554_, _19553_, _05997_);
  and _42370_ (_19555_, _19554_, _19552_);
  or _42371_ (_19556_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _42372_ (_19557_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and _42373_ (_19558_, _19557_, _05996_);
  and _42374_ (_19559_, _19558_, _19556_);
  or _42375_ (_19560_, _19559_, _19555_);
  or _42376_ (_19561_, _19560_, _06021_);
  or _42377_ (_19562_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _42378_ (_19563_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and _42379_ (_19564_, _19563_, _05997_);
  and _42380_ (_19565_, _19564_, _19562_);
  or _42381_ (_19566_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _42382_ (_19567_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and _42383_ (_19568_, _19567_, _05996_);
  and _42384_ (_19569_, _19568_, _19566_);
  or _42385_ (_19570_, _19569_, _19565_);
  or _42386_ (_19571_, _19570_, _05920_);
  and _42387_ (_19572_, _19571_, _05933_);
  and _42388_ (_19573_, _19572_, _19561_);
  or _42389_ (_19574_, _19573_, _19551_);
  and _42390_ (_19575_, _19574_, _06071_);
  and _42391_ (_19576_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and _42392_ (_19577_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _42393_ (_19578_, _19577_, _19576_);
  and _42394_ (_19579_, _19578_, _05996_);
  and _42395_ (_19580_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and _42396_ (_19581_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _42397_ (_19582_, _19581_, _19580_);
  and _42398_ (_19583_, _19582_, _05997_);
  or _42399_ (_19584_, _19583_, _19579_);
  or _42400_ (_19585_, _19584_, _06021_);
  and _42401_ (_19586_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _42402_ (_19587_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _42403_ (_19588_, _19587_, _19586_);
  and _42404_ (_19589_, _19588_, _05996_);
  and _42405_ (_19590_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _42406_ (_19591_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _42407_ (_19592_, _19591_, _19590_);
  and _42408_ (_19593_, _19592_, _05997_);
  or _42409_ (_19594_, _19593_, _19589_);
  or _42410_ (_19595_, _19594_, _05920_);
  and _42411_ (_19596_, _19595_, _06033_);
  and _42412_ (_19597_, _19596_, _19585_);
  or _42413_ (_19598_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _42414_ (_19599_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and _42415_ (_19600_, _19599_, _19598_);
  and _42416_ (_19601_, _19600_, _05996_);
  or _42417_ (_19602_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _42418_ (_19603_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and _42419_ (_19604_, _19603_, _19602_);
  and _42420_ (_19605_, _19604_, _05997_);
  or _42421_ (_19606_, _19605_, _19601_);
  or _42422_ (_19607_, _19606_, _06021_);
  or _42423_ (_19608_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _42424_ (_19609_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and _42425_ (_19610_, _19609_, _19608_);
  and _42426_ (_19611_, _19610_, _05996_);
  or _42427_ (_19612_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _42428_ (_19613_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and _42429_ (_19614_, _19613_, _19612_);
  and _42430_ (_19615_, _19614_, _05997_);
  or _42431_ (_19616_, _19615_, _19611_);
  or _42432_ (_19617_, _19616_, _05920_);
  and _42433_ (_19618_, _19617_, _05933_);
  and _42434_ (_19619_, _19618_, _19607_);
  or _42435_ (_19620_, _19619_, _19597_);
  and _42436_ (_19621_, _19620_, _05776_);
  or _42437_ (_19622_, _19621_, _19575_);
  and _42438_ (_19623_, _19622_, _06070_);
  or _42439_ (_19624_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _42440_ (_19625_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and _42441_ (_19626_, _19625_, _19624_);
  and _42442_ (_19627_, _19626_, _05996_);
  or _42443_ (_19628_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _42444_ (_19629_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and _42445_ (_19630_, _19629_, _19628_);
  and _42446_ (_19631_, _19630_, _05997_);
  or _42447_ (_19632_, _19631_, _19627_);
  and _42448_ (_19633_, _19632_, _06021_);
  or _42449_ (_19634_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _42450_ (_19635_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and _42451_ (_19636_, _19635_, _19634_);
  and _42452_ (_19637_, _19636_, _05996_);
  or _42453_ (_19638_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _42454_ (_19639_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and _42455_ (_19640_, _19639_, _19638_);
  and _42456_ (_19641_, _19640_, _05997_);
  or _42457_ (_19642_, _19641_, _19637_);
  and _42458_ (_19643_, _19642_, _05920_);
  or _42459_ (_19644_, _19643_, _19633_);
  and _42460_ (_19645_, _19644_, _05933_);
  and _42461_ (_19646_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and _42462_ (_19647_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _42463_ (_19648_, _19647_, _19646_);
  and _42464_ (_19649_, _19648_, _05996_);
  and _42465_ (_19650_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and _42466_ (_19651_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _42467_ (_19652_, _19651_, _19650_);
  and _42468_ (_19653_, _19652_, _05997_);
  or _42469_ (_19654_, _19653_, _19649_);
  and _42470_ (_19655_, _19654_, _06021_);
  and _42471_ (_19656_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and _42472_ (_19657_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _42473_ (_19658_, _19657_, _19656_);
  and _42474_ (_19659_, _19658_, _05996_);
  and _42475_ (_19660_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and _42476_ (_19661_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _42477_ (_19662_, _19661_, _19660_);
  and _42478_ (_19663_, _19662_, _05997_);
  or _42479_ (_19664_, _19663_, _19659_);
  and _42480_ (_19665_, _19664_, _05920_);
  or _42481_ (_19666_, _19665_, _19655_);
  and _42482_ (_19667_, _19666_, _06033_);
  or _42483_ (_19668_, _19667_, _19645_);
  and _42484_ (_19669_, _19668_, _05776_);
  or _42485_ (_19670_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _42486_ (_19671_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and _42487_ (_19672_, _19671_, _05997_);
  and _42488_ (_19673_, _19672_, _19670_);
  or _42489_ (_19674_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or _42490_ (_19675_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and _42491_ (_19676_, _19675_, _05996_);
  and _42492_ (_19677_, _19676_, _19674_);
  or _42493_ (_19678_, _19677_, _19673_);
  and _42494_ (_19679_, _19678_, _06021_);
  or _42495_ (_19680_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _42496_ (_19681_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and _42497_ (_19682_, _19681_, _05997_);
  and _42498_ (_19683_, _19682_, _19680_);
  or _42499_ (_19684_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or _42500_ (_19685_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and _42501_ (_19686_, _19685_, _05996_);
  and _42502_ (_19687_, _19686_, _19684_);
  or _42503_ (_19688_, _19687_, _19683_);
  and _42504_ (_19689_, _19688_, _05920_);
  or _42505_ (_19690_, _19689_, _19679_);
  and _42506_ (_19691_, _19690_, _05933_);
  and _42507_ (_19692_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and _42508_ (_19693_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or _42509_ (_19694_, _19693_, _19692_);
  and _42510_ (_19695_, _19694_, _05996_);
  and _42511_ (_19696_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and _42512_ (_19697_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or _42513_ (_19698_, _19697_, _19696_);
  and _42514_ (_19699_, _19698_, _05997_);
  or _42515_ (_19700_, _19699_, _19695_);
  and _42516_ (_19701_, _19700_, _06021_);
  and _42517_ (_19702_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and _42518_ (_19703_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or _42519_ (_19704_, _19703_, _19702_);
  and _42520_ (_19705_, _19704_, _05996_);
  and _42521_ (_19706_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and _42522_ (_19707_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _42523_ (_19708_, _19707_, _19706_);
  and _42524_ (_19709_, _19708_, _05997_);
  or _42525_ (_19710_, _19709_, _19705_);
  and _42526_ (_19711_, _19710_, _05920_);
  or _42527_ (_19712_, _19711_, _19701_);
  and _42528_ (_19713_, _19712_, _06033_);
  or _42529_ (_19714_, _19713_, _19691_);
  and _42530_ (_19715_, _19714_, _06071_);
  or _42531_ (_19716_, _19715_, _19669_);
  and _42532_ (_19717_, _19716_, _05822_);
  or _42533_ (_19718_, _19717_, _19623_);
  or _42534_ (_19719_, _19718_, _06616_);
  and _42535_ (_19720_, _19719_, _19529_);
  or _42536_ (_19721_, _19720_, _06020_);
  and _42537_ (_19722_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and _42538_ (_19723_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _42539_ (_19724_, _19723_, _19722_);
  and _42540_ (_19725_, _19724_, _05996_);
  and _42541_ (_19726_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and _42542_ (_19727_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _42543_ (_19728_, _19727_, _19726_);
  and _42544_ (_19729_, _19728_, _05997_);
  or _42545_ (_19730_, _19729_, _19725_);
  or _42546_ (_19731_, _19730_, _06021_);
  and _42547_ (_19732_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and _42548_ (_19733_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _42549_ (_19734_, _19733_, _19732_);
  and _42550_ (_19735_, _19734_, _05996_);
  and _42551_ (_19736_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and _42552_ (_19737_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _42553_ (_19738_, _19737_, _19736_);
  and _42554_ (_19739_, _19738_, _05997_);
  or _42555_ (_19740_, _19739_, _19735_);
  or _42556_ (_19741_, _19740_, _05920_);
  and _42557_ (_19742_, _19741_, _06033_);
  and _42558_ (_19743_, _19742_, _19731_);
  or _42559_ (_19744_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _42560_ (_19745_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and _42561_ (_19746_, _19745_, _19744_);
  and _42562_ (_19747_, _19746_, _05996_);
  or _42563_ (_19748_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _42564_ (_19749_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and _42565_ (_19750_, _19749_, _19748_);
  and _42566_ (_19751_, _19750_, _05997_);
  or _42567_ (_19752_, _19751_, _19747_);
  or _42568_ (_19753_, _19752_, _06021_);
  or _42569_ (_19754_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _42570_ (_19755_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and _42571_ (_19756_, _19755_, _19754_);
  and _42572_ (_19757_, _19756_, _05996_);
  or _42573_ (_19758_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _42574_ (_19759_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and _42575_ (_19760_, _19759_, _19758_);
  and _42576_ (_19761_, _19760_, _05997_);
  or _42577_ (_19762_, _19761_, _19757_);
  or _42578_ (_19763_, _19762_, _05920_);
  and _42579_ (_19764_, _19763_, _05933_);
  and _42580_ (_19765_, _19764_, _19753_);
  or _42581_ (_19766_, _19765_, _19743_);
  and _42582_ (_19767_, _19766_, _05776_);
  and _42583_ (_19768_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _42584_ (_19769_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or _42585_ (_19770_, _19769_, _19768_);
  and _42586_ (_19771_, _19770_, _05996_);
  and _42587_ (_19772_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _42588_ (_19773_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or _42589_ (_19774_, _19773_, _19772_);
  and _42590_ (_19775_, _19774_, _05997_);
  or _42591_ (_19776_, _19775_, _19771_);
  or _42592_ (_19777_, _19776_, _06021_);
  and _42593_ (_19778_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _42594_ (_19779_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _42595_ (_19780_, _19779_, _19778_);
  and _42596_ (_19781_, _19780_, _05996_);
  and _42597_ (_19782_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _42598_ (_19783_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or _42599_ (_19784_, _19783_, _19782_);
  and _42600_ (_19785_, _19784_, _05997_);
  or _42601_ (_19786_, _19785_, _19781_);
  or _42602_ (_19787_, _19786_, _05920_);
  and _42603_ (_19788_, _19787_, _06033_);
  and _42604_ (_19789_, _19788_, _19777_);
  or _42605_ (_19790_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or _42606_ (_19791_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _42607_ (_19792_, _19791_, _05997_);
  and _42608_ (_19793_, _19792_, _19790_);
  or _42609_ (_19794_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _42610_ (_19795_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and _42611_ (_19796_, _19795_, _05996_);
  and _42612_ (_19797_, _19796_, _19794_);
  or _42613_ (_19798_, _19797_, _19793_);
  or _42614_ (_19799_, _19798_, _06021_);
  or _42615_ (_19800_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or _42616_ (_19801_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _42617_ (_19802_, _19801_, _05997_);
  and _42618_ (_19803_, _19802_, _19800_);
  or _42619_ (_19804_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _42620_ (_19805_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _42621_ (_19806_, _19805_, _05996_);
  and _42622_ (_19807_, _19806_, _19804_);
  or _42623_ (_19808_, _19807_, _19803_);
  or _42624_ (_19809_, _19808_, _05920_);
  and _42625_ (_19810_, _19809_, _05933_);
  and _42626_ (_19811_, _19810_, _19799_);
  or _42627_ (_19812_, _19811_, _19789_);
  and _42628_ (_19813_, _19812_, _06071_);
  or _42629_ (_19814_, _19813_, _19767_);
  and _42630_ (_19815_, _19814_, _06070_);
  and _42631_ (_19816_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and _42632_ (_19817_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or _42633_ (_19818_, _19817_, _19816_);
  and _42634_ (_19819_, _19818_, _05996_);
  and _42635_ (_19820_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and _42636_ (_19821_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or _42637_ (_19822_, _19821_, _19820_);
  and _42638_ (_19823_, _19822_, _05997_);
  or _42639_ (_19824_, _19823_, _19819_);
  and _42640_ (_19825_, _19824_, _05920_);
  and _42641_ (_19826_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and _42642_ (_19827_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or _42643_ (_19828_, _19827_, _19826_);
  and _42644_ (_19829_, _19828_, _05996_);
  and _42645_ (_19830_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _42646_ (_19831_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or _42647_ (_19832_, _19831_, _19830_);
  and _42648_ (_19833_, _19832_, _05997_);
  or _42649_ (_19834_, _19833_, _19829_);
  and _42650_ (_19835_, _19834_, _06021_);
  or _42651_ (_19836_, _19835_, _19825_);
  and _42652_ (_19837_, _19836_, _06033_);
  or _42653_ (_19838_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or _42654_ (_19839_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and _42655_ (_19840_, _19839_, _05997_);
  and _42656_ (_19841_, _19840_, _19838_);
  or _42657_ (_19842_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or _42658_ (_19843_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and _42659_ (_19844_, _19843_, _05996_);
  and _42660_ (_19845_, _19844_, _19842_);
  or _42661_ (_19846_, _19845_, _19841_);
  and _42662_ (_19847_, _19846_, _05920_);
  or _42663_ (_19848_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or _42664_ (_19849_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and _42665_ (_19850_, _19849_, _05997_);
  and _42666_ (_19851_, _19850_, _19848_);
  or _42667_ (_19852_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or _42668_ (_19853_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and _42669_ (_19854_, _19853_, _05996_);
  and _42670_ (_19855_, _19854_, _19852_);
  or _42671_ (_19856_, _19855_, _19851_);
  and _42672_ (_19857_, _19856_, _06021_);
  or _42673_ (_19858_, _19857_, _19847_);
  and _42674_ (_19859_, _19858_, _05933_);
  or _42675_ (_19860_, _19859_, _19837_);
  and _42676_ (_19861_, _19860_, _06071_);
  and _42677_ (_19862_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _42678_ (_19863_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _42679_ (_19864_, _19863_, _19862_);
  and _42680_ (_19865_, _19864_, _05996_);
  and _42681_ (_19866_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and _42682_ (_19867_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _42683_ (_19868_, _19867_, _19866_);
  and _42684_ (_19869_, _19868_, _05997_);
  or _42685_ (_19870_, _19869_, _19865_);
  and _42686_ (_19871_, _19870_, _05920_);
  and _42687_ (_19872_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _42688_ (_19873_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _42689_ (_19874_, _19873_, _19872_);
  and _42690_ (_19875_, _19874_, _05996_);
  and _42691_ (_19876_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and _42692_ (_19877_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _42693_ (_19878_, _19877_, _19876_);
  and _42694_ (_19879_, _19878_, _05997_);
  or _42695_ (_19880_, _19879_, _19875_);
  and _42696_ (_19881_, _19880_, _06021_);
  or _42697_ (_19882_, _19881_, _19871_);
  and _42698_ (_19883_, _19882_, _06033_);
  or _42699_ (_19884_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _42700_ (_19885_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and _42701_ (_19886_, _19885_, _19884_);
  and _42702_ (_19887_, _19886_, _05996_);
  or _42703_ (_19888_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _42704_ (_19889_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _42705_ (_19890_, _19889_, _19888_);
  and _42706_ (_19891_, _19890_, _05997_);
  or _42707_ (_19892_, _19891_, _19887_);
  and _42708_ (_19893_, _19892_, _05920_);
  or _42709_ (_19894_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _42710_ (_19895_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and _42711_ (_19896_, _19895_, _19894_);
  and _42712_ (_19897_, _19896_, _05996_);
  or _42713_ (_19898_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _42714_ (_19899_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _42715_ (_19900_, _19899_, _19898_);
  and _42716_ (_19901_, _19900_, _05997_);
  or _42717_ (_19902_, _19901_, _19897_);
  and _42718_ (_19903_, _19902_, _06021_);
  or _42719_ (_19904_, _19903_, _19893_);
  and _42720_ (_19905_, _19904_, _05933_);
  or _42721_ (_19906_, _19905_, _19883_);
  and _42722_ (_19907_, _19906_, _05776_);
  or _42723_ (_19909_, _19907_, _19861_);
  and _42724_ (_19910_, _19909_, _05822_);
  or _42725_ (_19911_, _19910_, _19815_);
  or _42726_ (_19912_, _19911_, _05868_);
  and _42727_ (_19913_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and _42728_ (_19914_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _42729_ (_19915_, _19914_, _19913_);
  and _42730_ (_19916_, _19915_, _05996_);
  and _42731_ (_19917_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and _42732_ (_19918_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _42733_ (_19920_, _19918_, _19917_);
  and _42734_ (_19921_, _19920_, _05997_);
  or _42735_ (_19922_, _19921_, _19916_);
  or _42736_ (_19923_, _19922_, _06021_);
  and _42737_ (_19924_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and _42738_ (_19925_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _42739_ (_19926_, _19925_, _19924_);
  and _42740_ (_19927_, _19926_, _05996_);
  and _42741_ (_19928_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and _42742_ (_19929_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _42743_ (_19931_, _19929_, _19928_);
  and _42744_ (_19932_, _19931_, _05997_);
  or _42745_ (_19933_, _19932_, _19927_);
  or _42746_ (_19934_, _19933_, _05920_);
  and _42747_ (_19935_, _19934_, _06033_);
  and _42748_ (_19936_, _19935_, _19923_);
  or _42749_ (_19937_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _42750_ (_19938_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and _42751_ (_19939_, _19938_, _05997_);
  and _42752_ (_19940_, _19939_, _19937_);
  or _42753_ (_19942_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _42754_ (_19943_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and _42755_ (_19944_, _19943_, _05996_);
  and _42756_ (_19945_, _19944_, _19942_);
  or _42757_ (_19946_, _19945_, _19940_);
  or _42758_ (_19947_, _19946_, _06021_);
  or _42759_ (_19948_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _42760_ (_19949_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and _42761_ (_19950_, _19949_, _05997_);
  and _42762_ (_19951_, _19950_, _19948_);
  or _42763_ (_19953_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _42764_ (_19954_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and _42765_ (_19955_, _19954_, _05996_);
  and _42766_ (_19956_, _19955_, _19953_);
  or _42767_ (_19957_, _19956_, _19951_);
  or _42768_ (_19958_, _19957_, _05920_);
  and _42769_ (_19959_, _19958_, _05933_);
  and _42770_ (_19960_, _19959_, _19947_);
  or _42771_ (_19961_, _19960_, _19936_);
  and _42772_ (_19962_, _19961_, _06071_);
  and _42773_ (_19964_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _42774_ (_19965_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _42775_ (_19966_, _19965_, _19964_);
  and _42776_ (_19967_, _19966_, _05996_);
  and _42777_ (_19968_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _42778_ (_19969_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or _42779_ (_19970_, _19969_, _19968_);
  and _42780_ (_19971_, _19970_, _05997_);
  or _42781_ (_19972_, _19971_, _19967_);
  or _42782_ (_19973_, _19972_, _06021_);
  and _42783_ (_19974_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _42784_ (_19975_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or _42785_ (_19976_, _19975_, _19974_);
  and _42786_ (_19977_, _19976_, _05996_);
  and _42787_ (_19978_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _42788_ (_19979_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _42789_ (_19980_, _19979_, _19978_);
  and _42790_ (_19981_, _19980_, _05997_);
  or _42791_ (_19982_, _19981_, _19977_);
  or _42792_ (_19983_, _19982_, _05920_);
  and _42793_ (_19984_, _19983_, _06033_);
  and _42794_ (_19985_, _19984_, _19973_);
  or _42795_ (_19986_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or _42796_ (_19987_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _42797_ (_19988_, _19987_, _19986_);
  and _42798_ (_19989_, _19988_, _05996_);
  or _42799_ (_19990_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or _42800_ (_19991_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and _42801_ (_19992_, _19991_, _19990_);
  and _42802_ (_19993_, _19992_, _05997_);
  or _42803_ (_19994_, _19993_, _19989_);
  or _42804_ (_19995_, _19994_, _06021_);
  or _42805_ (_19996_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _42806_ (_19997_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _42807_ (_19998_, _19997_, _19996_);
  and _42808_ (_19999_, _19998_, _05996_);
  or _42809_ (_20000_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _42810_ (_20001_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and _42811_ (_20002_, _20001_, _20000_);
  and _42812_ (_20003_, _20002_, _05997_);
  or _42813_ (_20004_, _20003_, _19999_);
  or _42814_ (_20005_, _20004_, _05920_);
  and _42815_ (_20006_, _20005_, _05933_);
  and _42816_ (_20007_, _20006_, _19995_);
  or _42817_ (_20008_, _20007_, _19985_);
  and _42818_ (_20009_, _20008_, _05776_);
  or _42819_ (_20010_, _20009_, _19962_);
  and _42820_ (_20011_, _20010_, _06070_);
  or _42821_ (_20012_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _42822_ (_20013_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _42823_ (_20014_, _20013_, _20012_);
  and _42824_ (_20015_, _20014_, _05996_);
  or _42825_ (_20016_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _42826_ (_20017_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and _42827_ (_20018_, _20017_, _20016_);
  and _42828_ (_20019_, _20018_, _05997_);
  or _42829_ (_20020_, _20019_, _20015_);
  and _42830_ (_20021_, _20020_, _06021_);
  or _42831_ (_20022_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or _42832_ (_20023_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and _42833_ (_20024_, _20023_, _20022_);
  and _42834_ (_20025_, _20024_, _05996_);
  or _42835_ (_20026_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or _42836_ (_20027_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _42837_ (_20028_, _20027_, _20026_);
  and _42838_ (_20029_, _20028_, _05997_);
  or _42839_ (_20030_, _20029_, _20025_);
  and _42840_ (_20031_, _20030_, _05920_);
  or _42841_ (_20032_, _20031_, _20021_);
  and _42842_ (_20033_, _20032_, _05933_);
  and _42843_ (_20034_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _42844_ (_20035_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or _42845_ (_20036_, _20035_, _20034_);
  and _42846_ (_20037_, _20036_, _05996_);
  and _42847_ (_20038_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _42848_ (_20039_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _42849_ (_20040_, _20039_, _20038_);
  and _42850_ (_20041_, _20040_, _05997_);
  or _42851_ (_20042_, _20041_, _20037_);
  and _42852_ (_20043_, _20042_, _06021_);
  and _42853_ (_20044_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _42854_ (_20045_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or _42855_ (_20046_, _20045_, _20044_);
  and _42856_ (_20047_, _20046_, _05996_);
  and _42857_ (_20048_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and _42858_ (_20049_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _42859_ (_20050_, _20049_, _20048_);
  and _42860_ (_20051_, _20050_, _05997_);
  or _42861_ (_20052_, _20051_, _20047_);
  and _42862_ (_20053_, _20052_, _05920_);
  or _42863_ (_20054_, _20053_, _20043_);
  and _42864_ (_20055_, _20054_, _06033_);
  or _42865_ (_20056_, _20055_, _20033_);
  and _42866_ (_20057_, _20056_, _05776_);
  or _42867_ (_20058_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _42868_ (_20059_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and _42869_ (_20060_, _20059_, _05997_);
  and _42870_ (_20061_, _20060_, _20058_);
  or _42871_ (_20062_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _42872_ (_20063_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and _42873_ (_20064_, _20063_, _05996_);
  and _42874_ (_20065_, _20064_, _20062_);
  or _42875_ (_20066_, _20065_, _20061_);
  and _42876_ (_20067_, _20066_, _06021_);
  or _42877_ (_20068_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _42878_ (_20069_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _42879_ (_20070_, _20069_, _05997_);
  and _42880_ (_20071_, _20070_, _20068_);
  or _42881_ (_20072_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _42882_ (_20073_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and _42883_ (_20074_, _20073_, _05996_);
  and _42884_ (_20075_, _20074_, _20072_);
  or _42885_ (_20076_, _20075_, _20071_);
  and _42886_ (_20077_, _20076_, _05920_);
  or _42887_ (_20078_, _20077_, _20067_);
  and _42888_ (_20079_, _20078_, _05933_);
  and _42889_ (_20080_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _42890_ (_20081_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _42891_ (_20082_, _20081_, _20080_);
  and _42892_ (_20083_, _20082_, _05996_);
  and _42893_ (_20084_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and _42894_ (_20085_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _42895_ (_20086_, _20085_, _20084_);
  and _42896_ (_20087_, _20086_, _05997_);
  or _42897_ (_20088_, _20087_, _20083_);
  and _42898_ (_20089_, _20088_, _06021_);
  and _42899_ (_20090_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and _42900_ (_20091_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _42901_ (_20092_, _20091_, _20090_);
  and _42902_ (_20093_, _20092_, _05996_);
  and _42903_ (_20094_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and _42904_ (_20095_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _42905_ (_20096_, _20095_, _20094_);
  and _42906_ (_20097_, _20096_, _05997_);
  or _42907_ (_20098_, _20097_, _20093_);
  and _42908_ (_20099_, _20098_, _05920_);
  or _42909_ (_20100_, _20099_, _20089_);
  and _42910_ (_20101_, _20100_, _06033_);
  or _42911_ (_20102_, _20101_, _20079_);
  and _42912_ (_20103_, _20102_, _06071_);
  or _42913_ (_20104_, _20103_, _20057_);
  and _42914_ (_20105_, _20104_, _05822_);
  or _42915_ (_20106_, _20105_, _20011_);
  or _42916_ (_20107_, _20106_, _06616_);
  and _42917_ (_20108_, _20107_, _19912_);
  or _42918_ (_20109_, _20108_, _05584_);
  and _42919_ (_20110_, _20109_, _19721_);
  or _42920_ (_20111_, _20110_, _06019_);
  or _42921_ (_20112_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and _42922_ (_20113_, _20112_, _25365_);
  and _42923_ (_14807_, _20113_, _20111_);
  and _42924_ (_20114_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and _42925_ (_20115_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _42926_ (_20116_, _20115_, _20114_);
  and _42927_ (_20117_, _20116_, _05996_);
  and _42928_ (_20118_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and _42929_ (_20119_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _42930_ (_20120_, _20119_, _20118_);
  and _42931_ (_20121_, _20120_, _05997_);
  or _42932_ (_20122_, _20121_, _20117_);
  or _42933_ (_20123_, _20122_, _06021_);
  and _42934_ (_20124_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and _42935_ (_20125_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _42936_ (_20126_, _20125_, _20124_);
  and _42937_ (_20127_, _20126_, _05996_);
  and _42938_ (_20128_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and _42939_ (_20129_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _42940_ (_20130_, _20129_, _20128_);
  and _42941_ (_20131_, _20130_, _05997_);
  or _42942_ (_20132_, _20131_, _20127_);
  or _42943_ (_20133_, _20132_, _05920_);
  and _42944_ (_20134_, _20133_, _06033_);
  and _42945_ (_20135_, _20134_, _20123_);
  or _42946_ (_20136_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _42947_ (_20137_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and _42948_ (_20138_, _20137_, _20136_);
  and _42949_ (_20139_, _20138_, _05996_);
  or _42950_ (_20140_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _42951_ (_20141_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and _42952_ (_20142_, _20141_, _20140_);
  and _42953_ (_20143_, _20142_, _05997_);
  or _42954_ (_20144_, _20143_, _20139_);
  or _42955_ (_20145_, _20144_, _06021_);
  or _42956_ (_20146_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _42957_ (_20147_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and _42958_ (_20148_, _20147_, _20146_);
  and _42959_ (_20149_, _20148_, _05996_);
  or _42960_ (_20150_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _42961_ (_20151_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and _42962_ (_20152_, _20151_, _20150_);
  and _42963_ (_20153_, _20152_, _05997_);
  or _42964_ (_20154_, _20153_, _20149_);
  or _42965_ (_20155_, _20154_, _05920_);
  and _42966_ (_20156_, _20155_, _05933_);
  and _42967_ (_20157_, _20156_, _20145_);
  or _42968_ (_20158_, _20157_, _20135_);
  and _42969_ (_20159_, _20158_, _05776_);
  and _42970_ (_20160_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and _42971_ (_20161_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _42972_ (_20162_, _20161_, _20160_);
  and _42973_ (_20163_, _20162_, _05996_);
  and _42974_ (_20164_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and _42975_ (_20165_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _42976_ (_20166_, _20165_, _20164_);
  and _42977_ (_20167_, _20166_, _05997_);
  or _42978_ (_20168_, _20167_, _20163_);
  or _42979_ (_20169_, _20168_, _06021_);
  and _42980_ (_20170_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and _42981_ (_20171_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _42982_ (_20172_, _20171_, _20170_);
  and _42983_ (_20173_, _20172_, _05996_);
  and _42984_ (_20174_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and _42985_ (_20175_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _42986_ (_20176_, _20175_, _20174_);
  and _42987_ (_20177_, _20176_, _05997_);
  or _42988_ (_20178_, _20177_, _20173_);
  or _42989_ (_20179_, _20178_, _05920_);
  and _42990_ (_20180_, _20179_, _06033_);
  and _42991_ (_20181_, _20180_, _20169_);
  or _42992_ (_20182_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _42993_ (_20183_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and _42994_ (_20184_, _20183_, _05997_);
  and _42995_ (_20185_, _20184_, _20182_);
  or _42996_ (_20186_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _42997_ (_20187_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and _42998_ (_20188_, _20187_, _05996_);
  and _42999_ (_20189_, _20188_, _20186_);
  or _43000_ (_20190_, _20189_, _20185_);
  or _43001_ (_20191_, _20190_, _06021_);
  or _43002_ (_20192_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _43003_ (_20193_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and _43004_ (_20194_, _20193_, _05997_);
  and _43005_ (_20195_, _20194_, _20192_);
  or _43006_ (_20196_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _43007_ (_20197_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and _43008_ (_20198_, _20197_, _05996_);
  and _43009_ (_20199_, _20198_, _20196_);
  or _43010_ (_20200_, _20199_, _20195_);
  or _43011_ (_20201_, _20200_, _05920_);
  and _43012_ (_20202_, _20201_, _05933_);
  and _43013_ (_20203_, _20202_, _20191_);
  or _43014_ (_20204_, _20203_, _20181_);
  and _43015_ (_20205_, _20204_, _06071_);
  or _43016_ (_20206_, _20205_, _20159_);
  and _43017_ (_20207_, _20206_, _06070_);
  and _43018_ (_20208_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and _43019_ (_20209_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _43020_ (_20210_, _20209_, _20208_);
  and _43021_ (_20211_, _20210_, _05996_);
  and _43022_ (_20212_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _43023_ (_20213_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _43024_ (_20214_, _20213_, _20212_);
  and _43025_ (_20215_, _20214_, _05997_);
  or _43026_ (_20216_, _20215_, _20211_);
  and _43027_ (_20217_, _20216_, _05920_);
  and _43028_ (_20218_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _43029_ (_20219_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _43030_ (_20220_, _20219_, _20218_);
  and _43031_ (_20221_, _20220_, _05996_);
  and _43032_ (_20222_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and _43033_ (_20223_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _43034_ (_20224_, _20223_, _20222_);
  and _43035_ (_20225_, _20224_, _05997_);
  or _43036_ (_20226_, _20225_, _20221_);
  and _43037_ (_20227_, _20226_, _06021_);
  or _43038_ (_20228_, _20227_, _20217_);
  and _43039_ (_20229_, _20228_, _06033_);
  or _43040_ (_20230_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _43041_ (_20231_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _43042_ (_20232_, _20231_, _05997_);
  and _43043_ (_20233_, _20232_, _20230_);
  or _43044_ (_20234_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _43045_ (_20235_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _43046_ (_20236_, _20235_, _05996_);
  and _43047_ (_20237_, _20236_, _20234_);
  or _43048_ (_20238_, _20237_, _20233_);
  and _43049_ (_20239_, _20238_, _05920_);
  or _43050_ (_20240_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _43051_ (_20241_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _43052_ (_20242_, _20241_, _05997_);
  and _43053_ (_20243_, _20242_, _20240_);
  or _43054_ (_20244_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _43055_ (_20245_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _43056_ (_20246_, _20245_, _05996_);
  and _43057_ (_20247_, _20246_, _20244_);
  or _43058_ (_20248_, _20247_, _20243_);
  and _43059_ (_20249_, _20248_, _06021_);
  or _43060_ (_20250_, _20249_, _20239_);
  and _43061_ (_20251_, _20250_, _05933_);
  or _43062_ (_20252_, _20251_, _20229_);
  and _43063_ (_20253_, _20252_, _06071_);
  and _43064_ (_20254_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and _43065_ (_20255_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _43066_ (_20256_, _20255_, _20254_);
  and _43067_ (_20257_, _20256_, _05996_);
  and _43068_ (_20258_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and _43069_ (_20259_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _43070_ (_20260_, _20259_, _20258_);
  and _43071_ (_20261_, _20260_, _05997_);
  or _43072_ (_20262_, _20261_, _20257_);
  and _43073_ (_20263_, _20262_, _05920_);
  and _43074_ (_20264_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and _43075_ (_20265_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _43076_ (_20266_, _20265_, _20264_);
  and _43077_ (_20267_, _20266_, _05996_);
  and _43078_ (_20268_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and _43079_ (_20269_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _43080_ (_20270_, _20269_, _20268_);
  and _43081_ (_20271_, _20270_, _05997_);
  or _43082_ (_20272_, _20271_, _20267_);
  and _43083_ (_20273_, _20272_, _06021_);
  or _43084_ (_20274_, _20273_, _20263_);
  and _43085_ (_20275_, _20274_, _06033_);
  or _43086_ (_20276_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _43087_ (_20277_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and _43088_ (_20278_, _20277_, _20276_);
  and _43089_ (_20279_, _20278_, _05996_);
  or _43090_ (_20280_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _43091_ (_20281_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and _43092_ (_20282_, _20281_, _20280_);
  and _43093_ (_20283_, _20282_, _05997_);
  or _43094_ (_20284_, _20283_, _20279_);
  and _43095_ (_20285_, _20284_, _05920_);
  or _43096_ (_20286_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _43097_ (_20287_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and _43098_ (_20288_, _20287_, _20286_);
  and _43099_ (_20289_, _20288_, _05996_);
  or _43100_ (_20290_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _43101_ (_20291_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and _43102_ (_20292_, _20291_, _20290_);
  and _43103_ (_20293_, _20292_, _05997_);
  or _43104_ (_20294_, _20293_, _20289_);
  and _43105_ (_20295_, _20294_, _06021_);
  or _43106_ (_20296_, _20295_, _20285_);
  and _43107_ (_20297_, _20296_, _05933_);
  or _43108_ (_20298_, _20297_, _20275_);
  and _43109_ (_20299_, _20298_, _05776_);
  or _43110_ (_20300_, _20299_, _20253_);
  and _43111_ (_20301_, _20300_, _05822_);
  or _43112_ (_20302_, _20301_, _20207_);
  or _43113_ (_20303_, _20302_, _05868_);
  and _43114_ (_20304_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and _43115_ (_20305_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _43116_ (_20306_, _20305_, _20304_);
  and _43117_ (_20307_, _20306_, _05996_);
  and _43118_ (_20308_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and _43119_ (_20309_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _43120_ (_20310_, _20309_, _20308_);
  and _43121_ (_20311_, _20310_, _05997_);
  or _43122_ (_20312_, _20311_, _20307_);
  or _43123_ (_20313_, _20312_, _06021_);
  and _43124_ (_20314_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and _43125_ (_20315_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _43126_ (_20316_, _20315_, _20314_);
  and _43127_ (_20317_, _20316_, _05996_);
  and _43128_ (_20318_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and _43129_ (_20319_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _43130_ (_20320_, _20319_, _20318_);
  and _43131_ (_20321_, _20320_, _05997_);
  or _43132_ (_20322_, _20321_, _20317_);
  or _43133_ (_20323_, _20322_, _05920_);
  and _43134_ (_20324_, _20323_, _06033_);
  and _43135_ (_20325_, _20324_, _20313_);
  or _43136_ (_20326_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _43137_ (_20327_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and _43138_ (_20328_, _20327_, _05997_);
  and _43139_ (_20329_, _20328_, _20326_);
  or _43140_ (_20330_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _43141_ (_20331_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and _43142_ (_20332_, _20331_, _05996_);
  and _43143_ (_20333_, _20332_, _20330_);
  or _43144_ (_20334_, _20333_, _20329_);
  or _43145_ (_20335_, _20334_, _06021_);
  or _43146_ (_20336_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _43147_ (_20337_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and _43148_ (_20338_, _20337_, _05997_);
  and _43149_ (_20339_, _20338_, _20336_);
  or _43150_ (_20340_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _43151_ (_20341_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and _43152_ (_20342_, _20341_, _05996_);
  and _43153_ (_20343_, _20342_, _20340_);
  or _43154_ (_20344_, _20343_, _20339_);
  or _43155_ (_20345_, _20344_, _05920_);
  and _43156_ (_20346_, _20345_, _05933_);
  and _43157_ (_20347_, _20346_, _20335_);
  or _43158_ (_20348_, _20347_, _20325_);
  and _43159_ (_20349_, _20348_, _06071_);
  and _43160_ (_20350_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _43161_ (_20351_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _43162_ (_20352_, _20351_, _20350_);
  and _43163_ (_20353_, _20352_, _05996_);
  and _43164_ (_20354_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and _43165_ (_20355_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _43166_ (_20356_, _20355_, _20354_);
  and _43167_ (_20357_, _20356_, _05997_);
  or _43168_ (_20358_, _20357_, _20353_);
  or _43169_ (_20359_, _20358_, _06021_);
  and _43170_ (_20360_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and _43171_ (_20361_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _43172_ (_20362_, _20361_, _20360_);
  and _43173_ (_20363_, _20362_, _05996_);
  and _43174_ (_20364_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and _43175_ (_20365_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _43176_ (_20366_, _20365_, _20364_);
  and _43177_ (_20367_, _20366_, _05997_);
  or _43178_ (_20368_, _20367_, _20363_);
  or _43179_ (_20369_, _20368_, _05920_);
  and _43180_ (_20370_, _20369_, _06033_);
  and _43181_ (_20371_, _20370_, _20359_);
  or _43182_ (_20372_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _43183_ (_20373_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and _43184_ (_20374_, _20373_, _20372_);
  and _43185_ (_20375_, _20374_, _05996_);
  or _43186_ (_20376_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _43187_ (_20377_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and _43188_ (_20378_, _20377_, _20376_);
  and _43189_ (_20379_, _20378_, _05997_);
  or _43190_ (_20380_, _20379_, _20375_);
  or _43191_ (_20381_, _20380_, _06021_);
  or _43192_ (_20382_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _43193_ (_20383_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and _43194_ (_20384_, _20383_, _20382_);
  and _43195_ (_20385_, _20384_, _05996_);
  or _43196_ (_20386_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _43197_ (_20387_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and _43198_ (_20388_, _20387_, _20386_);
  and _43199_ (_20389_, _20388_, _05997_);
  or _43200_ (_20390_, _20389_, _20385_);
  or _43201_ (_20391_, _20390_, _05920_);
  and _43202_ (_20392_, _20391_, _05933_);
  and _43203_ (_20393_, _20392_, _20381_);
  or _43204_ (_20394_, _20393_, _20371_);
  and _43205_ (_20395_, _20394_, _05776_);
  or _43206_ (_20396_, _20395_, _20349_);
  and _43207_ (_20397_, _20396_, _06070_);
  or _43208_ (_20398_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _43209_ (_20399_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and _43210_ (_20400_, _20399_, _20398_);
  and _43211_ (_20401_, _20400_, _05996_);
  or _43212_ (_20402_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _43213_ (_20403_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and _43214_ (_20404_, _20403_, _20402_);
  and _43215_ (_20405_, _20404_, _05997_);
  or _43216_ (_20406_, _20405_, _20401_);
  and _43217_ (_20407_, _20406_, _06021_);
  or _43218_ (_20408_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _43219_ (_20409_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and _43220_ (_20410_, _20409_, _20408_);
  and _43221_ (_20411_, _20410_, _05996_);
  or _43222_ (_20412_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _43223_ (_20413_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and _43224_ (_20414_, _20413_, _20412_);
  and _43225_ (_20415_, _20414_, _05997_);
  or _43226_ (_20416_, _20415_, _20411_);
  and _43227_ (_20417_, _20416_, _05920_);
  or _43228_ (_20418_, _20417_, _20407_);
  and _43229_ (_20419_, _20418_, _05933_);
  and _43230_ (_20420_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and _43231_ (_20421_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _43232_ (_20422_, _20421_, _20420_);
  and _43233_ (_20423_, _20422_, _05996_);
  and _43234_ (_20424_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and _43235_ (_20425_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _43236_ (_20426_, _20425_, _20424_);
  and _43237_ (_20427_, _20426_, _05997_);
  or _43238_ (_20428_, _20427_, _20423_);
  and _43239_ (_20429_, _20428_, _06021_);
  and _43240_ (_20430_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and _43241_ (_20431_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _43242_ (_20432_, _20431_, _20430_);
  and _43243_ (_20433_, _20432_, _05996_);
  and _43244_ (_20434_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and _43245_ (_20435_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _43246_ (_20436_, _20435_, _20434_);
  and _43247_ (_20437_, _20436_, _05997_);
  or _43248_ (_20438_, _20437_, _20433_);
  and _43249_ (_20439_, _20438_, _05920_);
  or _43250_ (_20440_, _20439_, _20429_);
  and _43251_ (_20441_, _20440_, _06033_);
  or _43252_ (_20442_, _20441_, _20419_);
  and _43253_ (_20443_, _20442_, _05776_);
  or _43254_ (_20444_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or _43255_ (_20445_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and _43256_ (_20446_, _20445_, _05997_);
  and _43257_ (_20447_, _20446_, _20444_);
  or _43258_ (_20448_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _43259_ (_20449_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and _43260_ (_20450_, _20449_, _05996_);
  and _43261_ (_20451_, _20450_, _20448_);
  or _43262_ (_20452_, _20451_, _20447_);
  and _43263_ (_20453_, _20452_, _06021_);
  or _43264_ (_20454_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or _43265_ (_20455_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and _43266_ (_20456_, _20455_, _05997_);
  and _43267_ (_20457_, _20456_, _20454_);
  or _43268_ (_20458_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _43269_ (_20459_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and _43270_ (_20460_, _20459_, _05996_);
  and _43271_ (_20461_, _20460_, _20458_);
  or _43272_ (_20462_, _20461_, _20457_);
  and _43273_ (_20463_, _20462_, _05920_);
  or _43274_ (_20464_, _20463_, _20453_);
  and _43275_ (_20465_, _20464_, _05933_);
  and _43276_ (_20466_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and _43277_ (_20467_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _43278_ (_20468_, _20467_, _20466_);
  and _43279_ (_20469_, _20468_, _05996_);
  and _43280_ (_20470_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and _43281_ (_20471_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _43282_ (_20472_, _20471_, _20470_);
  and _43283_ (_20473_, _20472_, _05997_);
  or _43284_ (_20474_, _20473_, _20469_);
  and _43285_ (_20475_, _20474_, _06021_);
  and _43286_ (_20476_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and _43287_ (_20477_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _43288_ (_20478_, _20477_, _20476_);
  and _43289_ (_20479_, _20478_, _05996_);
  and _43290_ (_20480_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and _43291_ (_20481_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _43292_ (_20482_, _20481_, _20480_);
  and _43293_ (_20483_, _20482_, _05997_);
  or _43294_ (_20484_, _20483_, _20479_);
  and _43295_ (_20485_, _20484_, _05920_);
  or _43296_ (_20486_, _20485_, _20475_);
  and _43297_ (_20487_, _20486_, _06033_);
  or _43298_ (_20488_, _20487_, _20465_);
  and _43299_ (_20489_, _20488_, _06071_);
  or _43300_ (_20490_, _20489_, _20443_);
  and _43301_ (_20491_, _20490_, _05822_);
  or _43302_ (_20492_, _20491_, _20397_);
  or _43303_ (_20493_, _20492_, _06616_);
  and _43304_ (_20494_, _20493_, _20303_);
  or _43305_ (_20495_, _20494_, _06020_);
  and _43306_ (_20496_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and _43307_ (_20497_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _43308_ (_20498_, _20497_, _20496_);
  and _43309_ (_20499_, _20498_, _05996_);
  and _43310_ (_20500_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and _43311_ (_20501_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _43312_ (_20502_, _20501_, _20500_);
  and _43313_ (_20503_, _20502_, _05997_);
  or _43314_ (_20504_, _20503_, _20499_);
  or _43315_ (_20505_, _20504_, _06021_);
  and _43316_ (_20506_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and _43317_ (_20507_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _43318_ (_20508_, _20507_, _20506_);
  and _43319_ (_20509_, _20508_, _05996_);
  and _43320_ (_20510_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and _43321_ (_20511_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _43322_ (_20512_, _20511_, _20510_);
  and _43323_ (_20513_, _20512_, _05997_);
  or _43324_ (_20514_, _20513_, _20509_);
  or _43325_ (_20515_, _20514_, _05920_);
  and _43326_ (_20516_, _20515_, _06033_);
  and _43327_ (_20517_, _20516_, _20505_);
  or _43328_ (_20518_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _43329_ (_20519_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and _43330_ (_20520_, _20519_, _20518_);
  and _43331_ (_20521_, _20520_, _05996_);
  or _43332_ (_20522_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _43333_ (_20523_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and _43334_ (_20524_, _20523_, _20522_);
  and _43335_ (_20525_, _20524_, _05997_);
  or _43336_ (_20526_, _20525_, _20521_);
  or _43337_ (_20527_, _20526_, _06021_);
  or _43338_ (_20528_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _43339_ (_20529_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and _43340_ (_20530_, _20529_, _20528_);
  and _43341_ (_20531_, _20530_, _05996_);
  or _43342_ (_20532_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _43343_ (_20534_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and _43344_ (_20535_, _20534_, _20532_);
  and _43345_ (_20536_, _20535_, _05997_);
  or _43346_ (_20537_, _20536_, _20531_);
  or _43347_ (_20538_, _20537_, _05920_);
  and _43348_ (_20539_, _20538_, _05933_);
  and _43349_ (_20540_, _20539_, _20527_);
  or _43350_ (_20541_, _20540_, _20517_);
  and _43351_ (_20542_, _20541_, _05776_);
  and _43352_ (_20543_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _43353_ (_20544_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _43354_ (_20545_, _20544_, _20543_);
  and _43355_ (_20546_, _20545_, _05996_);
  and _43356_ (_20547_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _43357_ (_20548_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or _43358_ (_20549_, _20548_, _20547_);
  and _43359_ (_20550_, _20549_, _05997_);
  or _43360_ (_20551_, _20550_, _20546_);
  or _43361_ (_20552_, _20551_, _06021_);
  and _43362_ (_20553_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _43363_ (_20554_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _43364_ (_20555_, _20554_, _20553_);
  and _43365_ (_20556_, _20555_, _05996_);
  and _43366_ (_20557_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _43367_ (_20558_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _43368_ (_20559_, _20558_, _20557_);
  and _43369_ (_20560_, _20559_, _05997_);
  or _43370_ (_20561_, _20560_, _20556_);
  or _43371_ (_20562_, _20561_, _05920_);
  and _43372_ (_20563_, _20562_, _06033_);
  and _43373_ (_20564_, _20563_, _20552_);
  or _43374_ (_20565_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _43375_ (_20566_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _43376_ (_20567_, _20566_, _05997_);
  and _43377_ (_20568_, _20567_, _20565_);
  or _43378_ (_20569_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or _43379_ (_20570_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _43380_ (_20571_, _20570_, _05996_);
  and _43381_ (_20572_, _20571_, _20569_);
  or _43382_ (_20573_, _20572_, _20568_);
  or _43383_ (_20574_, _20573_, _06021_);
  or _43384_ (_20575_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _43385_ (_20576_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _43386_ (_20577_, _20576_, _05997_);
  and _43387_ (_20578_, _20577_, _20575_);
  or _43388_ (_20579_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or _43389_ (_20580_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _43390_ (_20581_, _20580_, _05996_);
  and _43391_ (_20582_, _20581_, _20579_);
  or _43392_ (_20583_, _20582_, _20578_);
  or _43393_ (_20584_, _20583_, _05920_);
  and _43394_ (_20585_, _20584_, _05933_);
  and _43395_ (_20586_, _20585_, _20574_);
  or _43396_ (_20587_, _20586_, _20564_);
  and _43397_ (_20588_, _20587_, _06071_);
  or _43398_ (_20589_, _20588_, _20542_);
  and _43399_ (_20590_, _20589_, _06070_);
  and _43400_ (_20591_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _43401_ (_20592_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or _43402_ (_20593_, _20592_, _20591_);
  and _43403_ (_20594_, _20593_, _05996_);
  and _43404_ (_20595_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _43405_ (_20596_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _43406_ (_20597_, _20596_, _20595_);
  and _43407_ (_20598_, _20597_, _05997_);
  or _43408_ (_20599_, _20598_, _20594_);
  and _43409_ (_20600_, _20599_, _05920_);
  and _43410_ (_20601_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _43411_ (_20602_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or _43412_ (_20603_, _20602_, _20601_);
  and _43413_ (_20604_, _20603_, _05996_);
  and _43414_ (_20605_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _43415_ (_20606_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or _43416_ (_20607_, _20606_, _20605_);
  and _43417_ (_20608_, _20607_, _05997_);
  or _43418_ (_20609_, _20608_, _20604_);
  and _43419_ (_20610_, _20609_, _06021_);
  or _43420_ (_20611_, _20610_, _20600_);
  and _43421_ (_20612_, _20611_, _06033_);
  or _43422_ (_20613_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _43423_ (_20614_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _43424_ (_20615_, _20614_, _05997_);
  and _43425_ (_20616_, _20615_, _20613_);
  or _43426_ (_20617_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _43427_ (_20618_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and _43428_ (_20619_, _20618_, _05996_);
  and _43429_ (_20620_, _20619_, _20617_);
  or _43430_ (_20621_, _20620_, _20616_);
  and _43431_ (_20622_, _20621_, _05920_);
  or _43432_ (_20623_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _43433_ (_20624_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _43434_ (_20625_, _20624_, _05997_);
  and _43435_ (_20626_, _20625_, _20623_);
  or _43436_ (_20627_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or _43437_ (_20628_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _43438_ (_20629_, _20628_, _05996_);
  and _43439_ (_20630_, _20629_, _20627_);
  or _43440_ (_20631_, _20630_, _20626_);
  and _43441_ (_20632_, _20631_, _06021_);
  or _43442_ (_20633_, _20632_, _20622_);
  and _43443_ (_20634_, _20633_, _05933_);
  or _43444_ (_20635_, _20634_, _20612_);
  and _43445_ (_20636_, _20635_, _06071_);
  and _43446_ (_20637_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and _43447_ (_20638_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _43448_ (_20639_, _20638_, _20637_);
  and _43449_ (_20640_, _20639_, _05996_);
  and _43450_ (_20641_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and _43451_ (_20642_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _43452_ (_20643_, _20642_, _20641_);
  and _43453_ (_20644_, _20643_, _05997_);
  or _43454_ (_20645_, _20644_, _20640_);
  and _43455_ (_20646_, _20645_, _05920_);
  and _43456_ (_20647_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and _43457_ (_20648_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _43458_ (_20649_, _20648_, _20647_);
  and _43459_ (_20650_, _20649_, _05996_);
  and _43460_ (_20651_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _43461_ (_20652_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _43462_ (_20653_, _20652_, _20651_);
  and _43463_ (_20654_, _20653_, _05997_);
  or _43464_ (_20655_, _20654_, _20650_);
  and _43465_ (_20656_, _20655_, _06021_);
  or _43466_ (_20657_, _20656_, _20646_);
  and _43467_ (_20658_, _20657_, _06033_);
  or _43468_ (_20659_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _43469_ (_20660_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _43470_ (_20661_, _20660_, _20659_);
  and _43471_ (_20662_, _20661_, _05996_);
  or _43472_ (_20663_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _43473_ (_20664_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and _43474_ (_20665_, _20664_, _20663_);
  and _43475_ (_20666_, _20665_, _05997_);
  or _43476_ (_20667_, _20666_, _20662_);
  and _43477_ (_20668_, _20667_, _05920_);
  or _43478_ (_20669_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _43479_ (_20670_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _43480_ (_20671_, _20670_, _20669_);
  and _43481_ (_20672_, _20671_, _05996_);
  or _43482_ (_20673_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _43483_ (_20674_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and _43484_ (_20675_, _20674_, _20673_);
  and _43485_ (_20676_, _20675_, _05997_);
  or _43486_ (_20677_, _20676_, _20672_);
  and _43487_ (_20678_, _20677_, _06021_);
  or _43488_ (_20679_, _20678_, _20668_);
  and _43489_ (_20680_, _20679_, _05933_);
  or _43490_ (_20681_, _20680_, _20658_);
  and _43491_ (_20682_, _20681_, _05776_);
  or _43492_ (_20683_, _20682_, _20636_);
  and _43493_ (_20684_, _20683_, _05822_);
  or _43494_ (_20685_, _20684_, _20590_);
  or _43495_ (_20686_, _20685_, _05868_);
  and _43496_ (_20687_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and _43497_ (_20688_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _43498_ (_20689_, _20688_, _20687_);
  and _43499_ (_20690_, _20689_, _05996_);
  and _43500_ (_20691_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and _43501_ (_20692_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _43502_ (_20693_, _20692_, _20691_);
  and _43503_ (_20694_, _20693_, _05997_);
  or _43504_ (_20695_, _20694_, _20690_);
  or _43505_ (_20696_, _20695_, _06021_);
  and _43506_ (_20697_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and _43507_ (_20698_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _43508_ (_20699_, _20698_, _20697_);
  and _43509_ (_20700_, _20699_, _05996_);
  and _43510_ (_20701_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and _43511_ (_20702_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _43512_ (_20703_, _20702_, _20701_);
  and _43513_ (_20704_, _20703_, _05997_);
  or _43514_ (_20705_, _20704_, _20700_);
  or _43515_ (_20706_, _20705_, _05920_);
  and _43516_ (_20707_, _20706_, _06033_);
  and _43517_ (_20708_, _20707_, _20696_);
  or _43518_ (_20709_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _43519_ (_20710_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and _43520_ (_20711_, _20710_, _05997_);
  and _43521_ (_20712_, _20711_, _20709_);
  or _43522_ (_20713_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _43523_ (_20714_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and _43524_ (_20715_, _20714_, _05996_);
  and _43525_ (_20716_, _20715_, _20713_);
  or _43526_ (_20717_, _20716_, _20712_);
  or _43527_ (_20718_, _20717_, _06021_);
  or _43528_ (_20719_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _43529_ (_20720_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and _43530_ (_20721_, _20720_, _05997_);
  and _43531_ (_20722_, _20721_, _20719_);
  or _43532_ (_20723_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _43533_ (_20724_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and _43534_ (_20725_, _20724_, _05996_);
  and _43535_ (_20726_, _20725_, _20723_);
  or _43536_ (_20727_, _20726_, _20722_);
  or _43537_ (_20728_, _20727_, _05920_);
  and _43538_ (_20729_, _20728_, _05933_);
  and _43539_ (_20730_, _20729_, _20718_);
  or _43540_ (_20731_, _20730_, _20708_);
  and _43541_ (_20732_, _20731_, _06071_);
  and _43542_ (_20733_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _43543_ (_20734_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _43544_ (_20735_, _20734_, _20733_);
  and _43545_ (_20736_, _20735_, _05996_);
  and _43546_ (_20737_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _43547_ (_20738_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or _43548_ (_20739_, _20738_, _20737_);
  and _43549_ (_20740_, _20739_, _05997_);
  or _43550_ (_20741_, _20740_, _20736_);
  or _43551_ (_20742_, _20741_, _06021_);
  and _43552_ (_20743_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and _43553_ (_20744_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or _43554_ (_20745_, _20744_, _20743_);
  and _43555_ (_20746_, _20745_, _05996_);
  and _43556_ (_20747_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _43557_ (_20748_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _43558_ (_20749_, _20748_, _20747_);
  and _43559_ (_20750_, _20749_, _05997_);
  or _43560_ (_20751_, _20750_, _20746_);
  or _43561_ (_20752_, _20751_, _05920_);
  and _43562_ (_20753_, _20752_, _06033_);
  and _43563_ (_20754_, _20753_, _20742_);
  or _43564_ (_20755_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _43565_ (_20756_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _43566_ (_20757_, _20756_, _20755_);
  and _43567_ (_20758_, _20757_, _05996_);
  or _43568_ (_20759_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _43569_ (_20760_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _43570_ (_20761_, _20760_, _20759_);
  and _43571_ (_20762_, _20761_, _05997_);
  or _43572_ (_20763_, _20762_, _20758_);
  or _43573_ (_20764_, _20763_, _06021_);
  or _43574_ (_20765_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or _43575_ (_20766_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _43576_ (_20767_, _20766_, _20765_);
  and _43577_ (_20768_, _20767_, _05996_);
  or _43578_ (_20769_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _43579_ (_20770_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _43580_ (_20771_, _20770_, _20769_);
  and _43581_ (_20772_, _20771_, _05997_);
  or _43582_ (_20773_, _20772_, _20768_);
  or _43583_ (_20774_, _20773_, _05920_);
  and _43584_ (_20775_, _20774_, _05933_);
  and _43585_ (_20776_, _20775_, _20764_);
  or _43586_ (_20777_, _20776_, _20754_);
  and _43587_ (_20778_, _20777_, _05776_);
  or _43588_ (_20779_, _20778_, _20732_);
  and _43589_ (_20780_, _20779_, _06070_);
  or _43590_ (_20781_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or _43591_ (_20782_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and _43592_ (_20783_, _20782_, _20781_);
  and _43593_ (_20784_, _20783_, _05996_);
  or _43594_ (_20785_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _43595_ (_20786_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _43596_ (_20787_, _20786_, _20785_);
  and _43597_ (_20788_, _20787_, _05997_);
  or _43598_ (_20789_, _20788_, _20784_);
  and _43599_ (_20790_, _20789_, _06021_);
  or _43600_ (_20791_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _43601_ (_20792_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and _43602_ (_20793_, _20792_, _20791_);
  and _43603_ (_20794_, _20793_, _05996_);
  or _43604_ (_20795_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _43605_ (_20796_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _43606_ (_20797_, _20796_, _20795_);
  and _43607_ (_20798_, _20797_, _05997_);
  or _43608_ (_20799_, _20798_, _20794_);
  and _43609_ (_20800_, _20799_, _05920_);
  or _43610_ (_20801_, _20800_, _20790_);
  and _43611_ (_20802_, _20801_, _05933_);
  and _43612_ (_20803_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and _43613_ (_20804_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _43614_ (_20805_, _20804_, _20803_);
  and _43615_ (_20806_, _20805_, _05996_);
  and _43616_ (_20807_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _43617_ (_20808_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _43618_ (_20809_, _20808_, _20807_);
  and _43619_ (_20810_, _20809_, _05997_);
  or _43620_ (_20811_, _20810_, _20806_);
  and _43621_ (_20812_, _20811_, _06021_);
  and _43622_ (_20813_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _43623_ (_20814_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _43624_ (_20815_, _20814_, _20813_);
  and _43625_ (_20816_, _20815_, _05996_);
  and _43626_ (_20817_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _43627_ (_20818_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or _43628_ (_20819_, _20818_, _20817_);
  and _43629_ (_20820_, _20819_, _05997_);
  or _43630_ (_20821_, _20820_, _20816_);
  and _43631_ (_20822_, _20821_, _05920_);
  or _43632_ (_20823_, _20822_, _20812_);
  and _43633_ (_20824_, _20823_, _06033_);
  or _43634_ (_20825_, _20824_, _20802_);
  and _43635_ (_20826_, _20825_, _05776_);
  or _43636_ (_20827_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _43637_ (_20828_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and _43638_ (_20829_, _20828_, _05997_);
  and _43639_ (_20830_, _20829_, _20827_);
  or _43640_ (_20831_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _43641_ (_20832_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and _43642_ (_20833_, _20832_, _05996_);
  and _43643_ (_20834_, _20833_, _20831_);
  or _43644_ (_20835_, _20834_, _20830_);
  and _43645_ (_20836_, _20835_, _06021_);
  or _43646_ (_20837_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _43647_ (_20838_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and _43648_ (_20839_, _20838_, _05997_);
  and _43649_ (_20840_, _20839_, _20837_);
  or _43650_ (_20841_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or _43651_ (_20842_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and _43652_ (_20843_, _20842_, _05996_);
  and _43653_ (_20844_, _20843_, _20841_);
  or _43654_ (_20845_, _20844_, _20840_);
  and _43655_ (_20846_, _20845_, _05920_);
  or _43656_ (_20847_, _20846_, _20836_);
  and _43657_ (_20848_, _20847_, _05933_);
  and _43658_ (_20849_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and _43659_ (_20850_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _43660_ (_20851_, _20850_, _20849_);
  and _43661_ (_20852_, _20851_, _05996_);
  and _43662_ (_20853_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and _43663_ (_20854_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _43664_ (_20855_, _20854_, _20853_);
  and _43665_ (_20856_, _20855_, _05997_);
  or _43666_ (_20857_, _20856_, _20852_);
  and _43667_ (_20858_, _20857_, _06021_);
  and _43668_ (_20859_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and _43669_ (_20860_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _43670_ (_20861_, _20860_, _20859_);
  and _43671_ (_20862_, _20861_, _05996_);
  and _43672_ (_20863_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and _43673_ (_20864_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _43674_ (_20865_, _20864_, _20863_);
  and _43675_ (_20866_, _20865_, _05997_);
  or _43676_ (_20867_, _20866_, _20862_);
  and _43677_ (_20868_, _20867_, _05920_);
  or _43678_ (_20869_, _20868_, _20858_);
  and _43679_ (_20870_, _20869_, _06033_);
  or _43680_ (_20871_, _20870_, _20848_);
  and _43681_ (_20872_, _20871_, _06071_);
  or _43682_ (_20873_, _20872_, _20826_);
  and _43683_ (_20874_, _20873_, _05822_);
  or _43684_ (_20875_, _20874_, _20780_);
  or _43685_ (_20876_, _20875_, _06616_);
  and _43686_ (_20877_, _20876_, _20686_);
  or _43687_ (_20878_, _20877_, _05584_);
  and _43688_ (_20879_, _20878_, _20495_);
  or _43689_ (_20880_, _20879_, _06019_);
  or _43690_ (_20881_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _43691_ (_20882_, _20881_, _25365_);
  and _43692_ (_14808_, _20882_, _20880_);
  and _43693_ (_20883_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and _43694_ (_20884_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _43695_ (_20885_, _20884_, _20883_);
  and _43696_ (_20886_, _20885_, _05996_);
  and _43697_ (_20887_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and _43698_ (_20888_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _43699_ (_20889_, _20888_, _20887_);
  and _43700_ (_20890_, _20889_, _05997_);
  or _43701_ (_20891_, _20890_, _20886_);
  or _43702_ (_20892_, _20891_, _06021_);
  and _43703_ (_20893_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and _43704_ (_20894_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _43705_ (_20895_, _20894_, _20893_);
  and _43706_ (_20896_, _20895_, _05996_);
  and _43707_ (_20897_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and _43708_ (_20898_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _43709_ (_20899_, _20898_, _20897_);
  and _43710_ (_20900_, _20899_, _05997_);
  or _43711_ (_20901_, _20900_, _20896_);
  or _43712_ (_20902_, _20901_, _05920_);
  and _43713_ (_20903_, _20902_, _06033_);
  and _43714_ (_20904_, _20903_, _20892_);
  or _43715_ (_20905_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _43716_ (_20906_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and _43717_ (_20907_, _20906_, _20905_);
  and _43718_ (_20908_, _20907_, _05996_);
  or _43719_ (_20909_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _43720_ (_20910_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and _43721_ (_20911_, _20910_, _20909_);
  and _43722_ (_20912_, _20911_, _05997_);
  or _43723_ (_20913_, _20912_, _20908_);
  or _43724_ (_20914_, _20913_, _06021_);
  or _43725_ (_20915_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _43726_ (_20916_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and _43727_ (_20917_, _20916_, _20915_);
  and _43728_ (_20918_, _20917_, _05996_);
  or _43729_ (_20919_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _43730_ (_20920_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and _43731_ (_20921_, _20920_, _20919_);
  and _43732_ (_20922_, _20921_, _05997_);
  or _43733_ (_20923_, _20922_, _20918_);
  or _43734_ (_20924_, _20923_, _05920_);
  and _43735_ (_20925_, _20924_, _05933_);
  and _43736_ (_20926_, _20925_, _20914_);
  or _43737_ (_20927_, _20926_, _20904_);
  and _43738_ (_20928_, _20927_, _05776_);
  and _43739_ (_20929_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and _43740_ (_20930_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _43741_ (_20931_, _20930_, _20929_);
  and _43742_ (_20932_, _20931_, _05996_);
  and _43743_ (_20933_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and _43744_ (_20934_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _43745_ (_20935_, _20934_, _20933_);
  and _43746_ (_20936_, _20935_, _05997_);
  or _43747_ (_20937_, _20936_, _20932_);
  or _43748_ (_20938_, _20937_, _06021_);
  and _43749_ (_20939_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and _43750_ (_20940_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _43751_ (_20941_, _20940_, _20939_);
  and _43752_ (_20942_, _20941_, _05996_);
  and _43753_ (_20943_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and _43754_ (_20944_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _43755_ (_20945_, _20944_, _20943_);
  and _43756_ (_20946_, _20945_, _05997_);
  or _43757_ (_20947_, _20946_, _20942_);
  or _43758_ (_20948_, _20947_, _05920_);
  and _43759_ (_20949_, _20948_, _06033_);
  and _43760_ (_20950_, _20949_, _20938_);
  or _43761_ (_20951_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _43762_ (_20952_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and _43763_ (_20953_, _20952_, _05997_);
  and _43764_ (_20954_, _20953_, _20951_);
  or _43765_ (_20955_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _43766_ (_20956_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and _43767_ (_20957_, _20956_, _05996_);
  and _43768_ (_20958_, _20957_, _20955_);
  or _43769_ (_20959_, _20958_, _20954_);
  or _43770_ (_20960_, _20959_, _06021_);
  or _43771_ (_20961_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _43772_ (_20962_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and _43773_ (_20963_, _20962_, _05997_);
  and _43774_ (_20964_, _20963_, _20961_);
  or _43775_ (_20965_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _43776_ (_20966_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and _43777_ (_20967_, _20966_, _05996_);
  and _43778_ (_20968_, _20967_, _20965_);
  or _43779_ (_20969_, _20968_, _20964_);
  or _43780_ (_20970_, _20969_, _05920_);
  and _43781_ (_20971_, _20970_, _05933_);
  and _43782_ (_20972_, _20971_, _20960_);
  or _43783_ (_20973_, _20972_, _20950_);
  and _43784_ (_20974_, _20973_, _06071_);
  or _43785_ (_20975_, _20974_, _20928_);
  and _43786_ (_20976_, _20975_, _06070_);
  and _43787_ (_20977_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _43788_ (_20978_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _43789_ (_20979_, _20978_, _20977_);
  and _43790_ (_20980_, _20979_, _05996_);
  and _43791_ (_20981_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _43792_ (_20982_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _43793_ (_20983_, _20982_, _20981_);
  and _43794_ (_20984_, _20983_, _05997_);
  or _43795_ (_20985_, _20984_, _20980_);
  and _43796_ (_20986_, _20985_, _05920_);
  and _43797_ (_20987_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _43798_ (_20988_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _43799_ (_20989_, _20988_, _20987_);
  and _43800_ (_20990_, _20989_, _05996_);
  and _43801_ (_20991_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _43802_ (_20992_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _43803_ (_20993_, _20992_, _20991_);
  and _43804_ (_20994_, _20993_, _05997_);
  or _43805_ (_20995_, _20994_, _20990_);
  and _43806_ (_20996_, _20995_, _06021_);
  or _43807_ (_20997_, _20996_, _20986_);
  and _43808_ (_20998_, _20997_, _06033_);
  or _43809_ (_20999_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _43810_ (_21000_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _43811_ (_21001_, _21000_, _05997_);
  and _43812_ (_21002_, _21001_, _20999_);
  or _43813_ (_21003_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _43814_ (_21004_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _43815_ (_21005_, _21004_, _05996_);
  and _43816_ (_21006_, _21005_, _21003_);
  or _43817_ (_21007_, _21006_, _21002_);
  and _43818_ (_21008_, _21007_, _05920_);
  or _43819_ (_21009_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _43820_ (_21010_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _43821_ (_21011_, _21010_, _05997_);
  and _43822_ (_21012_, _21011_, _21009_);
  or _43823_ (_21013_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _43824_ (_21014_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and _43825_ (_21015_, _21014_, _05996_);
  and _43826_ (_21016_, _21015_, _21013_);
  or _43827_ (_21017_, _21016_, _21012_);
  and _43828_ (_21018_, _21017_, _06021_);
  or _43829_ (_21019_, _21018_, _21008_);
  and _43830_ (_21020_, _21019_, _05933_);
  or _43831_ (_21021_, _21020_, _20998_);
  and _43832_ (_21022_, _21021_, _06071_);
  and _43833_ (_21023_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and _43834_ (_21024_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _43835_ (_21025_, _21024_, _21023_);
  and _43836_ (_21026_, _21025_, _05996_);
  and _43837_ (_21027_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and _43838_ (_21028_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _43839_ (_21029_, _21028_, _21027_);
  and _43840_ (_21030_, _21029_, _05997_);
  or _43841_ (_21031_, _21030_, _21026_);
  and _43842_ (_21032_, _21031_, _05920_);
  and _43843_ (_21033_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and _43844_ (_21034_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _43845_ (_21035_, _21034_, _21033_);
  and _43846_ (_21036_, _21035_, _05996_);
  and _43847_ (_21037_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and _43848_ (_21038_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _43849_ (_21039_, _21038_, _21037_);
  and _43850_ (_21040_, _21039_, _05997_);
  or _43851_ (_21041_, _21040_, _21036_);
  and _43852_ (_21042_, _21041_, _06021_);
  or _43853_ (_21043_, _21042_, _21032_);
  and _43854_ (_21044_, _21043_, _06033_);
  or _43855_ (_21045_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _43856_ (_21046_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and _43857_ (_21047_, _21046_, _21045_);
  and _43858_ (_21048_, _21047_, _05996_);
  or _43859_ (_21049_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _43860_ (_21050_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and _43861_ (_21051_, _21050_, _21049_);
  and _43862_ (_21052_, _21051_, _05997_);
  or _43863_ (_21053_, _21052_, _21048_);
  and _43864_ (_21054_, _21053_, _05920_);
  or _43865_ (_21055_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _43866_ (_21056_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and _43867_ (_21057_, _21056_, _21055_);
  and _43868_ (_21058_, _21057_, _05996_);
  or _43869_ (_21059_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _43870_ (_21060_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and _43871_ (_21061_, _21060_, _21059_);
  and _43872_ (_21062_, _21061_, _05997_);
  or _43873_ (_21063_, _21062_, _21058_);
  and _43874_ (_21064_, _21063_, _06021_);
  or _43875_ (_21065_, _21064_, _21054_);
  and _43876_ (_21066_, _21065_, _05933_);
  or _43877_ (_21067_, _21066_, _21044_);
  and _43878_ (_21068_, _21067_, _05776_);
  or _43879_ (_21069_, _21068_, _21022_);
  and _43880_ (_21070_, _21069_, _05822_);
  or _43881_ (_21071_, _21070_, _20976_);
  or _43882_ (_21072_, _21071_, _05868_);
  and _43883_ (_21073_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and _43884_ (_21074_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _43885_ (_21075_, _21074_, _21073_);
  and _43886_ (_21076_, _21075_, _05996_);
  and _43887_ (_21077_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and _43888_ (_21078_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _43889_ (_21079_, _21078_, _21077_);
  and _43890_ (_21080_, _21079_, _05997_);
  or _43891_ (_21081_, _21080_, _21076_);
  or _43892_ (_21082_, _21081_, _06021_);
  and _43893_ (_21083_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and _43894_ (_21084_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _43895_ (_21085_, _21084_, _21083_);
  and _43896_ (_21086_, _21085_, _05996_);
  and _43897_ (_21087_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and _43898_ (_21088_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _43899_ (_21089_, _21088_, _21087_);
  and _43900_ (_21090_, _21089_, _05997_);
  or _43901_ (_21091_, _21090_, _21086_);
  or _43902_ (_21092_, _21091_, _05920_);
  and _43903_ (_21093_, _21092_, _06033_);
  and _43904_ (_21094_, _21093_, _21082_);
  or _43905_ (_21095_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _43906_ (_21096_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and _43907_ (_21097_, _21096_, _05997_);
  and _43908_ (_21098_, _21097_, _21095_);
  or _43909_ (_21099_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _43910_ (_21100_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and _43911_ (_21101_, _21100_, _05996_);
  and _43912_ (_21102_, _21101_, _21099_);
  or _43913_ (_21103_, _21102_, _21098_);
  or _43914_ (_21104_, _21103_, _06021_);
  or _43915_ (_21105_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _43916_ (_21106_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and _43917_ (_21107_, _21106_, _05997_);
  and _43918_ (_21108_, _21107_, _21105_);
  or _43919_ (_21109_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _43920_ (_21110_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and _43921_ (_21111_, _21110_, _05996_);
  and _43922_ (_21112_, _21111_, _21109_);
  or _43923_ (_21113_, _21112_, _21108_);
  or _43924_ (_21114_, _21113_, _05920_);
  and _43925_ (_21115_, _21114_, _05933_);
  and _43926_ (_21116_, _21115_, _21104_);
  or _43927_ (_21117_, _21116_, _21094_);
  and _43928_ (_21118_, _21117_, _06071_);
  and _43929_ (_21119_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and _43930_ (_21120_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _43931_ (_21121_, _21120_, _21119_);
  and _43932_ (_21122_, _21121_, _05996_);
  and _43933_ (_21123_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and _43934_ (_21124_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _43935_ (_21125_, _21124_, _21123_);
  and _43936_ (_21126_, _21125_, _05997_);
  or _43937_ (_21127_, _21126_, _21122_);
  or _43938_ (_21128_, _21127_, _06021_);
  and _43939_ (_21129_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and _43940_ (_21130_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _43941_ (_21131_, _21130_, _21129_);
  and _43942_ (_21132_, _21131_, _05996_);
  and _43943_ (_21133_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _43944_ (_21134_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _43945_ (_21135_, _21134_, _21133_);
  and _43946_ (_21136_, _21135_, _05997_);
  or _43947_ (_21137_, _21136_, _21132_);
  or _43948_ (_21138_, _21137_, _05920_);
  and _43949_ (_21139_, _21138_, _06033_);
  and _43950_ (_21140_, _21139_, _21128_);
  or _43951_ (_21141_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _43952_ (_21142_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and _43953_ (_21143_, _21142_, _21141_);
  and _43954_ (_21144_, _21143_, _05996_);
  or _43955_ (_21145_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _43956_ (_21146_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and _43957_ (_21147_, _21146_, _21145_);
  and _43958_ (_21148_, _21147_, _05997_);
  or _43959_ (_21149_, _21148_, _21144_);
  or _43960_ (_21150_, _21149_, _06021_);
  or _43961_ (_21151_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _43962_ (_21152_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and _43963_ (_21153_, _21152_, _21151_);
  and _43964_ (_21154_, _21153_, _05996_);
  or _43965_ (_21155_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _43966_ (_21156_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _43967_ (_21157_, _21156_, _21155_);
  and _43968_ (_21158_, _21157_, _05997_);
  or _43969_ (_21159_, _21158_, _21154_);
  or _43970_ (_21160_, _21159_, _05920_);
  and _43971_ (_21161_, _21160_, _05933_);
  and _43972_ (_21162_, _21161_, _21150_);
  or _43973_ (_21163_, _21162_, _21140_);
  and _43974_ (_21164_, _21163_, _05776_);
  or _43975_ (_21165_, _21164_, _21118_);
  and _43976_ (_21166_, _21165_, _06070_);
  or _43977_ (_21167_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _43978_ (_21168_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and _43979_ (_21169_, _21168_, _21167_);
  and _43980_ (_21170_, _21169_, _05996_);
  or _43981_ (_21171_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _43982_ (_21172_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and _43983_ (_21173_, _21172_, _21171_);
  and _43984_ (_21174_, _21173_, _05997_);
  or _43985_ (_21175_, _21174_, _21170_);
  and _43986_ (_21176_, _21175_, _06021_);
  or _43987_ (_21177_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _43988_ (_21178_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and _43989_ (_21179_, _21178_, _21177_);
  and _43990_ (_21180_, _21179_, _05996_);
  or _43991_ (_21181_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _43992_ (_21182_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and _43993_ (_21183_, _21182_, _21181_);
  and _43994_ (_21184_, _21183_, _05997_);
  or _43995_ (_21185_, _21184_, _21180_);
  and _43996_ (_21186_, _21185_, _05920_);
  or _43997_ (_21187_, _21186_, _21176_);
  and _43998_ (_21188_, _21187_, _05933_);
  and _43999_ (_21189_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and _44000_ (_21190_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _44001_ (_21191_, _21190_, _21189_);
  and _44002_ (_21192_, _21191_, _05996_);
  and _44003_ (_21193_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and _44004_ (_21194_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _44005_ (_21195_, _21194_, _21193_);
  and _44006_ (_21196_, _21195_, _05997_);
  or _44007_ (_21197_, _21196_, _21192_);
  and _44008_ (_21198_, _21197_, _06021_);
  and _44009_ (_21199_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and _44010_ (_21200_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _44011_ (_21201_, _21200_, _21199_);
  and _44012_ (_21202_, _21201_, _05996_);
  and _44013_ (_21203_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and _44014_ (_21204_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _44015_ (_21205_, _21204_, _21203_);
  and _44016_ (_21206_, _21205_, _05997_);
  or _44017_ (_21207_, _21206_, _21202_);
  and _44018_ (_21208_, _21207_, _05920_);
  or _44019_ (_21209_, _21208_, _21198_);
  and _44020_ (_21210_, _21209_, _06033_);
  or _44021_ (_21211_, _21210_, _21188_);
  and _44022_ (_21212_, _21211_, _05776_);
  or _44023_ (_21213_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _44024_ (_21214_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and _44025_ (_21215_, _21214_, _05997_);
  and _44026_ (_21216_, _21215_, _21213_);
  or _44027_ (_21217_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _44028_ (_21218_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _44029_ (_21219_, _21218_, _05996_);
  and _44030_ (_21220_, _21219_, _21217_);
  or _44031_ (_21221_, _21220_, _21216_);
  and _44032_ (_21222_, _21221_, _06021_);
  or _44033_ (_21223_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _44034_ (_21224_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and _44035_ (_21225_, _21224_, _05997_);
  and _44036_ (_21226_, _21225_, _21223_);
  or _44037_ (_21227_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _44038_ (_21228_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and _44039_ (_21229_, _21228_, _05996_);
  and _44040_ (_21230_, _21229_, _21227_);
  or _44041_ (_21231_, _21230_, _21226_);
  and _44042_ (_21232_, _21231_, _05920_);
  or _44043_ (_21233_, _21232_, _21222_);
  and _44044_ (_21234_, _21233_, _05933_);
  and _44045_ (_21235_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and _44046_ (_21236_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _44047_ (_21237_, _21236_, _21235_);
  and _44048_ (_21238_, _21237_, _05996_);
  and _44049_ (_21239_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and _44050_ (_21240_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _44051_ (_21241_, _21240_, _21239_);
  and _44052_ (_21242_, _21241_, _05997_);
  or _44053_ (_21243_, _21242_, _21238_);
  and _44054_ (_21244_, _21243_, _06021_);
  and _44055_ (_21245_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and _44056_ (_21246_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _44057_ (_21247_, _21246_, _21245_);
  and _44058_ (_21248_, _21247_, _05996_);
  and _44059_ (_21249_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and _44060_ (_21250_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _44061_ (_21251_, _21250_, _21249_);
  and _44062_ (_21252_, _21251_, _05997_);
  or _44063_ (_21253_, _21252_, _21248_);
  and _44064_ (_21254_, _21253_, _05920_);
  or _44065_ (_21255_, _21254_, _21244_);
  and _44066_ (_21256_, _21255_, _06033_);
  or _44067_ (_21257_, _21256_, _21234_);
  and _44068_ (_21258_, _21257_, _06071_);
  or _44069_ (_21259_, _21258_, _21212_);
  and _44070_ (_21260_, _21259_, _05822_);
  or _44071_ (_21261_, _21260_, _21166_);
  or _44072_ (_21262_, _21261_, _06616_);
  and _44073_ (_21263_, _21262_, _21072_);
  or _44074_ (_21264_, _21263_, _06020_);
  and _44075_ (_21265_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and _44076_ (_21266_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _44077_ (_21267_, _21266_, _21265_);
  and _44078_ (_21268_, _21267_, _05996_);
  and _44079_ (_21269_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and _44080_ (_21270_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _44081_ (_21271_, _21270_, _21269_);
  and _44082_ (_21272_, _21271_, _05997_);
  or _44083_ (_21273_, _21272_, _21268_);
  or _44084_ (_21274_, _21273_, _06021_);
  and _44085_ (_21275_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and _44086_ (_21276_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _44087_ (_21277_, _21276_, _21275_);
  and _44088_ (_21278_, _21277_, _05996_);
  and _44089_ (_21279_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and _44090_ (_21280_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _44091_ (_21281_, _21280_, _21279_);
  and _44092_ (_21282_, _21281_, _05997_);
  or _44093_ (_21283_, _21282_, _21278_);
  or _44094_ (_21284_, _21283_, _05920_);
  and _44095_ (_21285_, _21284_, _06033_);
  and _44096_ (_21286_, _21285_, _21274_);
  or _44097_ (_21287_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _44098_ (_21288_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and _44099_ (_21289_, _21288_, _21287_);
  and _44100_ (_21290_, _21289_, _05996_);
  or _44101_ (_21291_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _44102_ (_21292_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and _44103_ (_21293_, _21292_, _21291_);
  and _44104_ (_21294_, _21293_, _05997_);
  or _44105_ (_21295_, _21294_, _21290_);
  or _44106_ (_21296_, _21295_, _06021_);
  or _44107_ (_21297_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _44108_ (_21298_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and _44109_ (_21299_, _21298_, _21297_);
  and _44110_ (_21300_, _21299_, _05996_);
  or _44111_ (_21301_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _44112_ (_21302_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and _44113_ (_21303_, _21302_, _21301_);
  and _44114_ (_21304_, _21303_, _05997_);
  or _44115_ (_21305_, _21304_, _21300_);
  or _44116_ (_21306_, _21305_, _05920_);
  and _44117_ (_21307_, _21306_, _05933_);
  and _44118_ (_21308_, _21307_, _21296_);
  or _44119_ (_21309_, _21308_, _21286_);
  and _44120_ (_21310_, _21309_, _05776_);
  and _44121_ (_21311_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and _44122_ (_21312_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _44123_ (_21313_, _21312_, _21311_);
  and _44124_ (_21314_, _21313_, _05996_);
  and _44125_ (_21315_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _44126_ (_21316_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or _44127_ (_21317_, _21316_, _21315_);
  and _44128_ (_21318_, _21317_, _05997_);
  or _44129_ (_21319_, _21318_, _21314_);
  or _44130_ (_21320_, _21319_, _06021_);
  and _44131_ (_21321_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _44132_ (_21322_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _44133_ (_21323_, _21322_, _21321_);
  and _44134_ (_21324_, _21323_, _05996_);
  and _44135_ (_21325_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _44136_ (_21326_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or _44137_ (_21327_, _21326_, _21325_);
  and _44138_ (_21328_, _21327_, _05997_);
  or _44139_ (_21329_, _21328_, _21324_);
  or _44140_ (_21330_, _21329_, _05920_);
  and _44141_ (_21331_, _21330_, _06033_);
  and _44142_ (_21332_, _21331_, _21320_);
  or _44143_ (_21333_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _44144_ (_21334_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _44145_ (_21335_, _21334_, _05997_);
  and _44146_ (_21336_, _21335_, _21333_);
  or _44147_ (_21337_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or _44148_ (_21338_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and _44149_ (_21339_, _21338_, _05996_);
  and _44150_ (_21340_, _21339_, _21337_);
  or _44151_ (_21341_, _21340_, _21336_);
  or _44152_ (_21342_, _21341_, _06021_);
  or _44153_ (_21343_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _44154_ (_21344_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _44155_ (_21345_, _21344_, _05997_);
  and _44156_ (_21346_, _21345_, _21343_);
  or _44157_ (_21347_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or _44158_ (_21348_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and _44159_ (_21349_, _21348_, _05996_);
  and _44160_ (_21350_, _21349_, _21347_);
  or _44161_ (_21351_, _21350_, _21346_);
  or _44162_ (_21352_, _21351_, _05920_);
  and _44163_ (_21353_, _21352_, _05933_);
  and _44164_ (_21354_, _21353_, _21342_);
  or _44165_ (_21355_, _21354_, _21332_);
  and _44166_ (_21356_, _21355_, _06071_);
  or _44167_ (_21357_, _21356_, _21310_);
  and _44168_ (_21358_, _21357_, _06070_);
  and _44169_ (_21359_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and _44170_ (_21360_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or _44171_ (_21361_, _21360_, _21359_);
  and _44172_ (_21362_, _21361_, _05996_);
  and _44173_ (_21363_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and _44174_ (_21364_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or _44175_ (_21365_, _21364_, _21363_);
  and _44176_ (_21366_, _21365_, _05997_);
  or _44177_ (_21367_, _21366_, _21362_);
  and _44178_ (_21368_, _21367_, _05920_);
  and _44179_ (_21369_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and _44180_ (_21370_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or _44181_ (_21371_, _21370_, _21369_);
  and _44182_ (_21372_, _21371_, _05996_);
  and _44183_ (_21373_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and _44184_ (_21374_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or _44185_ (_21375_, _21374_, _21373_);
  and _44186_ (_21376_, _21375_, _05997_);
  or _44187_ (_21377_, _21376_, _21372_);
  and _44188_ (_21378_, _21377_, _06021_);
  or _44189_ (_21379_, _21378_, _21368_);
  and _44190_ (_21380_, _21379_, _06033_);
  or _44191_ (_21381_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or _44192_ (_21382_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and _44193_ (_21383_, _21382_, _05997_);
  and _44194_ (_21384_, _21383_, _21381_);
  or _44195_ (_21385_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or _44196_ (_21386_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and _44197_ (_21387_, _21386_, _05996_);
  and _44198_ (_21388_, _21387_, _21385_);
  or _44199_ (_21389_, _21388_, _21384_);
  and _44200_ (_21390_, _21389_, _05920_);
  or _44201_ (_21391_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or _44202_ (_21392_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and _44203_ (_21393_, _21392_, _05997_);
  and _44204_ (_21394_, _21393_, _21391_);
  or _44205_ (_21395_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or _44206_ (_21396_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and _44207_ (_21397_, _21396_, _05996_);
  and _44208_ (_21398_, _21397_, _21395_);
  or _44209_ (_21399_, _21398_, _21394_);
  and _44210_ (_21400_, _21399_, _06021_);
  or _44211_ (_21401_, _21400_, _21390_);
  and _44212_ (_21402_, _21401_, _05933_);
  or _44213_ (_21403_, _21402_, _21380_);
  and _44214_ (_21404_, _21403_, _06071_);
  and _44215_ (_21405_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _44216_ (_21406_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _44217_ (_21407_, _21406_, _21405_);
  and _44218_ (_21408_, _21407_, _05996_);
  and _44219_ (_21409_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and _44220_ (_21410_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _44221_ (_21411_, _21410_, _21409_);
  and _44222_ (_21412_, _21411_, _05997_);
  or _44223_ (_21413_, _21412_, _21408_);
  and _44224_ (_21414_, _21413_, _05920_);
  and _44225_ (_21415_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _44226_ (_21416_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _44227_ (_21417_, _21416_, _21415_);
  and _44228_ (_21418_, _21417_, _05996_);
  and _44229_ (_21419_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and _44230_ (_21420_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _44231_ (_21421_, _21420_, _21419_);
  and _44232_ (_21422_, _21421_, _05997_);
  or _44233_ (_21423_, _21422_, _21418_);
  and _44234_ (_21424_, _21423_, _06021_);
  or _44235_ (_21425_, _21424_, _21414_);
  and _44236_ (_21426_, _21425_, _06033_);
  or _44237_ (_21427_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _44238_ (_21428_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and _44239_ (_21429_, _21428_, _21427_);
  and _44240_ (_21430_, _21429_, _05996_);
  or _44241_ (_21431_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _44242_ (_21432_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and _44243_ (_21433_, _21432_, _21431_);
  and _44244_ (_21434_, _21433_, _05997_);
  or _44245_ (_21435_, _21434_, _21430_);
  and _44246_ (_21436_, _21435_, _05920_);
  or _44247_ (_21437_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _44248_ (_21438_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and _44249_ (_21439_, _21438_, _21437_);
  and _44250_ (_21440_, _21439_, _05996_);
  or _44251_ (_21441_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _44252_ (_21442_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and _44253_ (_21443_, _21442_, _21441_);
  and _44254_ (_21444_, _21443_, _05997_);
  or _44255_ (_21445_, _21444_, _21440_);
  and _44256_ (_21446_, _21445_, _06021_);
  or _44257_ (_21447_, _21446_, _21436_);
  and _44258_ (_21448_, _21447_, _05933_);
  or _44259_ (_21449_, _21448_, _21426_);
  and _44260_ (_21450_, _21449_, _05776_);
  or _44261_ (_21451_, _21450_, _21404_);
  and _44262_ (_21452_, _21451_, _05822_);
  or _44263_ (_21453_, _21452_, _21358_);
  or _44264_ (_21454_, _21453_, _05868_);
  and _44265_ (_21455_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and _44266_ (_21456_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _44267_ (_21457_, _21456_, _21455_);
  and _44268_ (_21458_, _21457_, _05996_);
  and _44269_ (_21459_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and _44270_ (_21460_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _44271_ (_21461_, _21460_, _21459_);
  and _44272_ (_21462_, _21461_, _05997_);
  or _44273_ (_21463_, _21462_, _21458_);
  or _44274_ (_21464_, _21463_, _06021_);
  and _44275_ (_21465_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and _44276_ (_21466_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _44277_ (_21467_, _21466_, _21465_);
  and _44278_ (_21468_, _21467_, _05996_);
  and _44279_ (_21469_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and _44280_ (_21470_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _44281_ (_21471_, _21470_, _21469_);
  and _44282_ (_21472_, _21471_, _05997_);
  or _44283_ (_21473_, _21472_, _21468_);
  or _44284_ (_21474_, _21473_, _05920_);
  and _44285_ (_21475_, _21474_, _06033_);
  and _44286_ (_21476_, _21475_, _21464_);
  or _44287_ (_21477_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _44288_ (_21478_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and _44289_ (_21479_, _21478_, _05997_);
  and _44290_ (_21480_, _21479_, _21477_);
  or _44291_ (_21481_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _44292_ (_21482_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and _44293_ (_21483_, _21482_, _05996_);
  and _44294_ (_21484_, _21483_, _21481_);
  or _44295_ (_21485_, _21484_, _21480_);
  or _44296_ (_21486_, _21485_, _06021_);
  or _44297_ (_21487_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _44298_ (_21488_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and _44299_ (_21489_, _21488_, _05997_);
  and _44300_ (_21490_, _21489_, _21487_);
  or _44301_ (_21491_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _44302_ (_21492_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and _44303_ (_21493_, _21492_, _05996_);
  and _44304_ (_21494_, _21493_, _21491_);
  or _44305_ (_21495_, _21494_, _21490_);
  or _44306_ (_21496_, _21495_, _05920_);
  and _44307_ (_21497_, _21496_, _05933_);
  and _44308_ (_21498_, _21497_, _21486_);
  or _44309_ (_21499_, _21498_, _21476_);
  and _44310_ (_21500_, _21499_, _06071_);
  and _44311_ (_21501_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _44312_ (_21502_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _44313_ (_21503_, _21502_, _21501_);
  and _44314_ (_21504_, _21503_, _05996_);
  and _44315_ (_21505_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and _44316_ (_21506_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or _44317_ (_21507_, _21506_, _21505_);
  and _44318_ (_21508_, _21507_, _05997_);
  or _44319_ (_21509_, _21508_, _21504_);
  or _44320_ (_21510_, _21509_, _06021_);
  and _44321_ (_21511_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _44322_ (_21512_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or _44323_ (_21513_, _21512_, _21511_);
  and _44324_ (_21514_, _21513_, _05996_);
  and _44325_ (_21515_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _44326_ (_21516_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _44327_ (_21517_, _21516_, _21515_);
  and _44328_ (_21518_, _21517_, _05997_);
  or _44329_ (_21519_, _21518_, _21514_);
  or _44330_ (_21520_, _21519_, _05920_);
  and _44331_ (_21521_, _21520_, _06033_);
  and _44332_ (_21522_, _21521_, _21510_);
  or _44333_ (_21523_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or _44334_ (_21524_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and _44335_ (_21525_, _21524_, _21523_);
  and _44336_ (_21526_, _21525_, _05996_);
  or _44337_ (_21527_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _44338_ (_21528_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _44339_ (_21529_, _21528_, _21527_);
  and _44340_ (_21530_, _21529_, _05997_);
  or _44341_ (_21531_, _21530_, _21526_);
  or _44342_ (_21532_, _21531_, _06021_);
  or _44343_ (_21533_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or _44344_ (_21534_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _44345_ (_21535_, _21534_, _21533_);
  and _44346_ (_21536_, _21535_, _05996_);
  or _44347_ (_21537_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _44348_ (_21538_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _44349_ (_21539_, _21538_, _21537_);
  and _44350_ (_21540_, _21539_, _05997_);
  or _44351_ (_21541_, _21540_, _21536_);
  or _44352_ (_21542_, _21541_, _05920_);
  and _44353_ (_21543_, _21542_, _05933_);
  and _44354_ (_21544_, _21543_, _21532_);
  or _44355_ (_21545_, _21544_, _21522_);
  and _44356_ (_21546_, _21545_, _05776_);
  or _44357_ (_21547_, _21546_, _21500_);
  and _44358_ (_21548_, _21547_, _06070_);
  or _44359_ (_21549_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _44360_ (_21550_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and _44361_ (_21551_, _21550_, _21549_);
  and _44362_ (_21552_, _21551_, _05996_);
  or _44363_ (_21553_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or _44364_ (_21554_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _44365_ (_21555_, _21554_, _21553_);
  and _44366_ (_21556_, _21555_, _05997_);
  or _44367_ (_21557_, _21556_, _21552_);
  and _44368_ (_21558_, _21557_, _06021_);
  or _44369_ (_21559_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or _44370_ (_21560_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and _44371_ (_21561_, _21560_, _21559_);
  and _44372_ (_21562_, _21561_, _05996_);
  or _44373_ (_21563_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or _44374_ (_21564_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _44375_ (_21565_, _21564_, _21563_);
  and _44376_ (_21566_, _21565_, _05997_);
  or _44377_ (_21567_, _21566_, _21562_);
  and _44378_ (_21568_, _21567_, _05920_);
  or _44379_ (_21569_, _21568_, _21558_);
  and _44380_ (_21570_, _21569_, _05933_);
  and _44381_ (_21571_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _44382_ (_21572_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _44383_ (_21573_, _21572_, _21571_);
  and _44384_ (_21574_, _21573_, _05996_);
  and _44385_ (_21575_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and _44386_ (_21576_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or _44387_ (_21577_, _21576_, _21575_);
  and _44388_ (_21578_, _21577_, _05997_);
  or _44389_ (_21579_, _21578_, _21574_);
  and _44390_ (_21580_, _21579_, _06021_);
  and _44391_ (_21581_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and _44392_ (_21582_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or _44393_ (_21583_, _21582_, _21581_);
  and _44394_ (_21584_, _21583_, _05996_);
  and _44395_ (_21585_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _44396_ (_21586_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _44397_ (_21587_, _21586_, _21585_);
  and _44398_ (_21588_, _21587_, _05997_);
  or _44399_ (_21589_, _21588_, _21584_);
  and _44400_ (_21590_, _21589_, _05920_);
  or _44401_ (_21591_, _21590_, _21580_);
  and _44402_ (_21592_, _21591_, _06033_);
  or _44403_ (_21593_, _21592_, _21570_);
  and _44404_ (_21594_, _21593_, _05776_);
  or _44405_ (_21595_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _44406_ (_21596_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _44407_ (_21597_, _21596_, _05997_);
  and _44408_ (_21598_, _21597_, _21595_);
  or _44409_ (_21599_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _44410_ (_21600_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and _44411_ (_21601_, _21600_, _05996_);
  and _44412_ (_21602_, _21601_, _21599_);
  or _44413_ (_21603_, _21602_, _21598_);
  and _44414_ (_21604_, _21603_, _06021_);
  or _44415_ (_21605_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _44416_ (_21606_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and _44417_ (_21607_, _21606_, _05997_);
  and _44418_ (_21608_, _21607_, _21605_);
  or _44419_ (_21609_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _44420_ (_21610_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _44421_ (_21611_, _21610_, _05996_);
  and _44422_ (_21612_, _21611_, _21609_);
  or _44423_ (_21613_, _21612_, _21608_);
  and _44424_ (_21614_, _21613_, _05920_);
  or _44425_ (_21615_, _21614_, _21604_);
  and _44426_ (_21616_, _21615_, _05933_);
  and _44427_ (_21617_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and _44428_ (_21618_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _44429_ (_21619_, _21618_, _21617_);
  and _44430_ (_21620_, _21619_, _05996_);
  and _44431_ (_21621_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and _44432_ (_21622_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _44433_ (_21623_, _21622_, _21621_);
  and _44434_ (_21624_, _21623_, _05997_);
  or _44435_ (_21625_, _21624_, _21620_);
  and _44436_ (_21626_, _21625_, _06021_);
  and _44437_ (_21627_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and _44438_ (_21628_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _44439_ (_21629_, _21628_, _21627_);
  and _44440_ (_21630_, _21629_, _05996_);
  and _44441_ (_21631_, _06022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and _44442_ (_21632_, _05722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _44443_ (_21633_, _21632_, _21631_);
  and _44444_ (_21634_, _21633_, _05997_);
  or _44445_ (_21635_, _21634_, _21630_);
  and _44446_ (_21636_, _21635_, _05920_);
  or _44447_ (_21637_, _21636_, _21626_);
  and _44448_ (_21638_, _21637_, _06033_);
  or _44449_ (_21639_, _21638_, _21616_);
  and _44450_ (_21640_, _21639_, _06071_);
  or _44451_ (_21641_, _21640_, _21594_);
  and _44452_ (_21642_, _21641_, _05822_);
  or _44453_ (_21643_, _21642_, _21548_);
  or _44454_ (_21644_, _21643_, _06616_);
  and _44455_ (_21645_, _21644_, _21454_);
  or _44456_ (_21646_, _21645_, _05584_);
  and _44457_ (_21647_, _21646_, _21264_);
  or _44458_ (_21648_, _21647_, _06019_);
  or _44459_ (_21649_, _09249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _44460_ (_21650_, _21649_, _25365_);
  and _44461_ (_14809_, _21650_, _21648_);
  nor _44462_ (_05692_, _02153_, rst);
  and _44463_ (_21651_, _01760_, _25365_);
  nand _44464_ (_21652_, _21651_, _01989_);
  nor _44465_ (_21653_, _01998_, _01950_);
  or _44466_ (_05693_, _21653_, _21652_);
  not _44467_ (_21654_, _01823_);
  and _44468_ (_21655_, _01846_, _21654_);
  not _44469_ (_21656_, _01977_);
  not _44470_ (_21657_, _01898_);
  and _44471_ (_21658_, _01944_, _01920_);
  and _44472_ (_21659_, _21658_, _21657_);
  and _44473_ (_21660_, _21659_, _01872_);
  and _44474_ (_21661_, _21660_, _21656_);
  and _44475_ (_21662_, _21661_, _21655_);
  not _44476_ (_21663_, _01944_);
  nor _44477_ (_21664_, _21663_, _01920_);
  and _44478_ (_21665_, _21664_, _01898_);
  nor _44479_ (_21666_, _01977_, _01798_);
  nor _44480_ (_21667_, _01846_, _01823_);
  and _44481_ (_21668_, _21667_, _21666_);
  and _44482_ (_21669_, _21668_, _21665_);
  and _44483_ (_21670_, _01977_, _21663_);
  and _44484_ (_21671_, _21667_, _01798_);
  and _44485_ (_21672_, _21671_, _21670_);
  or _44486_ (_21673_, _21672_, _21669_);
  nor _44487_ (_21674_, _21656_, _01798_);
  and _44488_ (_21675_, _21674_, _21655_);
  and _44489_ (_21676_, _21675_, _21659_);
  and _44490_ (_21677_, _21674_, _21667_);
  and _44491_ (_21678_, _21677_, _21665_);
  or _44492_ (_21679_, _21678_, _21676_);
  or _44493_ (_21680_, _21679_, _21673_);
  and _44494_ (_21681_, _21655_, _01798_);
  not _44495_ (_21682_, _01872_);
  and _44496_ (_21683_, _21665_, _21682_);
  and _44497_ (_21684_, _21683_, _21681_);
  and _44498_ (_21685_, _21665_, _01872_);
  and _44499_ (_21686_, _01846_, _01823_);
  and _44500_ (_21687_, _21686_, _01798_);
  and _44501_ (_21688_, _21687_, _21685_);
  or _44502_ (_21689_, _21688_, _21684_);
  or _44503_ (_21690_, _21689_, _21680_);
  or _44504_ (_21691_, _21690_, _21662_);
  and _44505_ (_21692_, _21664_, _21657_);
  not _44506_ (_21693_, _21692_);
  not _44507_ (_21694_, _01846_);
  and _44508_ (_21695_, _21694_, _01823_);
  and _44509_ (_21696_, _21695_, _21666_);
  nor _44510_ (_21697_, _21696_, _21682_);
  nor _44511_ (_21698_, _21697_, _21693_);
  not _44512_ (_21699_, _21698_);
  and _44513_ (_21700_, _21692_, _01872_);
  and _44514_ (_21701_, _21686_, _21674_);
  and _44515_ (_21702_, _21701_, _21700_);
  and _44516_ (_21703_, _21656_, _01798_);
  and _44517_ (_21704_, _21695_, _21703_);
  and _44518_ (_21705_, _21704_, _21700_);
  nor _44519_ (_21706_, _21705_, _21702_);
  and _44520_ (_21707_, _21706_, _21699_);
  and _44521_ (_21708_, _21695_, _21674_);
  and _44522_ (_21709_, _21708_, _21683_);
  and _44523_ (_21710_, _01977_, _01798_);
  and _44524_ (_21711_, _21686_, _21710_);
  and _44525_ (_21712_, _21686_, _21666_);
  or _44526_ (_21713_, _21712_, _21711_);
  and _44527_ (_21714_, _21713_, _21700_);
  nor _44528_ (_21715_, _21714_, _21709_);
  not _44529_ (_21716_, _01798_);
  and _44530_ (_21717_, _21667_, _21716_);
  and _44531_ (_21718_, _21700_, _21717_);
  and _44532_ (_21719_, _21686_, _21716_);
  and _44533_ (_21720_, _21719_, _21685_);
  nor _44534_ (_21721_, _21720_, _21718_);
  and _44535_ (_21722_, _21721_, _21715_);
  and _44536_ (_21723_, _21703_, _21655_);
  and _44537_ (_21724_, _21700_, _21723_);
  and _44538_ (_21725_, _21695_, _01977_);
  and _44539_ (_21726_, _21725_, _21700_);
  nor _44540_ (_21727_, _21726_, _21724_);
  and _44541_ (_21728_, _21710_, _21667_);
  and _44542_ (_21729_, _21659_, _21682_);
  and _44543_ (_21730_, _21729_, _21728_);
  and _44544_ (_21731_, _21655_, _21716_);
  and _44545_ (_21732_, _01977_, _01898_);
  and _44546_ (_21733_, _21732_, _21658_);
  or _44547_ (_21734_, _21733_, _21670_);
  and _44548_ (_21735_, _21734_, _21731_);
  nor _44549_ (_21736_, _21735_, _21730_);
  and _44550_ (_21737_, _21736_, _21727_);
  and _44551_ (_21738_, _21737_, _21722_);
  nand _44552_ (_21739_, _21738_, _21707_);
  or _44553_ (_21740_, _21739_, _21691_);
  and _44554_ (_21741_, _21740_, _01761_);
  not _44555_ (_21742_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _44556_ (_21743_, _01759_, _00000_);
  and _44557_ (_21744_, _21743_, _02077_);
  nor _44558_ (_21745_, _21744_, _21742_);
  or _44559_ (_21746_, _21745_, rst);
  or _44560_ (_05694_, _21746_, _21741_);
  nand _44561_ (_21747_, _01823_, _01755_);
  or _44562_ (_21748_, _01755_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _44563_ (_21749_, _21748_, _25365_);
  and _44564_ (_05695_, _21749_, _21747_);
  and _44565_ (_21750_, \oc8051_top_1.oc8051_sfr1.wait_data , _25365_);
  and _44566_ (_21751_, _21750_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _44567_ (_21752_, _02125_, _02024_);
  and _44568_ (_21753_, _02125_, _02041_);
  and _44569_ (_21754_, _02041_, _02109_);
  or _44570_ (_21755_, _21754_, _21753_);
  or _44571_ (_21756_, _21755_, _21752_);
  and _44572_ (_21757_, _02147_, _01990_);
  and _44573_ (_21758_, _02006_, _02109_);
  or _44574_ (_21759_, _21758_, _21757_);
  and _44575_ (_21760_, _02006_, _01998_);
  and _44576_ (_21761_, _02024_, _02109_);
  or _44577_ (_21762_, _21761_, _21760_);
  or _44578_ (_21763_, _21762_, _02080_);
  or _44579_ (_21764_, _21763_, _21759_);
  or _44580_ (_21765_, _21764_, _21756_);
  or _44581_ (_21766_, _21765_, _02037_);
  and _44582_ (_21767_, _21766_, _21651_);
  or _44583_ (_05696_, _21767_, _21751_);
  and _44584_ (_21768_, _01998_, _02008_);
  or _44585_ (_21769_, _21768_, _02110_);
  and _44586_ (_21770_, _01987_, _01948_);
  and _44587_ (_21771_, _21770_, _02000_);
  or _44588_ (_21772_, _21771_, _02094_);
  and _44589_ (_21773_, _01954_, _01955_);
  and _44590_ (_21774_, _21773_, _02024_);
  or _44591_ (_21775_, _21774_, _21772_);
  or _44592_ (_21776_, _21775_, _21769_);
  and _44593_ (_21777_, _21776_, _01760_);
  and _44594_ (_21778_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _44595_ (_21779_, _02082_, _21742_);
  not _44596_ (_21780_, _02150_);
  and _44597_ (_21781_, _21780_, _21779_);
  or _44598_ (_21782_, _21781_, _21778_);
  or _44599_ (_21783_, _21782_, _21777_);
  and _44600_ (_05697_, _21783_, _25365_);
  and _44601_ (_21784_, _21750_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44602_ (_21785_, _01981_, _01948_);
  and _44603_ (_21786_, _21785_, _02011_);
  not _44604_ (_21787_, _02030_);
  and _44605_ (_21788_, _02147_, _21787_);
  or _44606_ (_21789_, _21788_, _02044_);
  and _44607_ (_21790_, _02147_, _02015_);
  or _44608_ (_21791_, _02042_, _02016_);
  or _44609_ (_21792_, _21791_, _21790_);
  or _44610_ (_21793_, _21792_, _21789_);
  nor _44611_ (_21794_, _02015_, _02041_);
  nor _44612_ (_21795_, _21794_, _01953_);
  and _44613_ (_21796_, _21785_, _02101_);
  nor _44614_ (_21797_, _21796_, _21795_);
  nand _44615_ (_21798_, _21797_, _02103_);
  and _44616_ (_21799_, _02147_, _02008_);
  and _44617_ (_21800_, _02147_, _02052_);
  or _44618_ (_21801_, _21800_, _21799_);
  or _44619_ (_21802_, _21801_, _21769_);
  or _44620_ (_21803_, _21802_, _21798_);
  or _44621_ (_21804_, _21803_, _21793_);
  or _44622_ (_21805_, _21804_, _21786_);
  and _44623_ (_21806_, _21805_, _21651_);
  or _44624_ (_05698_, _21806_, _21784_);
  and _44625_ (_21807_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _44626_ (_21808_, _21807_, _21781_);
  and _44627_ (_21809_, _02007_, _01760_);
  or _44628_ (_21810_, _21809_, _21808_);
  and _44629_ (_05699_, _21810_, _25365_);
  and _44630_ (_21811_, _02112_, _01987_);
  and _44631_ (_21812_, _01956_, _01949_);
  and _44632_ (_21813_, _02101_, _01951_);
  nor _44633_ (_21814_, _21813_, _21812_);
  nor _44634_ (_21815_, _21814_, _01987_);
  or _44635_ (_21816_, _21815_, _21811_);
  and _44636_ (_21817_, _21816_, _01756_);
  and _44637_ (_21818_, _21815_, _02079_);
  not _44638_ (_21819_, _01990_);
  nor _44639_ (_21820_, _21653_, _21819_);
  nor _44640_ (_21821_, _21820_, _02112_);
  not _44641_ (_21822_, _21821_);
  and _44642_ (_21823_, _21822_, _21779_);
  or _44643_ (_21824_, _21823_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _44644_ (_21825_, _21824_, _21818_);
  or _44645_ (_21826_, _21825_, _21817_);
  or _44646_ (_21827_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _00000_);
  and _44647_ (_21828_, _21827_, _25365_);
  and _44648_ (_05700_, _21828_, _21826_);
  and _44649_ (_21829_, _21750_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and _44650_ (_21830_, _02041_, _01950_);
  or _44651_ (_21831_, _21830_, _02064_);
  and _44652_ (_21832_, _02097_, _02101_);
  and _44653_ (_21833_, _02018_, _02024_);
  or _44654_ (_21834_, _21833_, _21832_);
  or _44655_ (_21835_, _21834_, _21831_);
  or _44656_ (_21836_, _02110_, _02042_);
  and _44657_ (_21837_, _02052_, _01951_);
  and _44658_ (_21838_, _21773_, _21787_);
  or _44659_ (_21839_, _21838_, _21837_);
  or _44660_ (_21840_, _21839_, _21836_);
  and _44661_ (_21841_, _21785_, _02000_);
  or _44662_ (_21842_, _21841_, _21796_);
  or _44663_ (_21843_, _21771_, _02025_);
  or _44664_ (_21844_, _21843_, _21842_);
  or _44665_ (_21845_, _21844_, _21840_);
  or _44666_ (_21846_, _21845_, _21835_);
  and _44667_ (_21847_, _21846_, _21651_);
  or _44668_ (_05701_, _21847_, _21829_);
  and _44669_ (_21848_, _21750_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _44670_ (_21849_, _02147_, _01995_);
  or _44671_ (_21850_, _21849_, _02023_);
  nor _44672_ (_21851_, _02102_, _01996_);
  nand _44673_ (_21852_, _21851_, _02050_);
  or _44674_ (_21853_, _21852_, _21850_);
  and _44675_ (_21854_, _02097_, _02000_);
  nor _44676_ (_21855_, _01982_, _01803_);
  and _44677_ (_21856_, _02118_, _21855_);
  or _44678_ (_21857_, _21856_, _02127_);
  or _44679_ (_21858_, _21857_, _21854_);
  not _44680_ (_21859_, _21797_);
  and _44681_ (_21860_, _02109_, _01851_);
  or _44682_ (_21861_, _21860_, _21859_);
  or _44683_ (_21862_, _21861_, _21858_);
  and _44684_ (_21863_, _02125_, _02058_);
  nor _44685_ (_21864_, _21863_, _02056_);
  not _44686_ (_21865_, _21864_);
  and _44687_ (_21866_, _02147_, _02047_);
  or _44688_ (_21867_, _21866_, _21865_);
  and _44689_ (_21868_, _21770_, _21855_);
  and _44690_ (_21869_, _21770_, _01994_);
  or _44691_ (_21870_, _21869_, _21868_);
  or _44692_ (_21871_, _21870_, _21774_);
  or _44693_ (_21872_, _21871_, _21867_);
  or _44694_ (_21873_, _21872_, _21862_);
  or _44695_ (_21874_, _21873_, _21853_);
  or _44696_ (_21875_, _21874_, _21793_);
  and _44697_ (_21876_, _21875_, _21651_);
  or _44698_ (_05702_, _21876_, _21848_);
  and _44699_ (_21877_, _21773_, _01852_);
  or _44700_ (_21878_, _21877_, _02098_);
  and _44701_ (_21879_, _21785_, _02005_);
  or _44702_ (_21880_, _21879_, _02105_);
  and _44703_ (_21881_, _01948_, _01852_);
  or _44704_ (_21882_, _21881_, _21880_);
  or _44705_ (_21883_, _21882_, _21878_);
  and _44706_ (_21884_, _21773_, _02008_);
  or _44707_ (_21885_, _21884_, _21780_);
  or _44708_ (_21886_, _21885_, _21883_);
  and _44709_ (_21887_, _21886_, _21651_);
  nor _44710_ (_21888_, _02150_, _01756_);
  and _44711_ (_21889_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _44712_ (_21890_, _21889_, _21888_);
  and _44713_ (_21891_, _21890_, _25365_);
  or _44714_ (_05703_, _21891_, _21887_);
  and _44715_ (_21892_, _01850_, _01803_);
  and _44716_ (_21893_, _21892_, _01981_);
  and _44717_ (_21894_, _21893_, _01957_);
  or _44718_ (_21895_, _02056_, _02044_);
  or _44719_ (_21896_, _21895_, _21894_);
  and _44720_ (_21897_, _21787_, _01951_);
  or _44721_ (_21898_, _21897_, _02002_);
  or _44722_ (_21899_, _21898_, _21896_);
  nand _44723_ (_21900_, _02055_, _02010_);
  nor _44724_ (_21901_, _21794_, _02043_);
  or _44725_ (_21902_, _21753_, _02025_);
  or _44726_ (_21903_, _21902_, _21901_);
  or _44727_ (_21904_, _21903_, _21900_);
  or _44728_ (_21905_, _21904_, _21899_);
  and _44729_ (_21906_, _21812_, _01981_);
  and _44730_ (_21907_, _21770_, _02005_);
  or _44731_ (_21908_, _21907_, _21906_);
  and _44732_ (_21909_, _21785_, _21892_);
  or _44733_ (_21910_, _21909_, _02013_);
  or _44734_ (_21911_, _21910_, _21772_);
  or _44735_ (_21912_, _21911_, _21908_);
  and _44736_ (_21913_, _02097_, _21892_);
  not _44737_ (_21914_, _02102_);
  nand _44738_ (_21915_, _21914_, _02019_);
  or _44739_ (_21916_, _21915_, _21913_);
  and _44740_ (_21917_, _02018_, _02006_);
  or _44741_ (_21918_, _21917_, _02069_);
  or _44742_ (_21919_, _21918_, _21916_);
  or _44743_ (_21920_, _21919_, _21912_);
  or _44744_ (_21921_, _21920_, _21859_);
  or _44745_ (_21922_, _21921_, _21905_);
  and _44746_ (_21923_, _21922_, _01760_);
  and _44747_ (_21924_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _44748_ (_21925_, _05597_, _02031_);
  and _44749_ (_21926_, _02125_, _21787_);
  or _44750_ (_21927_, _21926_, _21906_);
  and _44751_ (_21928_, _21927_, _02079_);
  or _44752_ (_21929_, _21928_, _21781_);
  or _44753_ (_21930_, _21929_, _21925_);
  or _44754_ (_21931_, _21930_, _21924_);
  or _44755_ (_21932_, _21931_, _21923_);
  and _44756_ (_05705_, _21932_, _25365_);
  and _44757_ (_05706_, _02136_, _25365_);
  and _44758_ (_05707_, _02086_, _25365_);
  not _44759_ (_21933_, _21651_);
  or _44760_ (_05708_, _21821_, _21933_);
  and _44761_ (_21934_, _01998_, _01989_);
  nor _44762_ (_21935_, _21934_, _02112_);
  or _44763_ (_05709_, _21935_, _21933_);
  or _44764_ (_21936_, _21684_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _44765_ (_21937_, _21936_, _21720_);
  or _44766_ (_21938_, _21937_, _21662_);
  and _44767_ (_21939_, _21938_, _21744_);
  nor _44768_ (_21940_, _21743_, _02077_);
  or _44769_ (_21941_, _21940_, rst);
  or _44770_ (_05710_, _21941_, _21939_);
  nand _44771_ (_21942_, _01872_, _01755_);
  or _44772_ (_21943_, _01755_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _44773_ (_21944_, _21943_, _25365_);
  and _44774_ (_05711_, _21944_, _21942_);
  not _44775_ (_21945_, _01755_);
  or _44776_ (_21946_, _01898_, _21945_);
  or _44777_ (_21947_, _01755_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _44778_ (_21948_, _21947_, _25365_);
  and _44779_ (_05712_, _21948_, _21946_);
  or _44780_ (_21949_, _01920_, _21945_);
  or _44781_ (_21950_, _01755_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _44782_ (_21951_, _21950_, _25365_);
  and _44783_ (_05713_, _21951_, _21949_);
  nand _44784_ (_21952_, _01944_, _01755_);
  or _44785_ (_21953_, _01755_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _44786_ (_21954_, _21953_, _25365_);
  and _44787_ (_05714_, _21954_, _21952_);
  or _44788_ (_21955_, _01977_, _21945_);
  or _44789_ (_21956_, _01755_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _44790_ (_21957_, _21956_, _25365_);
  and _44791_ (_05715_, _21957_, _21955_);
  nand _44792_ (_21958_, _01798_, _01755_);
  or _44793_ (_21959_, _01755_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _44794_ (_21960_, _21959_, _25365_);
  and _44795_ (_05716_, _21960_, _21958_);
  nand _44796_ (_21961_, _01846_, _01755_);
  or _44797_ (_21962_, _01755_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _44798_ (_21963_, _21962_, _25365_);
  and _44799_ (_05717_, _21963_, _21961_);
  and _44800_ (_21964_, _02147_, _02041_);
  or _44801_ (_21965_, _21964_, _21788_);
  or _44802_ (_21966_, _21965_, _21790_);
  and _44803_ (_21967_, _21785_, _02046_);
  or _44804_ (_21968_, _21967_, _21881_);
  and _44805_ (_21969_, _21773_, _02047_);
  or _44806_ (_21970_, _21969_, _21768_);
  or _44807_ (_21971_, _21970_, _21968_);
  or _44808_ (_21972_, _21971_, _21966_);
  or _44809_ (_21973_, _21757_, _01991_);
  and _44810_ (_21974_, _02147_, _02058_);
  or _44811_ (_21975_, _21974_, _21869_);
  or _44812_ (_21976_, _21975_, _21973_);
  or _44813_ (_21977_, _21850_, _02110_);
  and _44814_ (_21978_, _21773_, _02066_);
  or _44815_ (_21979_, _21978_, _02127_);
  or _44816_ (_21980_, _21979_, _21884_);
  or _44817_ (_21981_, _21980_, _21977_);
  or _44818_ (_21982_, _21981_, _21976_);
  and _44819_ (_21983_, _21770_, _02046_);
  and _44820_ (_21984_, _21770_, _01989_);
  or _44821_ (_21985_, _21984_, _21983_);
  or _44822_ (_21986_, _21985_, _21860_);
  and _44823_ (_21987_, _01989_, _01981_);
  and _44824_ (_21988_, _21987_, _02147_);
  or _44825_ (_21989_, _21877_, _21880_);
  or _44826_ (_21990_, _21989_, _21988_);
  or _44827_ (_21991_, _21990_, _21986_);
  or _44828_ (_21992_, _02123_, _02098_);
  or _44829_ (_21993_, _21992_, _02104_);
  or _44830_ (_21994_, _21993_, _21991_);
  or _44831_ (_21995_, _21994_, _21982_);
  or _44832_ (_21996_, _21995_, _21972_);
  and _44833_ (_21997_, _21996_, _01760_);
  and _44834_ (_21998_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _44835_ (_21999_, _21998_, _21823_);
  or _44836_ (_22000_, _21999_, _21997_);
  and _44837_ (_05951_, _22000_, _25365_);
  and _44838_ (_22001_, _21750_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _44839_ (_22002_, _21970_, _21858_);
  or _44840_ (_22003_, _22002_, _21759_);
  and _44841_ (_22004_, _02125_, _01993_);
  and _44842_ (_22005_, _22004_, _01987_);
  or _44843_ (_22006_, _21786_, _02100_);
  or _44844_ (_22007_, _22006_, _21870_);
  or _44845_ (_22008_, _22007_, _02026_);
  or _44846_ (_22009_, _22008_, _22005_);
  or _44847_ (_22010_, _02027_, _01995_);
  or _44848_ (_22011_, _02066_, _02033_);
  or _44849_ (_22012_, _22011_, _22010_);
  and _44850_ (_22013_, _22012_, _02147_);
  or _44851_ (_22014_, _22013_, _21801_);
  or _44852_ (_22015_, _22014_, _22009_);
  or _44853_ (_22016_, _22015_, _22003_);
  and _44854_ (_22017_, _22016_, _21651_);
  or _44855_ (_05952_, _22017_, _22001_);
  or _44856_ (_22018_, _21918_, _21908_);
  or _44857_ (_22019_, _22018_, _21905_);
  and _44858_ (_22020_, _22019_, _01760_);
  and _44859_ (_22021_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _44860_ (_22022_, _22021_, _21930_);
  or _44861_ (_22023_, _22022_, _22020_);
  and _44862_ (_05953_, _22023_, _25365_);
  and _44863_ (_22024_, _02001_, _01987_);
  or _44864_ (_22025_, _22024_, _21927_);
  or _44865_ (_22026_, _22025_, _21916_);
  or _44866_ (_22027_, _22026_, _02094_);
  and _44867_ (_22028_, _22027_, _01760_);
  and _44868_ (_22029_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _44869_ (_22030_, _22029_, _21929_);
  or _44870_ (_22031_, _22030_, _22028_);
  and _44871_ (_05954_, _22031_, _25365_);
  or _44872_ (_22032_, _21866_, _21927_);
  or _44873_ (_22033_, _21968_, _21860_);
  and _44874_ (_22034_, _21987_, _01957_);
  or _44875_ (_22035_, _21974_, _22034_);
  or _44876_ (_22036_, _21913_, _21849_);
  or _44877_ (_22037_, _22036_, _22035_);
  or _44878_ (_22038_, _22037_, _22033_);
  or _44879_ (_22039_, _22038_, _22032_);
  and _44880_ (_22040_, _21773_, _02027_);
  or _44881_ (_22041_, _22040_, _02112_);
  or _44882_ (_22042_, _21978_, _02149_);
  or _44883_ (_22043_, _22042_, _22041_);
  and _44884_ (_22044_, _02147_, _02024_);
  or _44885_ (_22045_, _21884_, _22044_);
  and _44886_ (_22046_, _21773_, _02052_);
  or _44887_ (_22047_, _22046_, _21757_);
  or _44888_ (_22048_, _21988_, _02148_);
  or _44889_ (_22049_, _22048_, _22047_);
  or _44890_ (_22050_, _22049_, _21966_);
  or _44891_ (_22051_, _22050_, _22045_);
  and _44892_ (_22052_, _21773_, _02033_);
  and _44893_ (_22053_, _02125_, _02066_);
  or _44894_ (_22054_, _22053_, _21909_);
  or _44895_ (_22055_, _21880_, _02104_);
  or _44896_ (_22056_, _02111_, _02098_);
  or _44897_ (_22057_, _22056_, _22055_);
  or _44898_ (_22058_, _22057_, _22054_);
  or _44899_ (_22059_, _22058_, _22052_);
  or _44900_ (_22060_, _22059_, _22051_);
  or _44901_ (_22061_, _22060_, _22043_);
  or _44902_ (_22062_, _22061_, _22039_);
  and _44903_ (_22063_, _22062_, _01760_);
  and _44904_ (_22064_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _44905_ (_22065_, _21823_, _21888_);
  or _44906_ (_22066_, _22065_, _22064_);
  or _44907_ (_22067_, _22066_, _22063_);
  and _44908_ (_05955_, _22067_, _25365_);
  and _44909_ (_22068_, _02056_, _01876_);
  and _44910_ (_22069_, _02109_, _01995_);
  or _44911_ (_22070_, _02069_, _22069_);
  or _44912_ (_22071_, _22070_, _22068_);
  and _44913_ (_22072_, _02018_, _02008_);
  or _44914_ (_22073_, _02149_, _22072_);
  or _44915_ (_22074_, _21894_, _21768_);
  or _44916_ (_22075_, _22074_, _22073_);
  or _44917_ (_22076_, _22075_, _02143_);
  or _44918_ (_22077_, _22076_, _22071_);
  or _44919_ (_22078_, _22077_, _22033_);
  or _44920_ (_22079_, _21785_, _02097_);
  and _44921_ (_22080_, _22079_, _01989_);
  or _44922_ (_22081_, _22055_, _02068_);
  or _44923_ (_22082_, _22081_, _22080_);
  or _44924_ (_22083_, _22082_, _22051_);
  or _44925_ (_22084_, _22083_, _22078_);
  and _44926_ (_22085_, _22084_, _01760_);
  and _44927_ (_22086_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _44928_ (_22087_, _22086_, _22065_);
  or _44929_ (_22088_, _22087_, _22085_);
  and _44930_ (_05956_, _22088_, _25365_);
  and _44931_ (_22089_, _21750_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _44932_ (_22090_, _02101_, _02109_);
  and _44933_ (_22091_, _22090_, _01981_);
  or _44934_ (_22092_, _22091_, _21754_);
  not _44935_ (_22093_, _05591_);
  or _44936_ (_22094_, _21884_, _22093_);
  and _44937_ (_22095_, _02109_, _02052_);
  or _44938_ (_22096_, _21879_, _21771_);
  or _44939_ (_22097_, _22096_, _22095_);
  and _44940_ (_22098_, _02027_, _02109_);
  and _44941_ (_22099_, _02097_, _01851_);
  or _44942_ (_22100_, _22099_, _22098_);
  or _44943_ (_22101_, _22100_, _22097_);
  or _44944_ (_22102_, _22101_, _22094_);
  or _44945_ (_22103_, _22102_, _22092_);
  or _44946_ (_22104_, _21964_, _21838_);
  or _44947_ (_22105_, _21902_, _21842_);
  or _44948_ (_22106_, _22105_, _22104_);
  and _44949_ (_22107_, _02027_, _01948_);
  or _44950_ (_22108_, _22107_, _22072_);
  or _44951_ (_22109_, _22108_, _02009_);
  and _44952_ (_22110_, _21877_, _01981_);
  or _44953_ (_22111_, _22110_, _21833_);
  or _44954_ (_22112_, _22111_, _22109_);
  not _44955_ (_22113_, _05589_);
  or _44956_ (_22114_, _21836_, _22113_);
  or _44957_ (_22115_, _22114_, _22112_);
  or _44958_ (_22116_, _22115_, _22106_);
  or _44959_ (_22117_, _22116_, _22103_);
  and _44960_ (_22118_, _22117_, _21651_);
  or _44961_ (_05957_, _22118_, _22089_);
  or _44962_ (_22119_, _22043_, _21867_);
  or _44963_ (_22120_, _22052_, _21856_);
  or _44964_ (_22121_, _22120_, _21774_);
  nor _44965_ (_22122_, _02030_, _02141_);
  and _44966_ (_22123_, _02109_, _01852_);
  and _44967_ (_22124_, _22123_, _01981_);
  or _44968_ (_22125_, _22124_, _21964_);
  or _44969_ (_22126_, _22125_, _22122_);
  or _44970_ (_22127_, _22126_, _22121_);
  or _44971_ (_22128_, _02106_, _02071_);
  or _44972_ (_22129_, _21868_, _21854_);
  or _44973_ (_22130_, _22129_, _02110_);
  or _44974_ (_22131_, _02111_, _02048_);
  or _44975_ (_22132_, _22131_, _22130_);
  or _44976_ (_22133_, _22132_, _22128_);
  or _44977_ (_22134_, _22133_, _21968_);
  or _44978_ (_22135_, _22134_, _22127_);
  or _44979_ (_22136_, _22135_, _22119_);
  and _44980_ (_22137_, _22136_, _21651_);
  and _44981_ (_22138_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _44982_ (_22139_, _02149_, _02140_);
  or _44983_ (_22140_, _22139_, _22138_);
  and _44984_ (_22141_, _22140_, _25365_);
  or _44985_ (_05958_, _22141_, _22137_);
  nor _44986_ (_22142_, _22072_, _02094_);
  nor _44987_ (_22143_, _21884_, _21786_);
  nand _44988_ (_22144_, _22143_, _22142_);
  or _44989_ (_22145_, _22144_, _22047_);
  and _44990_ (_22146_, _02052_, _01950_);
  or _44991_ (_22147_, _22146_, _21988_);
  or _44992_ (_22148_, _21967_, _02104_);
  or _44993_ (_22149_, _22148_, _22147_);
  or _44994_ (_22150_, _22149_, _22145_);
  nor _44995_ (_22151_, _21978_, _02071_);
  nor _44996_ (_22152_, _21774_, _05587_);
  nor _44997_ (_22153_, _22123_, _22096_);
  and _44998_ (_22154_, _22153_, _22152_);
  nand _44999_ (_22155_, _22154_, _22151_);
  or _45000_ (_22156_, _22155_, _22150_);
  or _45001_ (_22157_, _21901_, _21790_);
  or _45002_ (_22158_, _21838_, _22157_);
  or _45003_ (_22159_, _21798_, _22158_);
  or _45004_ (_22160_, _22159_, _22156_);
  and _45005_ (_22161_, _22160_, _01760_);
  and _45006_ (_22162_, _02149_, _00000_);
  and _45007_ (_22163_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _45008_ (_22164_, _22163_, _22162_);
  or _45009_ (_22165_, _22164_, _22161_);
  and _45010_ (_05959_, _22165_, _25365_);
  or _45011_ (_22166_, _22147_, _22104_);
  or _45012_ (_22167_, _22166_, _22148_);
  or _45013_ (_22168_, _02094_, _02102_);
  or _45014_ (_22169_, _22168_, _02069_);
  or _45015_ (_22170_, _22090_, _21978_);
  or _45016_ (_22171_, _22170_, _22169_);
  or _45017_ (_22172_, _21843_, _22093_);
  or _45018_ (_22173_, _22172_, _22171_);
  or _45019_ (_22174_, _21859_, _22157_);
  or _45020_ (_22175_, _22174_, _22173_);
  or _45021_ (_22176_, _22175_, _22167_);
  and _45022_ (_22177_, _22176_, _01760_);
  and _45023_ (_22178_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _45024_ (_22179_, _02148_, _00000_);
  or _45025_ (_22180_, _22179_, _22178_);
  or _45026_ (_22181_, _22180_, _22177_);
  and _45027_ (_05960_, _22181_, _25365_);
  and _45028_ (_22182_, _21750_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _45029_ (_22183_, _22046_, _22006_);
  nor _45030_ (_22184_, _21964_, _22098_);
  nand _45031_ (_22185_, _22184_, _05589_);
  or _45032_ (_22186_, _22185_, _22183_);
  or _45033_ (_22187_, _21761_, _02064_);
  or _45034_ (_22188_, _22187_, _22095_);
  or _45035_ (_22189_, _22188_, _21883_);
  or _45036_ (_22190_, _22094_, _22092_);
  or _45037_ (_22191_, _22190_, _22189_);
  or _45038_ (_22192_, _22191_, _22186_);
  and _45039_ (_22193_, _22192_, _21651_);
  or _45040_ (_05961_, _22193_, _22182_);
  nor _45041_ (_06079_, _01823_, rst);
  nor _45042_ (_06080_, _05579_, rst);
  and _45043_ (_22194_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _45044_ (_22195_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _45045_ (_22196_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _45046_ (_22197_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _45047_ (_22198_, _22197_, _22196_);
  and _45048_ (_22199_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  not _45049_ (_22200_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _45050_ (_22201_, _01789_, _22200_);
  nor _45051_ (_22202_, _22201_, _22199_);
  and _45052_ (_22203_, _22202_, _22198_);
  and _45053_ (_22205_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _45054_ (_22206_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _45055_ (_22207_, _22206_, _22205_);
  and _45056_ (_22208_, _22207_, _22203_);
  nor _45057_ (_22209_, _22208_, _01767_);
  nor _45058_ (_22210_, _22209_, _22195_);
  nor _45059_ (_22211_, _22210_, _05562_);
  nor _45060_ (_22212_, _22211_, _22194_);
  nor _45061_ (_06081_, _22212_, rst);
  nor _45062_ (_06083_, _01872_, rst);
  and _45063_ (_06084_, _01898_, _25365_);
  and _45064_ (_06085_, _01920_, _25365_);
  nor _45065_ (_06086_, _01944_, rst);
  and _45066_ (_06087_, _01977_, _25365_);
  nor _45067_ (_06088_, _01798_, rst);
  nor _45068_ (_06089_, _01846_, rst);
  nor _45069_ (_06090_, _05669_, rst);
  nor _45070_ (_06091_, _05966_, rst);
  nor _45071_ (_06092_, _05891_, rst);
  nor _45072_ (_06093_, _05620_, rst);
  nor _45073_ (_06094_, _05745_, rst);
  nor _45074_ (_06096_, _05813_, rst);
  nor _45075_ (_06097_, _05863_, rst);
  and _45076_ (_22215_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _45077_ (_22216_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _45078_ (_22217_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _45079_ (_22218_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _45080_ (_22219_, _22218_, _22217_);
  and _45081_ (_22220_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  not _45082_ (_22221_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _45083_ (_22223_, _01789_, _22221_);
  nor _45084_ (_22224_, _22223_, _22220_);
  and _45085_ (_22225_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _45086_ (_22226_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _45087_ (_22227_, _22226_, _22225_);
  and _45088_ (_22228_, _22227_, _22224_);
  and _45089_ (_22229_, _22228_, _22219_);
  nor _45090_ (_22230_, _22229_, _01767_);
  nor _45091_ (_22231_, _22230_, _22216_);
  nor _45092_ (_22232_, _22231_, _05562_);
  nor _45093_ (_22234_, _22232_, _22215_);
  nor _45094_ (_06098_, _22234_, rst);
  and _45095_ (_22235_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _45096_ (_22236_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _45097_ (_22237_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _45098_ (_22238_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _45099_ (_22239_, _22238_, _22237_);
  and _45100_ (_22240_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _45101_ (_22241_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _45102_ (_22242_, _22241_, _22240_);
  and _45103_ (_22244_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  not _45104_ (_22245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _45105_ (_22246_, _01789_, _22245_);
  nor _45106_ (_22247_, _22246_, _22244_);
  and _45107_ (_22248_, _22247_, _22242_);
  and _45108_ (_22249_, _22248_, _22239_);
  nor _45109_ (_22250_, _22249_, _01767_);
  nor _45110_ (_22251_, _22250_, _22236_);
  nor _45111_ (_22252_, _22251_, _05562_);
  nor _45112_ (_22253_, _22252_, _22235_);
  nor _45113_ (_06099_, _22253_, rst);
  and _45114_ (_22255_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _45115_ (_22256_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _45116_ (_22257_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _45117_ (_22258_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _45118_ (_22259_, _22258_, _22257_);
  and _45119_ (_22260_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not _45120_ (_22261_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _45121_ (_22262_, _01789_, _22261_);
  nor _45122_ (_22263_, _22262_, _22260_);
  and _45123_ (_22264_, _22263_, _22259_);
  and _45124_ (_22265_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _45125_ (_22266_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _45126_ (_22267_, _22266_, _22265_);
  and _45127_ (_22268_, _22267_, _22264_);
  nor _45128_ (_22269_, _22268_, _01767_);
  nor _45129_ (_22270_, _22269_, _22256_);
  nor _45130_ (_22271_, _22270_, _05562_);
  nor _45131_ (_22272_, _22271_, _22255_);
  nor _45132_ (_06100_, _22272_, rst);
  and _45133_ (_22273_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _45134_ (_22274_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _45135_ (_22275_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _45136_ (_22276_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _45137_ (_22277_, _22276_, _22275_);
  and _45138_ (_22278_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _45139_ (_22279_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _45140_ (_22280_, _22279_, _22278_);
  and _45141_ (_22281_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not _45142_ (_22282_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _45143_ (_22283_, _01789_, _22282_);
  nor _45144_ (_22284_, _22283_, _22281_);
  and _45145_ (_22285_, _22284_, _22280_);
  and _45146_ (_22286_, _22285_, _22277_);
  nor _45147_ (_22287_, _22286_, _01767_);
  nor _45148_ (_22288_, _22287_, _22274_);
  nor _45149_ (_22289_, _22288_, _05562_);
  nor _45150_ (_22290_, _22289_, _22273_);
  nor _45151_ (_06101_, _22290_, rst);
  and _45152_ (_22291_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _45153_ (_22292_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _45154_ (_22293_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _45155_ (_22294_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _45156_ (_22295_, _22294_, _22293_);
  and _45157_ (_22296_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _45158_ (_22297_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _45159_ (_22298_, _22297_, _22296_);
  and _45160_ (_22299_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  not _45161_ (_22300_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _45162_ (_22301_, _01789_, _22300_);
  nor _45163_ (_22302_, _22301_, _22299_);
  and _45164_ (_22303_, _22302_, _22298_);
  and _45165_ (_22304_, _22303_, _22295_);
  nor _45166_ (_22305_, _22304_, _01767_);
  nor _45167_ (_22306_, _22305_, _22292_);
  nor _45168_ (_22307_, _22306_, _05562_);
  nor _45169_ (_22308_, _22307_, _22291_);
  nor _45170_ (_06102_, _22308_, rst);
  and _45171_ (_22309_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _45172_ (_22310_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _45173_ (_22311_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _45174_ (_22312_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _45175_ (_22313_, _22312_, _22311_);
  and _45176_ (_22314_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  not _45177_ (_22315_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _45178_ (_22316_, _01789_, _22315_);
  nor _45179_ (_22317_, _22316_, _22314_);
  and _45180_ (_22318_, _22317_, _22313_);
  and _45181_ (_22319_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _45182_ (_22320_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _45183_ (_22321_, _22320_, _22319_);
  and _45184_ (_22322_, _22321_, _22318_);
  nor _45185_ (_22323_, _22322_, _01767_);
  nor _45186_ (_22324_, _22323_, _22310_);
  nor _45187_ (_22325_, _22324_, _05562_);
  nor _45188_ (_22326_, _22325_, _22309_);
  nor _45189_ (_06103_, _22326_, rst);
  and _45190_ (_22327_, _05562_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _45191_ (_22328_, _01767_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _45192_ (_22329_, _01781_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _45193_ (_22330_, _01775_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _45194_ (_22331_, _22330_, _22329_);
  and _45195_ (_22332_, _01779_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  not _45196_ (_22333_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _45197_ (_22334_, _01789_, _22333_);
  nor _45198_ (_22335_, _22334_, _22332_);
  and _45199_ (_22336_, _01784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _45200_ (_22337_, _01771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _45201_ (_22338_, _22337_, _22336_);
  and _45202_ (_22339_, _22338_, _22335_);
  and _45203_ (_22340_, _22339_, _22331_);
  nor _45204_ (_22341_, _22340_, _01767_);
  nor _45205_ (_22342_, _22341_, _22328_);
  nor _45206_ (_22343_, _22342_, _05562_);
  nor _45207_ (_22344_, _22343_, _22327_);
  nor _45208_ (_06104_, _22344_, rst);
  and _45209_ (_22345_, _01761_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _45210_ (_22346_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _45211_ (_22347_, _22345_, _02402_);
  and _45212_ (_22348_, _22347_, _25365_);
  and _45213_ (_06107_, _22348_, _22346_);
  and _45214_ (_22349_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _45215_ (_22350_, _22345_);
  and _45216_ (_22351_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  or _45217_ (_22352_, _22351_, _22349_);
  and _45218_ (_06108_, _22352_, _25365_);
  nor _45219_ (_06113_, _05584_, rst);
  and _45220_ (_06115_, _05559_, _25365_);
  or _45221_ (_22353_, _05597_, _02036_);
  not _45222_ (_22354_, _22353_);
  nor _45223_ (_22355_, _22354_, _05599_);
  not _45224_ (_22356_, _22355_);
  nor _45225_ (_22357_, _05653_, _00921_);
  and _45226_ (_22358_, _05653_, _00921_);
  nor _45227_ (_22359_, _22358_, _22357_);
  nor _45228_ (_22360_, _05775_, _00938_);
  and _45229_ (_22361_, _05775_, _00938_);
  nor _45230_ (_22362_, _22361_, _22360_);
  or _45231_ (_22363_, _22362_, _22359_);
  nor _45232_ (_22364_, _05821_, _00892_);
  and _45233_ (_22365_, _05821_, _00892_);
  nor _45234_ (_22366_, _22365_, _22364_);
  nor _45235_ (_22367_, _05867_, _00879_);
  and _45236_ (_22368_, _05867_, _00879_);
  nor _45237_ (_22369_, _22368_, _22367_);
  or _45238_ (_22370_, _22369_, _22366_);
  or _45239_ (_22371_, _22370_, _22363_);
  nor _45240_ (_22372_, _22371_, _06012_);
  nor _45241_ (_22373_, _01294_, _03341_);
  and _45242_ (_22374_, _22373_, _22372_);
  and _45243_ (_22375_, _22374_, _22356_);
  not _45244_ (_22376_, _22375_);
  nor _45245_ (_22377_, _05918_, _00835_);
  and _45246_ (_22378_, _05918_, _00835_);
  nor _45247_ (_22379_, _22378_, _22377_);
  and _45248_ (_22380_, _05720_, _01405_);
  nor _45249_ (_22381_, _22380_, _22379_);
  nor _45250_ (_22382_, _05994_, _00847_);
  and _45251_ (_22383_, _05994_, _00847_);
  nor _45252_ (_22384_, _22383_, _22382_);
  nor _45253_ (_22385_, _05720_, _01405_);
  nor _45254_ (_22386_, _22385_, _22384_);
  and _45255_ (_22387_, _22386_, _22381_);
  and _45256_ (_22388_, _22387_, _01189_);
  and _45257_ (_22389_, _22388_, _22372_);
  nor _45258_ (_22390_, _00906_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _45259_ (_22391_, _22390_, _22389_);
  not _45260_ (_22392_, _22391_);
  nor _45261_ (_22393_, _21814_, _02140_);
  nor _45262_ (_22394_, _02084_, _02079_);
  nor _45263_ (_22395_, _21760_, _02111_);
  and _45264_ (_22396_, _22356_, _00997_);
  not _45265_ (_22397_, _22396_);
  and _45266_ (_22398_, _22355_, _02146_);
  or _45267_ (_22399_, _01081_, _01060_);
  or _45268_ (_22400_, _22399_, _01306_);
  nor _45269_ (_22401_, _22400_, _01075_);
  nand _45270_ (_22402_, _22401_, _01427_);
  nor _45271_ (_22403_, _22402_, _01548_);
  and _45272_ (_22404_, _22403_, _01613_);
  and _45273_ (_22405_, _22404_, _22398_);
  and _45274_ (_22406_, _22405_, _01099_);
  and _45275_ (_22407_, _02081_, _01999_);
  and _45276_ (_22408_, _22407_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _45277_ (_22409_, _22408_, _22406_);
  and _45278_ (_22410_, _01998_, _01994_);
  and _45279_ (_22411_, _22410_, _02079_);
  nor _45280_ (_22412_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _45281_ (_22413_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _45282_ (_22414_, _22413_, _22412_);
  nor _45283_ (_22415_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _45284_ (_22416_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _45285_ (_22417_, _22416_, _22415_);
  and _45286_ (_22418_, _22417_, _22414_);
  nand _45287_ (_22419_, _22418_, _22411_);
  and _45288_ (_22420_, _22419_, _22409_);
  and _45289_ (_22421_, _22420_, _22397_);
  not _45290_ (_22422_, _22006_);
  not _45291_ (_22423_, _21841_);
  nor _45292_ (_22424_, _22046_, _02042_);
  and _45293_ (_22425_, _22424_, _22423_);
  and _45294_ (_22426_, _22425_, _22422_);
  not _45295_ (_22427_, _02066_);
  nor _45296_ (_22428_, _02058_, _02027_);
  and _45297_ (_22429_, _22428_, _22427_);
  nor _45298_ (_22430_, _22429_, _02029_);
  not _45299_ (_22431_, _22430_);
  and _45300_ (_22432_, _22431_, _22426_);
  not _45301_ (_22433_, _22432_);
  and _45302_ (_22434_, _22433_, _22421_);
  nand _45303_ (_22435_, _02080_, _01987_);
  and _45304_ (_22436_, _22435_, _02031_);
  and _45305_ (_22437_, _22436_, _02035_);
  nor _45306_ (_22438_, _22437_, _22421_);
  nor _45307_ (_22439_, _22438_, _22434_);
  nand _45308_ (_22440_, _22439_, _22395_);
  nor _45309_ (_22441_, _22440_, _02126_);
  nor _45310_ (_22442_, _22441_, _22394_);
  nor _45311_ (_22443_, _22442_, _22393_);
  not _45312_ (_22444_, _02851_);
  and _45313_ (_22445_, _22444_, _02093_);
  and _45314_ (_22446_, _22355_, _01803_);
  nor _45315_ (_22447_, _22446_, _02146_);
  nor _45316_ (_22448_, _02684_, _02675_);
  and _45317_ (_22449_, _22448_, _02726_);
  not _45318_ (_22450_, _22449_);
  and _45319_ (_22451_, _22450_, _22447_);
  nor _45320_ (_22452_, _22451_, _22445_);
  not _45321_ (_22453_, _22452_);
  nor _45322_ (_22454_, _22453_, _22443_);
  and _45323_ (_22455_, _22454_, _22392_);
  and _45324_ (_22456_, _22455_, _22376_);
  nor _45325_ (_22457_, _02084_, rst);
  and _45326_ (_06118_, _22457_, _22456_);
  and _45327_ (_06119_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _25365_);
  and _45328_ (_06120_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _25365_);
  nor _45329_ (_22458_, _01770_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _45330_ (_22459_, _22458_, _05562_);
  nor _45331_ (_22460_, _22459_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _45332_ (_22461_, _22460_);
  and _45333_ (_22462_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _45334_ (_22463_, _22462_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _45335_ (_22464_, _22463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _45336_ (_22465_, _22464_, _22461_);
  and _45337_ (_22466_, _22465_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _45338_ (_22467_, _22466_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _45339_ (_22468_, _22467_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _45340_ (_22469_, _22468_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _45341_ (_22470_, _22469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _45342_ (_22471_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _45343_ (_22472_, _22471_, _22470_);
  and _45344_ (_22473_, _22472_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _45345_ (_22474_, _22473_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _45346_ (_22475_, _22474_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _45347_ (_22476_, _22474_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _45348_ (_22477_, _22476_, _22475_);
  or _45349_ (_22478_, _22477_, _22456_);
  and _45350_ (_22479_, _22478_, _25365_);
  and _45351_ (_22480_, _01998_, _01852_);
  nand _45352_ (_22481_, _22480_, _01756_);
  and _45353_ (_22482_, _22481_, _22353_);
  or _45354_ (_22483_, _22183_, _02042_);
  nand _45355_ (_22484_, _22483_, _02079_);
  and _45356_ (_22485_, _21813_, _01756_);
  nor _45357_ (_22486_, _22485_, _02084_);
  and _45358_ (_22487_, _22486_, _22484_);
  and _45359_ (_22488_, _22487_, _22482_);
  and _45360_ (_22489_, _22488_, _05579_);
  nand _45361_ (_22490_, _22487_, _22482_);
  and _45362_ (_22491_, _22490_, _22212_);
  nor _45363_ (_22492_, _22491_, _22489_);
  and _45364_ (_22493_, _22492_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _45365_ (_22494_, _22492_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _45366_ (_22495_, _22494_);
  and _45367_ (_22496_, _22488_, _05863_);
  and _45368_ (_22497_, _22490_, _22344_);
  nor _45369_ (_22498_, _22497_, _22496_);
  and _45370_ (_22499_, _22498_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _45371_ (_22500_, _22499_);
  nor _45372_ (_22501_, _22498_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _45373_ (_22502_, _22501_, _22499_);
  and _45374_ (_22503_, _22488_, _05813_);
  and _45375_ (_22504_, _22490_, _22326_);
  nor _45376_ (_22505_, _22504_, _22503_);
  nor _45377_ (_22506_, _22505_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _45378_ (_22507_, _22505_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _45379_ (_22508_, _22488_, _05745_);
  and _45380_ (_22509_, _22490_, _22308_);
  nor _45381_ (_22510_, _22509_, _22508_);
  nand _45382_ (_22511_, _22510_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _45383_ (_22512_, _22488_, _05620_);
  and _45384_ (_22513_, _22490_, _22290_);
  nor _45385_ (_22514_, _22513_, _22512_);
  nor _45386_ (_22515_, _22514_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _45387_ (_22516_, _22514_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _45388_ (_22517_, _22490_, _05892_);
  not _45389_ (_22518_, _22272_);
  or _45390_ (_22519_, _22488_, _22518_);
  nand _45391_ (_22520_, _22519_, _22517_);
  or _45392_ (_22521_, _22520_, _00317_);
  or _45393_ (_22522_, _22490_, _05967_);
  not _45394_ (_22523_, _22253_);
  or _45395_ (_22524_, _22488_, _22523_);
  and _45396_ (_22525_, _22524_, _22522_);
  nand _45397_ (_22526_, _22525_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _45398_ (_22527_, _22490_, _05670_);
  not _45399_ (_22528_, _22234_);
  or _45400_ (_22529_, _22488_, _22528_);
  and _45401_ (_22530_, _22529_, _22527_);
  and _45402_ (_22531_, _22530_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _45403_ (_22532_, _22525_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _45404_ (_22533_, _22532_, _22526_);
  and _45405_ (_22534_, _22533_, _22531_);
  not _45406_ (_22535_, _22534_);
  nand _45407_ (_22536_, _22535_, _22526_);
  nand _45408_ (_22537_, _22520_, _00317_);
  and _45409_ (_22538_, _22537_, _22521_);
  and _45410_ (_22539_, _22538_, _22536_);
  not _45411_ (_22540_, _22539_);
  nand _45412_ (_22541_, _22540_, _22521_);
  nor _45413_ (_22542_, _22541_, _22516_);
  nor _45414_ (_22543_, _22542_, _22515_);
  or _45415_ (_22544_, _22510_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _45416_ (_22545_, _22544_, _22511_);
  nand _45417_ (_22546_, _22545_, _22543_);
  nand _45418_ (_22547_, _22546_, _22511_);
  nor _45419_ (_22548_, _22547_, _22507_);
  nor _45420_ (_22549_, _22548_, _22506_);
  nand _45421_ (_22550_, _22549_, _22502_);
  nand _45422_ (_22551_, _22550_, _22500_);
  and _45423_ (_22552_, _22551_, _22495_);
  or _45424_ (_22553_, _22552_, _22493_);
  and _45425_ (_22554_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _45426_ (_22555_, _22554_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _45427_ (_22556_, _22555_, _22553_);
  and _45428_ (_22557_, _22556_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _45429_ (_22558_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _45430_ (_22559_, _22558_, _22557_);
  or _45431_ (_22560_, _22559_, _22492_);
  not _45432_ (_22561_, _22492_);
  or _45433_ (_22562_, _22553_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _45434_ (_22563_, _22562_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _45435_ (_22564_, _22563_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _45436_ (_22565_, _22564_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _45437_ (_22566_, _22565_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _45438_ (_22567_, _22566_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _45439_ (_22568_, _22567_, _22561_);
  and _45440_ (_22569_, _22568_, _22560_);
  or _45441_ (_22570_, _22492_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _45442_ (_22571_, _22492_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _45443_ (_22572_, _22571_, _22570_);
  and _45444_ (_22573_, _22572_, _22569_);
  nand _45445_ (_22574_, _22573_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _45446_ (_22575_, _22573_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _45447_ (_22576_, _22395_, _22426_);
  and _45448_ (_22577_, _22576_, _02079_);
  not _45449_ (_22578_, _22577_);
  and _45450_ (_22579_, _22482_, _02146_);
  and _45451_ (_22580_, _22579_, _22578_);
  and _45452_ (_22581_, _02111_, _02079_);
  nor _45453_ (_22582_, _22581_, _22393_);
  not _45454_ (_22583_, _22582_);
  and _45455_ (_22584_, _22583_, _22488_);
  nor _45456_ (_22585_, _22584_, _22580_);
  and _45457_ (_22586_, _22585_, _22575_);
  and _45458_ (_22587_, _22586_, _22574_);
  and _45459_ (_22588_, _02084_, _01184_);
  and _45460_ (_22589_, _22581_, _02413_);
  and _45461_ (_22590_, _22582_, _22488_);
  and _45462_ (_22591_, _22590_, _22580_);
  and _45463_ (_22592_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _45464_ (_22593_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _45465_ (_22594_, _22593_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _45466_ (_22595_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _45467_ (_22596_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _45468_ (_22597_, _22596_, _22595_);
  and _45469_ (_22598_, _22597_, _22594_);
  and _45470_ (_22599_, _22598_, _22555_);
  and _45471_ (_22600_, _22599_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _45472_ (_22601_, _22600_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _45473_ (_22602_, _22601_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _45474_ (_22603_, _22602_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _45475_ (_22604_, _22603_, _02402_);
  or _45476_ (_22605_, _22603_, _02402_);
  and _45477_ (_22606_, _22605_, _22604_);
  and _45478_ (_22607_, _22584_, _22580_);
  and _45479_ (_22608_, _22607_, _22606_);
  and _45480_ (_22609_, _22485_, _05580_);
  or _45481_ (_22610_, _22609_, _22608_);
  or _45482_ (_22611_, _22610_, _22592_);
  nor _45483_ (_22612_, _22611_, _22589_);
  nand _45484_ (_22613_, _22612_, _22456_);
  or _45485_ (_22614_, _22613_, _22588_);
  or _45486_ (_22615_, _22614_, _22587_);
  and _45487_ (_06121_, _22615_, _22479_);
  not _45488_ (_22616_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _45489_ (_22617_, _01760_, _22616_);
  not _45490_ (_22618_, _22617_);
  not _45491_ (_22619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _45492_ (_22620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _45493_ (_22621_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _45494_ (_22622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _45495_ (_22623_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _45496_ (_22624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _45497_ (_22625_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _45498_ (_22626_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45499_ (_22627_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _45500_ (_22628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _45501_ (_22629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _45502_ (_22630_, _22629_, _22627_);
  and _45503_ (_22631_, _22630_, _22628_);
  nor _45504_ (_22632_, _22631_, _22627_);
  nor _45505_ (_22633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _45506_ (_22634_, _22633_, _22626_);
  not _45507_ (_22635_, _22634_);
  nor _45508_ (_22636_, _22635_, _22632_);
  nor _45509_ (_22637_, _22636_, _22626_);
  not _45510_ (_22638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _45511_ (_22639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _45512_ (_22640_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _45513_ (_22641_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _45514_ (_22642_, _22641_, _22640_);
  and _45515_ (_22643_, _22642_, _22639_);
  and _45516_ (_22644_, _22643_, _22638_);
  and _45517_ (_22645_, _22644_, _22637_);
  and _45518_ (_22646_, _22645_, _22625_);
  and _45519_ (_22647_, _22646_, _22624_);
  and _45520_ (_22648_, _22647_, _22623_);
  and _45521_ (_22649_, _22648_, _22622_);
  and _45522_ (_22650_, _22649_, _22621_);
  and _45523_ (_22651_, _22650_, _22620_);
  and _45524_ (_22652_, _22651_, _22619_);
  nor _45525_ (_22653_, _22651_, _22619_);
  nor _45526_ (_22654_, _22653_, _22652_);
  not _45527_ (_22655_, _22654_);
  nor _45528_ (_22656_, _22650_, _22620_);
  nor _45529_ (_22657_, _22656_, _22651_);
  not _45530_ (_22658_, _22657_);
  nor _45531_ (_22659_, _22649_, _22621_);
  nor _45532_ (_22660_, _22659_, _22650_);
  not _45533_ (_22661_, _22660_);
  nor _45534_ (_22662_, _22648_, _22622_);
  nor _45535_ (_22663_, _22662_, _22649_);
  not _45536_ (_22664_, _22663_);
  nor _45537_ (_22665_, _22647_, _22623_);
  or _45538_ (_22666_, _22665_, _22648_);
  nor _45539_ (_22667_, _22646_, _22624_);
  nor _45540_ (_22668_, _22667_, _22647_);
  not _45541_ (_22669_, _22668_);
  and _45542_ (_22670_, _22637_, _22643_);
  nor _45543_ (_22671_, _22670_, _22638_);
  nor _45544_ (_22672_, _22671_, _22645_);
  not _45545_ (_22673_, _22672_);
  and _45546_ (_22674_, _22637_, _22642_);
  nor _45547_ (_22675_, _22674_, _22639_);
  nor _45548_ (_22676_, _22675_, _22670_);
  not _45549_ (_22677_, _22676_);
  and _45550_ (_22678_, _22637_, _22641_);
  nor _45551_ (_22679_, _22678_, _22640_);
  nor _45552_ (_22680_, _22679_, _22674_);
  not _45553_ (_22681_, _22680_);
  not _45554_ (_22682_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _45555_ (_22683_, _22637_, _22682_);
  nor _45556_ (_22684_, _22637_, _22682_);
  nor _45557_ (_22685_, _22684_, _22683_);
  not _45558_ (_22686_, _22685_);
  and _45559_ (_22687_, _21685_, _21723_);
  not _45560_ (_22688_, _21729_);
  nor _45561_ (_22689_, _21686_, _21668_);
  nor _45562_ (_22690_, _22689_, _22688_);
  nor _45563_ (_22691_, _22690_, _22687_);
  and _45564_ (_22692_, _21710_, _21655_);
  and _45565_ (_22693_, _22692_, _21660_);
  nor _45566_ (_22694_, _21665_, _21659_);
  not _45567_ (_22695_, _22694_);
  and _45568_ (_22696_, _21704_, _01872_);
  and _45569_ (_22697_, _22696_, _22695_);
  nor _45570_ (_22698_, _22697_, _22693_);
  and _45571_ (_22699_, _22698_, _22691_);
  and _45572_ (_22700_, _21704_, _21683_);
  nor _45573_ (_22701_, _21708_, _21723_);
  nor _45574_ (_22702_, _22701_, _22688_);
  nor _45575_ (_22703_, _22702_, _22700_);
  and _45576_ (_22704_, _22695_, _21696_);
  not _45577_ (_22705_, _21660_);
  nor _45578_ (_22706_, _21708_, _21701_);
  nor _45579_ (_22707_, _22706_, _22705_);
  nor _45580_ (_22708_, _22707_, _22704_);
  and _45581_ (_22709_, _22708_, _22703_);
  and _45582_ (_22710_, _22709_, _22699_);
  not _45583_ (_22711_, _21707_);
  nor _45584_ (_22712_, _21685_, _21659_);
  and _45585_ (_22713_, _21695_, _21710_);
  not _45586_ (_22714_, _21685_);
  nor _45587_ (_22715_, _21708_, _21728_);
  nor _45588_ (_22716_, _22715_, _22714_);
  nor _45589_ (_22717_, _22716_, _22713_);
  nor _45590_ (_22718_, _22717_, _22712_);
  nor _45591_ (_22719_, _22718_, _22711_);
  and _45592_ (_22720_, _22719_, _22710_);
  nor _45593_ (_22721_, _21730_, _21714_);
  nand _45594_ (_22722_, _21676_, _21682_);
  and _45595_ (_22723_, _21675_, _21660_);
  and _45596_ (_22724_, _22713_, _21683_);
  nor _45597_ (_22725_, _22724_, _22723_);
  and _45598_ (_22726_, _22725_, _22722_);
  and _45599_ (_22727_, _22726_, _22721_);
  and _45600_ (_22728_, _21712_, _21660_);
  and _45601_ (_22729_, _21666_, _21655_);
  or _45602_ (_22730_, _22692_, _22729_);
  not _45603_ (_22731_, _22730_);
  and _45604_ (_22732_, _21667_, _21703_);
  nor _45605_ (_22733_, _22732_, _21675_);
  and _45606_ (_22734_, _22733_, _22731_);
  nor _45607_ (_22735_, _22734_, _22714_);
  nor _45608_ (_22736_, _22735_, _22728_);
  and _45609_ (_22737_, _21700_, _21655_);
  and _45610_ (_22738_, _22737_, _01977_);
  nor _45611_ (_22739_, _22732_, _22692_);
  nor _45612_ (_22740_, _21704_, _21677_);
  and _45613_ (_22741_, _22740_, _22739_);
  nor _45614_ (_22742_, _22741_, _22688_);
  nor _45615_ (_22743_, _22742_, _22738_);
  and _45616_ (_22744_, _22743_, _22736_);
  nor _45617_ (_22745_, _21735_, _21724_);
  nor _45618_ (_22746_, _21671_, _22729_);
  not _45619_ (_22747_, _22746_);
  and _45620_ (_22748_, _22747_, _21700_);
  and _45621_ (_22749_, _21655_, _21656_);
  nor _45622_ (_22750_, _22749_, _21708_);
  nor _45623_ (_22751_, _22750_, _01944_);
  nor _45624_ (_22752_, _22751_, _22748_);
  and _45625_ (_22753_, _22752_, _22745_);
  and _45626_ (_22754_, _21658_, _01898_);
  and _45627_ (_22755_, _22754_, _22749_);
  not _45628_ (_22756_, _22755_);
  and _45629_ (_22757_, _21695_, _21716_);
  and _45630_ (_22758_, _21733_, _22757_);
  nor _45631_ (_22759_, _22758_, _21672_);
  and _45632_ (_22760_, _22759_, _22756_);
  nor _45633_ (_22761_, _21726_, _21688_);
  and _45634_ (_22762_, _22761_, _22760_);
  and _45635_ (_22763_, _22762_, _22753_);
  and _45636_ (_22764_, _22763_, _22744_);
  and _45637_ (_22765_, _22764_, _22727_);
  and _45638_ (_22766_, _22765_, _22720_);
  not _45639_ (_22767_, _22766_);
  nor _45640_ (_22768_, _22630_, _22628_);
  nor _45641_ (_22769_, _22768_, _22631_);
  nand _45642_ (_22770_, _22769_, _22767_);
  or _45643_ (_22771_, _21735_, _21688_);
  or _45644_ (_22772_, _22771_, _22702_);
  or _45645_ (_22773_, _22700_, _21702_);
  and _45646_ (_22774_, _21696_, _21683_);
  and _45647_ (_22775_, _21700_, _22692_);
  or _45648_ (_22776_, _22775_, _22774_);
  or _45649_ (_22777_, _22776_, _22773_);
  nor _45650_ (_22778_, _22777_, _22772_);
  nand _45651_ (_22779_, _22778_, _22727_);
  nor _45652_ (_22780_, _22779_, _22766_);
  not _45653_ (_22781_, _22780_);
  nor _45654_ (_22782_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _45655_ (_22783_, _22782_, _22628_);
  and _45656_ (_22784_, _22783_, _22781_);
  or _45657_ (_22785_, _22769_, _22767_);
  and _45658_ (_22786_, _22785_, _22770_);
  nand _45659_ (_22787_, _22786_, _22784_);
  and _45660_ (_22788_, _22787_, _22770_);
  not _45661_ (_22789_, _22788_);
  and _45662_ (_22790_, _22635_, _22632_);
  nor _45663_ (_22791_, _22790_, _22636_);
  and _45664_ (_22792_, _22791_, _22789_);
  and _45665_ (_22793_, _22792_, _22686_);
  not _45666_ (_22794_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _45667_ (_22795_, _22683_, _22794_);
  or _45668_ (_22796_, _22795_, _22678_);
  and _45669_ (_22797_, _22796_, _22793_);
  and _45670_ (_22798_, _22797_, _22681_);
  and _45671_ (_22799_, _22798_, _22677_);
  and _45672_ (_22800_, _22799_, _22673_);
  nor _45673_ (_22801_, _22645_, _22625_);
  or _45674_ (_22802_, _22801_, _22646_);
  and _45675_ (_22803_, _22802_, _22800_);
  and _45676_ (_22804_, _22803_, _22669_);
  and _45677_ (_22805_, _22804_, _22666_);
  and _45678_ (_22806_, _22805_, _22664_);
  and _45679_ (_22807_, _22806_, _22661_);
  and _45680_ (_22808_, _22807_, _22658_);
  and _45681_ (_22809_, _22808_, _22655_);
  nor _45682_ (_22810_, _22809_, _22618_);
  nor _45683_ (_22811_, _22617_, _02402_);
  not _45684_ (_22812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _45685_ (_22813_, _22652_, _22812_);
  nor _45686_ (_22814_, _22652_, _22812_);
  nor _45687_ (_22815_, _22814_, _22813_);
  and _45688_ (_22816_, _22815_, _22617_);
  or _45689_ (_22817_, _22816_, _22811_);
  or _45690_ (_22818_, _22817_, _22810_);
  nand _45691_ (_22819_, _22815_, _22810_);
  nor _45692_ (_22820_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _45693_ (_22821_, _22820_, _22819_);
  and _45694_ (_22822_, _22821_, _22818_);
  and _45695_ (_22823_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _25365_);
  and _45696_ (_22824_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _45697_ (_06122_, _22824_, _22822_);
  nor _45698_ (_22825_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _45699_ (_06123_, _22825_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _45700_ (_06124_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _25365_);
  nor _45701_ (_22826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _45702_ (_22827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _45703_ (_22828_, _22827_, _22826_);
  nor _45704_ (_22829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _45705_ (_22830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _45706_ (_22831_, _22830_, _22829_);
  and _45707_ (_22832_, _22831_, _22828_);
  nor _45708_ (_22833_, _22832_, rst);
  and _45709_ (_22834_, \oc8051_top_1.oc8051_rom1.ea_int , _01757_);
  nand _45710_ (_22835_, _22834_, _01760_);
  and _45711_ (_22836_, _22835_, _06124_);
  or _45712_ (_06125_, _22836_, _22833_);
  and _45713_ (_22837_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _45714_ (_22838_, _22837_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _45715_ (_06126_, _22838_, _25365_);
  nor _45716_ (_22839_, _22460_, _05562_);
  or _45717_ (_22840_, _22766_, _01773_);
  nor _45718_ (_22841_, _22780_, _01787_);
  nand _45719_ (_22842_, _22766_, _01773_);
  and _45720_ (_22843_, _22842_, _22840_);
  nand _45721_ (_22844_, _22843_, _22841_);
  and _45722_ (_22845_, _22844_, _22840_);
  nor _45723_ (_22846_, _22845_, _05562_);
  and _45724_ (_22847_, _22846_, _01769_);
  nor _45725_ (_22848_, _22846_, _01769_);
  nor _45726_ (_22849_, _22848_, _22847_);
  nor _45727_ (_22850_, _22849_, _22839_);
  and _45728_ (_22851_, _01774_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45729_ (_22852_, _22851_, _22839_);
  and _45730_ (_22853_, _22852_, _22779_);
  or _45731_ (_22854_, _22853_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _45732_ (_22855_, _22854_, _22850_);
  and _45733_ (_06127_, _22855_, _25365_);
  and _45734_ (_22856_, _01891_, _01818_);
  and _45735_ (_22857_, _01970_, _01842_);
  and _45736_ (_22858_, _22857_, _22856_);
  and _45737_ (_22859_, _01761_, _25365_);
  and _45738_ (_22860_, _22859_, _01916_);
  and _45739_ (_22861_, _22860_, _01939_);
  and _45740_ (_22862_, _01868_, _01794_);
  and _45741_ (_22863_, _22862_, _22861_);
  and _45742_ (_06130_, _22863_, _22858_);
  nor _45743_ (_22864_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _45744_ (_22865_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _45745_ (_22866_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _45746_ (_06132_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _25365_);
  and _45747_ (_22867_, _06132_, _22866_);
  or _45748_ (_06131_, _22867_, _22865_);
  not _45749_ (_22868_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _45750_ (_22869_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _45751_ (_22870_, _22869_, _22868_);
  and _45752_ (_22871_, _22869_, _22868_);
  nor _45753_ (_22872_, _22871_, _22870_);
  not _45754_ (_22873_, _22872_);
  and _45755_ (_22874_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _45756_ (_22875_, _22874_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _45757_ (_22876_, _22874_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _45758_ (_22877_, _22876_, _22875_);
  or _45759_ (_22878_, _22877_, _22869_);
  and _45760_ (_22879_, _22878_, _22873_);
  nor _45761_ (_22880_, _22870_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _45762_ (_22881_, _22870_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _45763_ (_22882_, _22881_, _22880_);
  or _45764_ (_22883_, _22875_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _45765_ (_06135_, _22883_, _25365_);
  and _45766_ (_22884_, _06135_, _22882_);
  and _45767_ (_06134_, _22884_, _22879_);
  not _45768_ (_22885_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _45769_ (_22886_, _22460_, _22885_);
  and _45770_ (_22887_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _45771_ (_22888_, _22886_);
  and _45772_ (_22889_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _45773_ (_22890_, _22889_, _22887_);
  and _45774_ (_06136_, _22890_, _25365_);
  and _45775_ (_22891_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor _45776_ (_22892_, _22886_, _05565_);
  or _45777_ (_22893_, _22892_, _22891_);
  and _45778_ (_06137_, _22893_, _25365_);
  and _45779_ (_22894_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _45780_ (_22895_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _45781_ (_22896_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _22895_);
  and _45782_ (_22897_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _45783_ (_22898_, _22897_, _22894_);
  and _45784_ (_06138_, _22898_, _25365_);
  and _45785_ (_22899_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  or _45786_ (_22900_, _22899_, _22896_);
  and _45787_ (_06139_, _22900_, _25365_);
  or _45788_ (_22901_, _22895_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _45789_ (_06140_, _22901_, _25365_);
  not _45790_ (_22902_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _45791_ (_22903_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _45792_ (_22904_, _22903_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _45793_ (_22905_, _22895_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _45794_ (_22906_, _22905_, _25365_);
  and _45795_ (_06141_, _22906_, _22904_);
  or _45796_ (_22907_, _22895_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _45797_ (_06142_, _22907_, _25365_);
  nor _45798_ (_22908_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _45799_ (_22909_, _22908_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _45800_ (_22910_, _22909_, _25365_);
  and _45801_ (_22911_, _06132_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _45802_ (_06143_, _22911_, _22910_);
  and _45803_ (_22912_, _22885_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _45804_ (_22913_, _22912_, _22909_);
  and _45805_ (_06144_, _22913_, _25365_);
  not _45806_ (_22914_, _22909_);
  or _45807_ (_22915_, _22914_, _02413_);
  or _45808_ (_22916_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _45809_ (_22917_, _22916_, _25365_);
  and _45810_ (_06145_, _22917_, _22915_);
  or _45811_ (_22918_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand _45812_ (_22919_, _22345_, _00349_);
  and _45813_ (_22920_, _22919_, _25365_);
  and _45814_ (_06150_, _22920_, _22918_);
  or _45815_ (_22921_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _45816_ (_22922_, _22345_, _00299_);
  and _45817_ (_22923_, _22922_, _25365_);
  and _45818_ (_06151_, _22923_, _22921_);
  or _45819_ (_22924_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _45820_ (_22925_, _22345_, _00317_);
  and _45821_ (_22926_, _22925_, _25365_);
  and _45822_ (_06152_, _22926_, _22924_);
  or _45823_ (_22927_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _45824_ (_22928_, _22345_, _00202_);
  and _45825_ (_22929_, _22928_, _25365_);
  and _45826_ (_06154_, _22929_, _22927_);
  or _45827_ (_22930_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand _45828_ (_22931_, _22345_, _00031_);
  and _45829_ (_22932_, _22931_, _25365_);
  and _45830_ (_06155_, _22932_, _22930_);
  or _45831_ (_22933_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _45832_ (_22934_, _22345_, _00220_);
  and _45833_ (_22935_, _22934_, _25365_);
  and _45834_ (_06156_, _22935_, _22933_);
  or _45835_ (_22936_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _45836_ (_22937_, _22345_, _00241_);
  and _45837_ (_22938_, _22937_, _25365_);
  and _45838_ (_06157_, _22938_, _22936_);
  or _45839_ (_22939_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand _45840_ (_22940_, _22345_, _00271_);
  and _45841_ (_22941_, _22940_, _25365_);
  and _45842_ (_06158_, _22941_, _22939_);
  or _45843_ (_22942_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _45844_ (_22943_, _22345_, _02374_);
  and _45845_ (_22944_, _22943_, _25365_);
  and _45846_ (_06159_, _22944_, _22942_);
  or _45847_ (_22945_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _45848_ (_22946_, _22345_, _02380_);
  and _45849_ (_22947_, _22946_, _25365_);
  and _45850_ (_06160_, _22947_, _22945_);
  or _45851_ (_22948_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _45852_ (_22949_, _22345_, _02385_);
  and _45853_ (_22950_, _22949_, _25365_);
  and _45854_ (_06161_, _22950_, _22948_);
  or _45855_ (_22951_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _45856_ (_22952_, _22345_, _02370_);
  and _45857_ (_22953_, _22952_, _25365_);
  and _45858_ (_06162_, _22953_, _22951_);
  or _45859_ (_22954_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _45860_ (_22955_, _22345_, _02391_);
  and _45861_ (_22956_, _22955_, _25365_);
  and _45862_ (_06163_, _22956_, _22954_);
  or _45863_ (_22957_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _45864_ (_22958_, _22345_, _02366_);
  and _45865_ (_22959_, _22958_, _25365_);
  and _45866_ (_06164_, _22959_, _22957_);
  or _45867_ (_22960_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _45868_ (_22961_, _22345_, _02397_);
  and _45869_ (_22962_, _22961_, _25365_);
  and _45870_ (_06165_, _22962_, _22960_);
  and _45871_ (_22963_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _45872_ (_22964_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _45873_ (_22965_, _22964_, _22963_);
  and _45874_ (_06166_, _22965_, _25365_);
  and _45875_ (_22966_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _45876_ (_22967_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _45877_ (_22968_, _22967_, _22966_);
  and _45878_ (_06167_, _22968_, _25365_);
  and _45879_ (_22969_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _45880_ (_22970_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _45881_ (_22971_, _22970_, _22969_);
  and _45882_ (_06168_, _22971_, _25365_);
  and _45883_ (_22972_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _45884_ (_22973_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _45885_ (_22974_, _22973_, _22972_);
  and _45886_ (_06169_, _22974_, _25365_);
  and _45887_ (_22975_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _45888_ (_22976_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or _45889_ (_22977_, _22976_, _22975_);
  and _45890_ (_06170_, _22977_, _25365_);
  and _45891_ (_22978_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _45892_ (_22979_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or _45893_ (_22980_, _22979_, _22978_);
  and _45894_ (_06171_, _22980_, _25365_);
  and _45895_ (_22981_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _45896_ (_22982_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or _45897_ (_22983_, _22982_, _22981_);
  and _45898_ (_06172_, _22983_, _25365_);
  and _45899_ (_22984_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _45900_ (_22985_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or _45901_ (_22986_, _22985_, _22984_);
  and _45902_ (_06173_, _22986_, _25365_);
  and _45903_ (_22987_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _45904_ (_22988_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or _45905_ (_22989_, _22988_, _22987_);
  and _45906_ (_06174_, _22989_, _25365_);
  and _45907_ (_22990_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _45908_ (_22991_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _45909_ (_22992_, _22991_, _22990_);
  and _45910_ (_06175_, _22992_, _25365_);
  and _45911_ (_22993_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _45912_ (_22994_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or _45913_ (_22995_, _22994_, _22993_);
  and _45914_ (_06176_, _22995_, _25365_);
  and _45915_ (_22996_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _45916_ (_22997_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or _45917_ (_22998_, _22997_, _22996_);
  and _45918_ (_06177_, _22998_, _25365_);
  and _45919_ (_22999_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _45920_ (_23000_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or _45921_ (_23001_, _23000_, _22999_);
  and _45922_ (_06178_, _23001_, _25365_);
  and _45923_ (_23002_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _45924_ (_23003_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or _45925_ (_23004_, _23003_, _23002_);
  and _45926_ (_06179_, _23004_, _25365_);
  and _45927_ (_23005_, _22345_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _45928_ (_23006_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or _45929_ (_23007_, _23006_, _23005_);
  and _45930_ (_06180_, _23007_, _25365_);
  and _45931_ (_06200_, _01876_, _25365_);
  and _45932_ (_06201_, _01902_, _25365_);
  and _45933_ (_06202_, _01924_, _25365_);
  nor _45934_ (_06203_, _05508_, rst);
  nor _45935_ (_23008_, _22886_, _22221_);
  and _45936_ (_23009_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _45937_ (_23010_, _23009_, _22886_);
  or _45938_ (_23011_, _23010_, _23008_);
  and _45939_ (_06204_, _23011_, _25365_);
  and _45940_ (_23012_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nor _45941_ (_23013_, _22886_, _22245_);
  or _45942_ (_23014_, _23013_, _23012_);
  and _45943_ (_06205_, _23014_, _25365_);
  nor _45944_ (_23015_, _22886_, _22261_);
  and _45945_ (_23016_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _45946_ (_23017_, _23016_, _23015_);
  and _45947_ (_06206_, _23017_, _25365_);
  nor _45948_ (_23018_, _22886_, _22282_);
  and _45949_ (_23019_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or _45950_ (_23020_, _23019_, _23018_);
  and _45951_ (_06207_, _23020_, _25365_);
  and _45952_ (_23021_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nor _45953_ (_23022_, _22886_, _22300_);
  or _45954_ (_23023_, _23022_, _23021_);
  and _45955_ (_06208_, _23023_, _25365_);
  and _45956_ (_23024_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nor _45957_ (_23025_, _22886_, _22315_);
  or _45958_ (_23026_, _23025_, _23024_);
  and _45959_ (_06209_, _23026_, _25365_);
  nor _45960_ (_23027_, _22886_, _22333_);
  and _45961_ (_23028_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _45962_ (_23029_, _23028_, _22886_);
  or _45963_ (_23030_, _23029_, _23027_);
  and _45964_ (_06210_, _23030_, _25365_);
  nor _45965_ (_23031_, _22886_, _22200_);
  and _45966_ (_23032_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _45967_ (_23033_, _23032_, _23031_);
  and _45968_ (_06211_, _23033_, _25365_);
  and _45969_ (_23034_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _45970_ (_23035_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _45971_ (_23036_, _23035_, _23034_);
  and _45972_ (_06212_, _23036_, _25365_);
  and _45973_ (_23037_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _45974_ (_23038_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _45975_ (_23039_, _23038_, _23037_);
  and _45976_ (_06213_, _23039_, _25365_);
  and _45977_ (_23040_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _45978_ (_23041_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _45979_ (_23042_, _23041_, _23040_);
  and _45980_ (_06214_, _23042_, _25365_);
  and _45981_ (_23043_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _45982_ (_23044_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _45983_ (_23045_, _23044_, _23043_);
  and _45984_ (_06215_, _23045_, _25365_);
  and _45985_ (_23046_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _45986_ (_23047_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _45987_ (_23048_, _23047_, _23046_);
  and _45988_ (_06216_, _23048_, _25365_);
  and _45989_ (_23049_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _45990_ (_23050_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _45991_ (_23051_, _23050_, _23049_);
  and _45992_ (_06217_, _23051_, _25365_);
  and _45993_ (_23052_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _45994_ (_23053_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _45995_ (_23054_, _23053_, _23052_);
  and _45996_ (_06218_, _23054_, _25365_);
  and _45997_ (_23055_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _45998_ (_23056_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _45999_ (_23057_, _23056_, _23055_);
  and _46000_ (_06219_, _23057_, _25365_);
  and _46001_ (_23058_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _46002_ (_23059_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _46003_ (_23060_, _23059_, _23058_);
  and _46004_ (_06220_, _23060_, _25365_);
  and _46005_ (_23061_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _46006_ (_23062_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _46007_ (_23063_, _23062_, _23061_);
  and _46008_ (_06221_, _23063_, _25365_);
  and _46009_ (_23064_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _46010_ (_23065_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _46011_ (_23066_, _23065_, _23064_);
  and _46012_ (_06222_, _23066_, _25365_);
  and _46013_ (_23067_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _46014_ (_23068_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _46015_ (_23069_, _23068_, _23067_);
  and _46016_ (_06223_, _23069_, _25365_);
  and _46017_ (_23070_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _46018_ (_23071_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _46019_ (_23072_, _23071_, _23070_);
  and _46020_ (_06224_, _23072_, _25365_);
  and _46021_ (_23073_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _46022_ (_23074_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _46023_ (_23075_, _23074_, _23073_);
  and _46024_ (_06225_, _23075_, _25365_);
  and _46025_ (_23076_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _46026_ (_23077_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _46027_ (_23078_, _23077_, _23076_);
  and _46028_ (_06226_, _23078_, _25365_);
  and _46029_ (_23079_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _46030_ (_23080_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _46031_ (_23081_, _23080_, _23079_);
  and _46032_ (_06227_, _23081_, _25365_);
  and _46033_ (_23082_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _46034_ (_23083_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _46035_ (_23084_, _23083_, _23082_);
  and _46036_ (_06228_, _23084_, _25365_);
  and _46037_ (_23085_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _46038_ (_23086_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _46039_ (_23087_, _23086_, _23085_);
  and _46040_ (_06229_, _23087_, _25365_);
  and _46041_ (_23088_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _46042_ (_23089_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _46043_ (_23090_, _23089_, _23088_);
  and _46044_ (_06230_, _23090_, _25365_);
  and _46045_ (_23091_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _46046_ (_23092_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _46047_ (_23093_, _23092_, _23091_);
  and _46048_ (_06231_, _23093_, _25365_);
  and _46049_ (_23094_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _46050_ (_23095_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _46051_ (_23096_, _23095_, _23094_);
  and _46052_ (_06232_, _23096_, _25365_);
  and _46053_ (_23097_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _46054_ (_23098_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _46055_ (_23099_, _23098_, _23097_);
  and _46056_ (_06233_, _23099_, _25365_);
  and _46057_ (_23100_, _22886_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _46058_ (_23101_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _46059_ (_23102_, _23101_, _23100_);
  and _46060_ (_06234_, _23102_, _25365_);
  nor _46061_ (_06235_, _05689_, rst);
  nor _46062_ (_06236_, _05987_, rst);
  nor _46063_ (_06237_, _05911_, rst);
  nor _46064_ (_06238_, _05642_, rst);
  nor _46065_ (_06239_, _05767_, rst);
  nor _46066_ (_06240_, _05797_, rst);
  nor _46067_ (_06241_, _05844_, rst);
  and _46068_ (_06256_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _25365_);
  and _46069_ (_06258_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _25365_);
  and _46070_ (_06259_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _25365_);
  and _46071_ (_06260_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _25365_);
  and _46072_ (_06261_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _25365_);
  and _46073_ (_06262_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _25365_);
  and _46074_ (_06263_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _25365_);
  or _46075_ (_23103_, _22591_, _22581_);
  and _46076_ (_23104_, _23103_, _01337_);
  and _46077_ (_23105_, _02083_, _02126_);
  and _46078_ (_23106_, _23105_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _46079_ (_23107_, _02125_, _02101_);
  and _46080_ (_23108_, _23107_, _01756_);
  and _46081_ (_23109_, _23108_, _22528_);
  nor _46082_ (_23110_, _22006_, _02080_);
  and _46083_ (_23111_, _23110_, _22395_);
  and _46084_ (_23112_, _23111_, _22425_);
  nor _46085_ (_23113_, _23112_, _05597_);
  not _46086_ (_23114_, _23113_);
  and _46087_ (_23115_, _01998_, _01756_);
  and _46088_ (_23116_, _23115_, _01852_);
  not _46089_ (_23117_, _23116_);
  and _46090_ (_23118_, _23117_, _22353_);
  and _46091_ (_23119_, _23118_, _23114_);
  nor _46092_ (_23120_, _23108_, _23105_);
  and _46093_ (_23121_, _23120_, _23117_);
  and _46094_ (_23122_, _23121_, _22484_);
  and _46095_ (_23123_, _23122_, _22353_);
  and _46096_ (_23124_, _22583_, _23123_);
  and _46097_ (_23125_, _23124_, _23119_);
  and _46098_ (_23126_, _23125_, _05670_);
  or _46099_ (_23127_, _23126_, _23109_);
  or _46100_ (_23128_, _23127_, _23106_);
  or _46101_ (_23129_, _23128_, _23104_);
  and _46102_ (_23130_, _22389_, _00907_);
  and _46103_ (_23131_, _23130_, _01186_);
  and _46104_ (_23132_, _22444_, _22411_);
  nor _46105_ (_23133_, _23132_, _22443_);
  not _46106_ (_23134_, _23133_);
  nor _46107_ (_23135_, _23134_, _23131_);
  and _46108_ (_23136_, _22450_, _22407_);
  nor _46109_ (_23137_, _23136_, _22375_);
  and _46110_ (_23138_, _23137_, _23135_);
  or _46111_ (_23139_, _22530_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _46112_ (_23140_, _22531_);
  nor _46113_ (_23141_, _23124_, _23119_);
  and _46114_ (_23142_, _23141_, _23140_);
  nand _46115_ (_23143_, _23142_, _23139_);
  nand _46116_ (_23144_, _23143_, _23138_);
  or _46117_ (_23145_, _23144_, _23129_);
  or _46118_ (_23146_, _23138_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _46119_ (_23147_, _23146_, _25365_);
  and _46120_ (_06264_, _23147_, _23145_);
  not _46121_ (_23148_, _23138_);
  and _46122_ (_23149_, _23103_, _01397_);
  or _46123_ (_23150_, _22533_, _22531_);
  and _46124_ (_23151_, _22585_, _22535_);
  and _46125_ (_23152_, _23151_, _23150_);
  and _46126_ (_23153_, _22485_, _22523_);
  and _46127_ (_23154_, _02084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _46128_ (_23155_, _22607_, _05967_);
  or _46129_ (_23156_, _23155_, _23154_);
  or _46130_ (_23157_, _23156_, _23153_);
  or _46131_ (_23158_, _23157_, _23152_);
  or _46132_ (_23159_, _23158_, _23149_);
  or _46133_ (_23160_, _23159_, _23148_);
  or _46134_ (_23161_, _23138_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _46135_ (_23162_, _23161_, _25365_);
  and _46136_ (_06265_, _23162_, _23160_);
  and _46137_ (_23163_, _22461_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _46138_ (_23164_, _22461_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _46139_ (_23165_, _23164_, _23163_);
  nor _46140_ (_23166_, _23165_, _22456_);
  and _46141_ (_23167_, _23103_, _01457_);
  or _46142_ (_23168_, _22538_, _22536_);
  and _46143_ (_23169_, _22585_, _22540_);
  and _46144_ (_23170_, _23169_, _23168_);
  and _46145_ (_23171_, _22485_, _22518_);
  and _46146_ (_23172_, _02084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _46147_ (_23173_, _22607_, _05892_);
  or _46148_ (_23174_, _23173_, _23172_);
  or _46149_ (_23175_, _23174_, _23171_);
  or _46150_ (_23176_, _23175_, _23170_);
  or _46151_ (_23177_, _23176_, _23167_);
  and _46152_ (_23178_, _23177_, _22456_);
  or _46153_ (_23179_, _23178_, _23166_);
  and _46154_ (_06266_, _23179_, _25365_);
  and _46155_ (_23180_, _23163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _46156_ (_23181_, _23163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _46157_ (_23182_, _23181_, _23180_);
  nor _46158_ (_23183_, _23182_, _22456_);
  and _46159_ (_23184_, _23103_, _01522_);
  or _46160_ (_23185_, _22515_, _22516_);
  not _46161_ (_23186_, _23185_);
  nand _46162_ (_23187_, _23186_, _22541_);
  or _46163_ (_23188_, _23186_, _22541_);
  and _46164_ (_23189_, _23188_, _22585_);
  and _46165_ (_23190_, _23189_, _23187_);
  not _46166_ (_23191_, _22290_);
  and _46167_ (_23192_, _22485_, _23191_);
  and _46168_ (_23193_, _02084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _46169_ (_23194_, _22607_, _05621_);
  or _46170_ (_23195_, _23194_, _23193_);
  or _46171_ (_23196_, _23195_, _23192_);
  or _46172_ (_23197_, _23196_, _23190_);
  or _46173_ (_23198_, _23197_, _23184_);
  and _46174_ (_23199_, _23198_, _22456_);
  or _46175_ (_23200_, _23199_, _23183_);
  and _46176_ (_06267_, _23200_, _25365_);
  and _46177_ (_23201_, _23103_, _01589_);
  or _46178_ (_23202_, _22545_, _22543_);
  and _46179_ (_23203_, _22585_, _22546_);
  and _46180_ (_23204_, _23203_, _23202_);
  not _46181_ (_23205_, _22308_);
  and _46182_ (_23206_, _22485_, _23205_);
  and _46183_ (_23207_, _22607_, _05746_);
  and _46184_ (_23208_, _02084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _46185_ (_23209_, _23208_, _23207_);
  or _46186_ (_23210_, _23209_, _23206_);
  nor _46187_ (_23211_, _23210_, _23204_);
  nand _46188_ (_23212_, _23211_, _22456_);
  or _46189_ (_23213_, _23212_, _23201_);
  and _46190_ (_23214_, _22463_, _22461_);
  nor _46191_ (_23215_, _23180_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _46192_ (_23216_, _23215_, _23214_);
  or _46193_ (_23217_, _23216_, _22456_);
  and _46194_ (_23218_, _23217_, _25365_);
  and _46195_ (_06268_, _23218_, _23213_);
  nor _46196_ (_23219_, _23214_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _46197_ (_23220_, _23219_, _22465_);
  nor _46198_ (_23221_, _23220_, _22456_);
  and _46199_ (_23222_, _23103_, _01673_);
  or _46200_ (_23223_, _22506_, _22507_);
  not _46201_ (_23224_, _23223_);
  nand _46202_ (_23225_, _23224_, _22547_);
  or _46203_ (_23226_, _23224_, _22547_);
  and _46204_ (_23227_, _23226_, _22585_);
  and _46205_ (_23228_, _23227_, _23225_);
  and _46206_ (_23229_, _22607_, _05814_);
  not _46207_ (_23230_, _22326_);
  and _46208_ (_23231_, _22485_, _23230_);
  and _46209_ (_23232_, _02084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _46210_ (_23233_, _23232_, _23231_);
  or _46211_ (_23234_, _23233_, _23229_);
  or _46212_ (_23235_, _23234_, _23228_);
  or _46213_ (_23236_, _23235_, _23222_);
  and _46214_ (_23237_, _23236_, _22456_);
  or _46215_ (_23238_, _23237_, _23221_);
  and _46216_ (_06269_, _23238_, _25365_);
  nor _46217_ (_23239_, _22465_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _46218_ (_23240_, _23239_, _22466_);
  nor _46219_ (_23241_, _23240_, _22456_);
  and _46220_ (_23242_, _23103_, _01737_);
  and _46221_ (_23243_, _23105_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _46222_ (_23244_, _22344_);
  and _46223_ (_23245_, _23108_, _23244_);
  and _46224_ (_23246_, _23125_, _05864_);
  or _46225_ (_23247_, _23246_, _23245_);
  or _46226_ (_23248_, _23247_, _23243_);
  or _46227_ (_23249_, _22549_, _22502_);
  and _46228_ (_23250_, _23249_, _22550_);
  and _46229_ (_23251_, _23250_, _23141_);
  or _46230_ (_23252_, _23251_, _23248_);
  or _46231_ (_23253_, _23252_, _23242_);
  and _46232_ (_23254_, _23253_, _22456_);
  or _46233_ (_23255_, _23254_, _23241_);
  and _46234_ (_06270_, _23255_, _25365_);
  nor _46235_ (_23256_, _22466_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _46236_ (_23257_, _23256_, _22467_);
  or _46237_ (_23258_, _23257_, _22456_);
  and _46238_ (_23259_, _23258_, _25365_);
  and _46239_ (_23260_, _23105_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _46240_ (_23261_, _23103_, _01184_);
  not _46241_ (_23262_, _22212_);
  and _46242_ (_23263_, _23108_, _23262_);
  and _46243_ (_23264_, _23125_, _05580_);
  or _46244_ (_23265_, _23264_, _23263_);
  or _46245_ (_23266_, _22493_, _22494_);
  not _46246_ (_23267_, _23266_);
  nand _46247_ (_23268_, _23267_, _22551_);
  or _46248_ (_23269_, _23267_, _22551_);
  and _46249_ (_23270_, _23269_, _23141_);
  and _46250_ (_23271_, _23270_, _23268_);
  or _46251_ (_23272_, _23271_, _23265_);
  or _46252_ (_23273_, _23272_, _23261_);
  nor _46253_ (_23274_, _23273_, _23260_);
  nand _46254_ (_23275_, _23274_, _23138_);
  and _46255_ (_06271_, _23275_, _23259_);
  nor _46256_ (_23276_, _22467_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _46257_ (_23277_, _23276_, _22468_);
  or _46258_ (_23278_, _23277_, _22456_);
  and _46259_ (_23279_, _23278_, _25365_);
  and _46260_ (_23280_, _22553_, _02374_);
  nor _46261_ (_23281_, _22553_, _02374_);
  nor _46262_ (_23282_, _23281_, _23280_);
  nor _46263_ (_23283_, _23282_, _22492_);
  and _46264_ (_23284_, _23282_, _22492_);
  or _46265_ (_23285_, _23284_, _23283_);
  and _46266_ (_23286_, _23285_, _23141_);
  and _46267_ (_23287_, _23105_, _01337_);
  and _46268_ (_23288_, _23125_, _21716_);
  and _46269_ (_23289_, _22581_, _02451_);
  and _46270_ (_23290_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _46271_ (_23291_, _23108_, _05670_);
  or _46272_ (_23292_, _23291_, _23290_);
  or _46273_ (_23293_, _23292_, _23289_);
  or _46274_ (_23294_, _23293_, _23288_);
  or _46275_ (_23295_, _23294_, _23287_);
  or _46276_ (_23296_, _23295_, _23286_);
  or _46277_ (_23297_, _23296_, _23148_);
  and _46278_ (_06272_, _23297_, _23279_);
  nor _46279_ (_23298_, _22468_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _46280_ (_23299_, _23298_, _22469_);
  or _46281_ (_23300_, _23299_, _22456_);
  and _46282_ (_23301_, _23300_, _25365_);
  and _46283_ (_23302_, _22553_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _46284_ (_23303_, _23302_, _22561_);
  nor _46285_ (_23304_, _22562_, _22561_);
  nor _46286_ (_23305_, _23304_, _23303_);
  nand _46287_ (_23306_, _23305_, _02380_);
  or _46288_ (_23307_, _23305_, _02380_);
  and _46289_ (_23308_, _23307_, _22585_);
  and _46290_ (_23309_, _23308_, _23306_);
  and _46291_ (_23310_, _02084_, _01397_);
  not _46292_ (_23311_, _22581_);
  nor _46293_ (_23312_, _23311_, _02481_);
  and _46294_ (_23313_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _46295_ (_23314_, _22485_, _05967_);
  and _46296_ (_23315_, _22607_, _21694_);
  or _46297_ (_23316_, _23315_, _23314_);
  or _46298_ (_23317_, _23316_, _23313_);
  nor _46299_ (_23318_, _23317_, _23312_);
  nand _46300_ (_23319_, _23318_, _22456_);
  or _46301_ (_23320_, _23319_, _23310_);
  or _46302_ (_23321_, _23320_, _23309_);
  and _46303_ (_06273_, _23321_, _23301_);
  nor _46304_ (_23322_, _22469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _46305_ (_23323_, _23322_, _22470_);
  or _46306_ (_23324_, _23323_, _22456_);
  and _46307_ (_23325_, _23324_, _25365_);
  and _46308_ (_23326_, _23304_, _02380_);
  and _46309_ (_23327_, _23303_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _46310_ (_23328_, _23327_, _23326_);
  nand _46311_ (_23329_, _23328_, _02385_);
  or _46312_ (_23330_, _23328_, _02385_);
  and _46313_ (_23331_, _23330_, _22585_);
  and _46314_ (_23332_, _23331_, _23329_);
  and _46315_ (_23333_, _02084_, _01457_);
  nor _46316_ (_23334_, _23311_, _02511_);
  and _46317_ (_23335_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _46318_ (_23336_, _22485_, _05892_);
  and _46319_ (_23337_, _22607_, _21654_);
  or _46320_ (_23338_, _23337_, _23336_);
  or _46321_ (_23339_, _23338_, _23335_);
  nor _46322_ (_23340_, _23339_, _23334_);
  nand _46323_ (_23341_, _23340_, _22456_);
  or _46324_ (_23342_, _23341_, _23333_);
  or _46325_ (_23343_, _23342_, _23332_);
  and _46326_ (_06274_, _23343_, _23325_);
  nor _46327_ (_23344_, _22470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _46328_ (_23345_, _22470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _46329_ (_23346_, _23345_, _23344_);
  or _46330_ (_23347_, _23346_, _22456_);
  and _46331_ (_23348_, _23347_, _25365_);
  and _46332_ (_23349_, _22556_, _22561_);
  nor _46333_ (_23350_, _22564_, _22561_);
  or _46334_ (_23351_, _23350_, _23349_);
  nand _46335_ (_23352_, _23351_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _46336_ (_23353_, _23351_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _46337_ (_23354_, _23353_, _22585_);
  and _46338_ (_23355_, _23354_, _23352_);
  and _46339_ (_23356_, _02084_, _01522_);
  nor _46340_ (_23357_, _23311_, _02540_);
  and _46341_ (_23358_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _46342_ (_23359_, _22599_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _46343_ (_23360_, _23359_, _22600_);
  and _46344_ (_23361_, _23360_, _22607_);
  and _46345_ (_23362_, _22485_, _05621_);
  or _46346_ (_23363_, _23362_, _23361_);
  or _46347_ (_23364_, _23363_, _23358_);
  nor _46348_ (_23365_, _23364_, _23357_);
  nand _46349_ (_23366_, _23365_, _22456_);
  or _46350_ (_23367_, _23366_, _23356_);
  or _46351_ (_23368_, _23367_, _23355_);
  and _46352_ (_06275_, _23368_, _23348_);
  nor _46353_ (_23369_, _23345_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _46354_ (_23370_, _23369_, _22472_);
  or _46355_ (_23371_, _23370_, _22456_);
  and _46356_ (_23372_, _23371_, _25365_);
  and _46357_ (_23373_, _22557_, _22561_);
  nor _46358_ (_23374_, _22565_, _22561_);
  nor _46359_ (_23375_, _23374_, _23373_);
  nand _46360_ (_23376_, _23375_, _02391_);
  or _46361_ (_23377_, _23375_, _02391_);
  and _46362_ (_23378_, _23377_, _23376_);
  and _46363_ (_23379_, _23378_, _23141_);
  nor _46364_ (_23380_, _22600_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _46365_ (_23381_, _23380_, _22601_);
  and _46366_ (_23382_, _23381_, _23125_);
  and _46367_ (_23383_, _23105_, _01589_);
  nor _46368_ (_23384_, _23311_, _02572_);
  and _46369_ (_23385_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _46370_ (_23386_, _23108_, _05746_);
  or _46371_ (_23387_, _23386_, _23385_);
  or _46372_ (_23388_, _23387_, _23384_);
  or _46373_ (_23389_, _23388_, _23383_);
  nor _46374_ (_23390_, _23389_, _23382_);
  nand _46375_ (_23391_, _23390_, _23138_);
  or _46376_ (_23392_, _23391_, _23379_);
  and _46377_ (_06276_, _23392_, _23372_);
  and _46378_ (_23393_, _02084_, _01673_);
  nor _46379_ (_23394_, _23311_, _02604_);
  and _46380_ (_23395_, _22485_, _05814_);
  and _46381_ (_23396_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _46382_ (_23397_, _22601_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _46383_ (_23398_, _23397_, _22602_);
  and _46384_ (_23399_, _23398_, _22607_);
  or _46385_ (_23400_, _23399_, _23396_);
  or _46386_ (_23401_, _23400_, _23395_);
  or _46387_ (_23402_, _23401_, _23394_);
  or _46388_ (_23403_, _23402_, _23393_);
  nand _46389_ (_23404_, _23373_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _46390_ (_23405_, _22566_, _22561_);
  and _46391_ (_23406_, _23405_, _23404_);
  nor _46392_ (_23407_, _23406_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _46393_ (_23408_, _23406_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _46394_ (_23409_, _23408_, _23407_);
  and _46395_ (_23410_, _23409_, _22585_);
  or _46396_ (_23411_, _23410_, _23403_);
  or _46397_ (_23412_, _23411_, _23148_);
  nor _46398_ (_23413_, _22472_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _46399_ (_23414_, _23413_, _22473_);
  or _46400_ (_23415_, _23414_, _23138_);
  and _46401_ (_23416_, _23415_, _25365_);
  and _46402_ (_06277_, _23416_, _23412_);
  and _46403_ (_23417_, _02084_, _01737_);
  nor _46404_ (_23418_, _23311_, _02634_);
  and _46405_ (_23419_, _22591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _46406_ (_23420_, _22485_, _05864_);
  or _46407_ (_23421_, _23420_, _23419_);
  or _46408_ (_23422_, _22602_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _46409_ (_23423_, _23422_, _22603_);
  and _46410_ (_23424_, _23423_, _22607_);
  or _46411_ (_23425_, _23424_, _23421_);
  or _46412_ (_23426_, _23425_, _23418_);
  or _46413_ (_23427_, _23426_, _23417_);
  nor _46414_ (_23428_, _22569_, _02397_);
  and _46415_ (_23429_, _22569_, _02397_);
  or _46416_ (_23430_, _23429_, _23428_);
  and _46417_ (_23431_, _23430_, _22585_);
  or _46418_ (_23432_, _23431_, _23427_);
  or _46419_ (_23433_, _23432_, _23148_);
  nor _46420_ (_23434_, _22473_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _46421_ (_23435_, _23434_, _22474_);
  or _46422_ (_23436_, _23435_, _23138_);
  and _46423_ (_23437_, _23436_, _25365_);
  and _46424_ (_06278_, _23437_, _23433_);
  and _46425_ (_23438_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _46426_ (_23439_, _22783_, _22781_);
  nor _46427_ (_23440_, _23439_, _22784_);
  or _46428_ (_23441_, _23440_, _22618_);
  or _46429_ (_23442_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _46430_ (_23443_, _23442_, _22820_);
  and _46431_ (_23444_, _23443_, _23441_);
  or _46432_ (_06279_, _23444_, _23438_);
  and _46433_ (_23445_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _46434_ (_23446_, _22786_, _22784_);
  and _46435_ (_23447_, _23446_, _22787_);
  or _46436_ (_23448_, _23447_, _22618_);
  or _46437_ (_23449_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _46438_ (_23450_, _23449_, _22820_);
  and _46439_ (_23451_, _23450_, _23448_);
  or _46440_ (_06280_, _23451_, _23445_);
  or _46441_ (_23452_, _22791_, _22789_);
  nor _46442_ (_23453_, _22792_, _22618_);
  and _46443_ (_23454_, _23453_, _23452_);
  nor _46444_ (_23455_, _22617_, _00317_);
  or _46445_ (_23456_, _23455_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _46446_ (_23457_, _23456_, _23454_);
  or _46447_ (_23458_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _01757_);
  and _46448_ (_23459_, _23458_, _25365_);
  and _46449_ (_06281_, _23459_, _23457_);
  and _46450_ (_23460_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _46451_ (_23461_, _22792_, _22686_);
  nor _46452_ (_23462_, _23461_, _22793_);
  or _46453_ (_23463_, _23462_, _22618_);
  or _46454_ (_23464_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _46455_ (_23465_, _23464_, _22820_);
  and _46456_ (_23466_, _23465_, _23463_);
  or _46457_ (_06282_, _23466_, _23460_);
  and _46458_ (_23467_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _46459_ (_23468_, _22796_, _22793_);
  nor _46460_ (_23469_, _23468_, _22797_);
  or _46461_ (_23470_, _23469_, _22618_);
  or _46462_ (_23471_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _46463_ (_23472_, _23471_, _22820_);
  and _46464_ (_23473_, _23472_, _23470_);
  or _46465_ (_06283_, _23473_, _23467_);
  and _46466_ (_23474_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _46467_ (_23475_, _22797_, _22681_);
  nor _46468_ (_23476_, _23475_, _22798_);
  or _46469_ (_23477_, _23476_, _22618_);
  or _46470_ (_23478_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _46471_ (_23479_, _23478_, _22820_);
  and _46472_ (_23480_, _23479_, _23477_);
  or _46473_ (_06284_, _23480_, _23474_);
  nor _46474_ (_23481_, _22798_, _22677_);
  nor _46475_ (_23482_, _23481_, _22799_);
  or _46476_ (_23483_, _23482_, _22618_);
  or _46477_ (_23484_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _46478_ (_23485_, _23484_, _22820_);
  and _46479_ (_23486_, _23485_, _23483_);
  and _46480_ (_23487_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _46481_ (_06285_, _23487_, _23486_);
  nor _46482_ (_23488_, _22799_, _22673_);
  nor _46483_ (_23489_, _23488_, _22800_);
  or _46484_ (_23490_, _23489_, _22618_);
  or _46485_ (_23491_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _46486_ (_23492_, _23491_, _22820_);
  and _46487_ (_23493_, _23492_, _23490_);
  and _46488_ (_23494_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _46489_ (_06286_, _23494_, _23493_);
  and _46490_ (_23495_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _46491_ (_23496_, _22802_, _22800_);
  nor _46492_ (_23497_, _23496_, _22803_);
  or _46493_ (_23498_, _23497_, _22618_);
  or _46494_ (_23499_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _46495_ (_23500_, _23499_, _22820_);
  and _46496_ (_23501_, _23500_, _23498_);
  or _46497_ (_06287_, _23501_, _23495_);
  nor _46498_ (_23502_, _22803_, _22669_);
  nor _46499_ (_23503_, _23502_, _22804_);
  or _46500_ (_23504_, _23503_, _22618_);
  or _46501_ (_23505_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _46502_ (_23506_, _23505_, _22820_);
  and _46503_ (_23507_, _23506_, _23504_);
  and _46504_ (_23508_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _46505_ (_06288_, _23508_, _23507_);
  and _46506_ (_23509_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _46507_ (_23510_, _22804_, _22666_);
  nor _46508_ (_23511_, _23510_, _22805_);
  or _46509_ (_23512_, _23511_, _22618_);
  or _46510_ (_23513_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _46511_ (_23514_, _23513_, _22820_);
  and _46512_ (_23515_, _23514_, _23512_);
  or _46513_ (_06289_, _23515_, _23509_);
  nor _46514_ (_23516_, _22805_, _22664_);
  nor _46515_ (_23517_, _23516_, _22806_);
  or _46516_ (_23518_, _23517_, _22618_);
  or _46517_ (_23519_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _46518_ (_23520_, _23519_, _22820_);
  and _46519_ (_23521_, _23520_, _23518_);
  and _46520_ (_23522_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _46521_ (_06290_, _23522_, _23521_);
  nor _46522_ (_23523_, _22806_, _22661_);
  nor _46523_ (_23524_, _23523_, _22807_);
  or _46524_ (_23525_, _23524_, _22618_);
  or _46525_ (_23526_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _46526_ (_23527_, _23526_, _22820_);
  and _46527_ (_23528_, _23527_, _23525_);
  and _46528_ (_23529_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _46529_ (_06291_, _23529_, _23528_);
  nor _46530_ (_23530_, _22807_, _22658_);
  nor _46531_ (_23531_, _23530_, _22808_);
  or _46532_ (_23532_, _23531_, _22618_);
  or _46533_ (_23533_, _22617_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _46534_ (_23534_, _23533_, _22820_);
  and _46535_ (_23535_, _23534_, _23532_);
  and _46536_ (_23536_, _22823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _46537_ (_06292_, _23536_, _23535_);
  or _46538_ (_23537_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _01757_);
  and _46539_ (_23538_, _23537_, _25365_);
  or _46540_ (_23539_, _22808_, _22655_);
  and _46541_ (_23540_, _23539_, _22810_);
  nor _46542_ (_23541_, _22617_, _02397_);
  or _46543_ (_23542_, _23541_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _46544_ (_23543_, _23542_, _23540_);
  and _46545_ (_06293_, _23543_, _23538_);
  and _46546_ (_23544_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _46547_ (_23545_, _23544_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _46548_ (_06294_, _23545_, _25365_);
  and _46549_ (_23546_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _46550_ (_23547_, _23546_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _46551_ (_06295_, _23547_, _25365_);
  and _46552_ (_23548_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _46553_ (_23549_, _23548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _46554_ (_06296_, _23549_, _25365_);
  and _46555_ (_23550_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _46556_ (_23551_, _23550_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _46557_ (_06297_, _23551_, _25365_);
  and _46558_ (_23552_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _46559_ (_23553_, _23552_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _46560_ (_06298_, _23553_, _25365_);
  and _46561_ (_23554_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _46562_ (_23555_, _23554_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _46563_ (_06299_, _23555_, _25365_);
  and _46564_ (_23556_, _22832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _46565_ (_23557_, _23556_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _46566_ (_06300_, _23557_, _25365_);
  nor _46567_ (_23558_, _22780_, _05562_);
  and _46568_ (_23559_, _23558_, _01787_);
  nor _46569_ (_23560_, _23558_, _01787_);
  or _46570_ (_23561_, _23560_, _23559_);
  and _46571_ (_06301_, _23561_, _22820_);
  or _46572_ (_23562_, _22843_, _22841_);
  and _46573_ (_23563_, _23562_, _22844_);
  or _46574_ (_23564_, _23563_, _05562_);
  or _46575_ (_23565_, _01760_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _46576_ (_23566_, _23565_, _22820_);
  and _46577_ (_06302_, _23566_, _23564_);
  and _46578_ (_23567_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _46579_ (_23568_, _23009_, _06132_);
  or _46580_ (_06317_, _23568_, _23567_);
  and _46581_ (_23569_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _46582_ (_23570_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _46583_ (_23571_, _23570_, _06132_);
  or _46584_ (_06318_, _23571_, _23569_);
  and _46585_ (_23572_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _46586_ (_23573_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _46587_ (_23574_, _23573_, _06132_);
  or _46588_ (_06319_, _23574_, _23572_);
  and _46589_ (_23575_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _46590_ (_23576_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _46591_ (_23577_, _23576_, _06132_);
  or _46592_ (_06320_, _23577_, _23575_);
  and _46593_ (_23578_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _46594_ (_23579_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _46595_ (_23580_, _23579_, _06132_);
  or _46596_ (_06321_, _23580_, _23578_);
  and _46597_ (_23581_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _46598_ (_23582_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _46599_ (_23583_, _23582_, _06132_);
  or _46600_ (_06322_, _23583_, _23581_);
  and _46601_ (_23584_, _22864_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _46602_ (_23585_, _23028_, _06132_);
  or _46603_ (_06323_, _23585_, _23584_);
  and _46604_ (_06324_, _22872_, _25365_);
  nor _46605_ (_06325_, _22882_, rst);
  and _46606_ (_06326_, _22878_, _25365_);
  or _46607_ (_23586_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand _46608_ (_23587_, _22886_, _22221_);
  and _46609_ (_23588_, _23587_, _25365_);
  and _46610_ (_06327_, _23588_, _23586_);
  or _46611_ (_23589_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nand _46612_ (_23590_, _22886_, _22245_);
  and _46613_ (_23591_, _23590_, _25365_);
  and _46614_ (_06328_, _23591_, _23589_);
  or _46615_ (_23592_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand _46616_ (_23593_, _22886_, _22261_);
  and _46617_ (_23594_, _23593_, _25365_);
  and _46618_ (_06329_, _23594_, _23592_);
  or _46619_ (_23595_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _46620_ (_23596_, _22886_, _22282_);
  and _46621_ (_23597_, _23596_, _25365_);
  and _46622_ (_06330_, _23597_, _23595_);
  or _46623_ (_23598_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand _46624_ (_23599_, _22886_, _22300_);
  and _46625_ (_23600_, _23599_, _25365_);
  and _46626_ (_06331_, _23600_, _23598_);
  or _46627_ (_23601_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _46628_ (_23602_, _22886_, _22315_);
  and _46629_ (_23603_, _23602_, _25365_);
  and _46630_ (_06332_, _23603_, _23601_);
  or _46631_ (_23604_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _46632_ (_23605_, _22886_, _22333_);
  and _46633_ (_23606_, _23605_, _25365_);
  and _46634_ (_06333_, _23606_, _23604_);
  or _46635_ (_23607_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _46636_ (_23608_, _22886_, _22200_);
  and _46637_ (_23609_, _23608_, _25365_);
  and _46638_ (_06334_, _23609_, _23607_);
  and _46639_ (_23610_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _46640_ (_23611_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _46641_ (_23612_, _23611_, _23610_);
  and _46642_ (_06335_, _23612_, _25365_);
  and _46643_ (_23613_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _46644_ (_23614_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _46645_ (_23615_, _23614_, _23613_);
  and _46646_ (_06336_, _23615_, _25365_);
  and _46647_ (_23616_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _46648_ (_23617_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _46649_ (_23618_, _23617_, _23616_);
  and _46650_ (_06337_, _23618_, _25365_);
  and _46651_ (_23619_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _46652_ (_23620_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _46653_ (_23621_, _23620_, _23619_);
  and _46654_ (_06338_, _23621_, _25365_);
  and _46655_ (_23622_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _46656_ (_23623_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _46657_ (_23624_, _23623_, _23622_);
  and _46658_ (_06339_, _23624_, _25365_);
  and _46659_ (_23625_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _46660_ (_23626_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _46661_ (_23627_, _23626_, _23625_);
  and _46662_ (_06340_, _23627_, _25365_);
  and _46663_ (_23628_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _46664_ (_23629_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _46665_ (_23630_, _23629_, _23628_);
  and _46666_ (_06341_, _23630_, _25365_);
  and _46667_ (_23631_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _46668_ (_23632_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _46669_ (_23633_, _23632_, _23631_);
  and _46670_ (_06342_, _23633_, _25365_);
  and _46671_ (_23634_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _46672_ (_23635_, _22886_, _01863_);
  or _46673_ (_23636_, _23635_, _23634_);
  and _46674_ (_06343_, _23636_, _25365_);
  and _46675_ (_23637_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor _46676_ (_23638_, _22886_, _01887_);
  or _46677_ (_23639_, _23638_, _23637_);
  and _46678_ (_06344_, _23639_, _25365_);
  and _46679_ (_23640_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _46680_ (_23641_, _22886_, _01908_);
  or _46681_ (_23642_, _23641_, _23640_);
  and _46682_ (_06345_, _23642_, _25365_);
  and _46683_ (_23643_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _46684_ (_23644_, _22886_, _01934_);
  or _46685_ (_23645_, _23644_, _23643_);
  and _46686_ (_06346_, _23645_, _25365_);
  and _46687_ (_23646_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _46688_ (_23647_, _22886_, _01961_);
  or _46689_ (_23648_, _23647_, _23646_);
  and _46690_ (_06347_, _23648_, _25365_);
  and _46691_ (_23649_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _46692_ (_23650_, _22886_, _01786_);
  or _46693_ (_23651_, _23650_, _23649_);
  and _46694_ (_06348_, _23651_, _25365_);
  and _46695_ (_23652_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _46696_ (_23653_, _22886_, _01835_);
  or _46697_ (_23654_, _23653_, _23652_);
  and _46698_ (_06349_, _23654_, _25365_);
  and _46699_ (_23655_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _46700_ (_23656_, _22886_, _01811_);
  or _46701_ (_23657_, _23656_, _23655_);
  and _46702_ (_06350_, _23657_, _25365_);
  and _46703_ (_23658_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor _46704_ (_23659_, _22886_, _05660_);
  or _46705_ (_23660_, _23659_, _23658_);
  and _46706_ (_06351_, _23660_, _25365_);
  and _46707_ (_23661_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor _46708_ (_23662_, _22886_, _05946_);
  or _46709_ (_23663_, _23662_, _23661_);
  and _46710_ (_06352_, _23663_, _25365_);
  and _46711_ (_23664_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _46712_ (_23665_, _22888_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _46713_ (_23666_, _23665_, _23664_);
  and _46714_ (_06353_, _23666_, _25365_);
  and _46715_ (_23667_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor _46716_ (_23668_, _22886_, _05611_);
  or _46717_ (_23669_, _23668_, _23667_);
  and _46718_ (_06354_, _23669_, _25365_);
  and _46719_ (_23670_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _46720_ (_23671_, _22886_, _05733_);
  or _46721_ (_23672_, _23671_, _23670_);
  and _46722_ (_06355_, _23672_, _25365_);
  and _46723_ (_23673_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _46724_ (_23674_, _22886_, _05801_);
  or _46725_ (_23675_, _23674_, _23673_);
  and _46726_ (_06356_, _23675_, _25365_);
  and _46727_ (_23676_, _22886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor _46728_ (_23677_, _22886_, _05851_);
  or _46729_ (_23678_, _23677_, _23676_);
  and _46730_ (_06357_, _23678_, _25365_);
  and _46731_ (_23679_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _46732_ (_23680_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _46733_ (_23681_, _23680_, _23679_);
  and _46734_ (_06359_, _23681_, _25365_);
  and _46735_ (_23682_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _46736_ (_23683_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _46737_ (_23684_, _23683_, _23682_);
  and _46738_ (_06360_, _23684_, _25365_);
  and _46739_ (_23685_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _46740_ (_23686_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _46741_ (_23687_, _23686_, _23685_);
  and _46742_ (_06361_, _23687_, _25365_);
  and _46743_ (_23688_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _46744_ (_23689_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _46745_ (_23690_, _23689_, _23688_);
  and _46746_ (_06362_, _23690_, _25365_);
  and _46747_ (_23691_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _46748_ (_23692_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _46749_ (_23693_, _23692_, _23691_);
  and _46750_ (_06363_, _23693_, _25365_);
  and _46751_ (_23694_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _46752_ (_23695_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _46753_ (_23696_, _23695_, _23694_);
  and _46754_ (_06364_, _23696_, _25365_);
  and _46755_ (_23697_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _46756_ (_23698_, _22896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _46757_ (_23699_, _23698_, _23697_);
  and _46758_ (_06365_, _23699_, _25365_);
  and _46759_ (_23700_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _46760_ (_23701_, _05689_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _46761_ (_23702_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _46762_ (_23703_, _23702_, _22895_);
  and _46763_ (_23704_, _23703_, _23701_);
  or _46764_ (_23705_, _23704_, _23700_);
  and _46765_ (_06366_, _23705_, _25365_);
  and _46766_ (_23706_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _46767_ (_23707_, _05987_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _46768_ (_23708_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _46769_ (_23709_, _23708_, _22895_);
  and _46770_ (_23710_, _23709_, _23707_);
  or _46771_ (_23711_, _23710_, _23706_);
  and _46772_ (_06367_, _23711_, _25365_);
  and _46773_ (_23712_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _46774_ (_23713_, _05911_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _46775_ (_23714_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _46776_ (_23715_, _23714_, _22895_);
  and _46777_ (_23716_, _23715_, _23713_);
  or _46778_ (_23717_, _23716_, _23712_);
  and _46779_ (_06368_, _23717_, _25365_);
  and _46780_ (_23718_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _46781_ (_23719_, _05642_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _46782_ (_23720_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _46783_ (_23721_, _23720_, _22895_);
  and _46784_ (_23722_, _23721_, _23719_);
  or _46785_ (_23723_, _23722_, _23718_);
  and _46786_ (_06369_, _23723_, _25365_);
  and _46787_ (_23724_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _46788_ (_23725_, _05767_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _46789_ (_23726_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _46790_ (_23727_, _23726_, _22895_);
  and _46791_ (_23728_, _23727_, _23725_);
  or _46792_ (_23729_, _23728_, _23724_);
  and _46793_ (_06370_, _23729_, _25365_);
  and _46794_ (_23730_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _46795_ (_23731_, _05797_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _46796_ (_23732_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _46797_ (_23733_, _23732_, _22895_);
  and _46798_ (_23734_, _23733_, _23731_);
  or _46799_ (_23735_, _23734_, _23730_);
  and _46800_ (_06371_, _23735_, _25365_);
  and _46801_ (_23736_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _46802_ (_23737_, _05844_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _46803_ (_23738_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _46804_ (_23739_, _23738_, _22895_);
  and _46805_ (_23740_, _23739_, _23737_);
  or _46806_ (_23741_, _23740_, _23736_);
  and _46807_ (_06372_, _23741_, _25365_);
  and _46808_ (_23742_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46809_ (_23743_, _05559_, _22902_);
  or _46810_ (_23744_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _46811_ (_23745_, _23744_, _22895_);
  and _46812_ (_23746_, _23745_, _23743_);
  or _46813_ (_23747_, _23746_, _23742_);
  and _46814_ (_06373_, _23747_, _25365_);
  and _46815_ (_23748_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _46816_ (_23749_, _23748_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46817_ (_23750_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _22895_);
  and _46818_ (_23751_, _23750_, _25365_);
  and _46819_ (_06374_, _23751_, _23749_);
  and _46820_ (_23752_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _46821_ (_23753_, _23752_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46822_ (_23754_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _22895_);
  and _46823_ (_23755_, _23754_, _25365_);
  and _46824_ (_06375_, _23755_, _23753_);
  and _46825_ (_23756_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _46826_ (_23757_, _23756_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46827_ (_23758_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _22895_);
  and _46828_ (_23759_, _23758_, _25365_);
  and _46829_ (_06376_, _23759_, _23757_);
  and _46830_ (_23760_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _46831_ (_23761_, _23760_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46832_ (_23762_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _22895_);
  and _46833_ (_23763_, _23762_, _25365_);
  and _46834_ (_06377_, _23763_, _23761_);
  and _46835_ (_23764_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _46836_ (_23765_, _23764_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46837_ (_23766_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _22895_);
  and _46838_ (_23767_, _23766_, _25365_);
  and _46839_ (_06378_, _23767_, _23765_);
  and _46840_ (_23768_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _46841_ (_23769_, _23768_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46842_ (_23770_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _22895_);
  and _46843_ (_23771_, _23770_, _25365_);
  and _46844_ (_06379_, _23771_, _23769_);
  and _46845_ (_23772_, _22902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _46846_ (_23773_, _23772_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _46847_ (_23774_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _22895_);
  and _46848_ (_23775_, _23774_, _25365_);
  and _46849_ (_06380_, _23775_, _23773_);
  or _46850_ (_23776_, _22914_, _01337_);
  or _46851_ (_23777_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _46852_ (_23778_, _23777_, _25365_);
  and _46853_ (_06381_, _23778_, _23776_);
  or _46854_ (_23779_, _22914_, _01397_);
  or _46855_ (_23780_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _46856_ (_23781_, _23780_, _25365_);
  and _46857_ (_06382_, _23781_, _23779_);
  or _46858_ (_23782_, _22914_, _01457_);
  or _46859_ (_23783_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _46860_ (_23784_, _23783_, _25365_);
  and _46861_ (_06383_, _23784_, _23782_);
  or _46862_ (_23785_, _22914_, _01522_);
  or _46863_ (_23786_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _46864_ (_23787_, _23786_, _25365_);
  and _46865_ (_06384_, _23787_, _23785_);
  or _46866_ (_23788_, _22914_, _01589_);
  or _46867_ (_23789_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _46868_ (_23790_, _23789_, _25365_);
  and _46869_ (_06385_, _23790_, _23788_);
  or _46870_ (_23791_, _22914_, _01673_);
  or _46871_ (_23792_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _46872_ (_23793_, _23792_, _25365_);
  and _46873_ (_06386_, _23793_, _23791_);
  or _46874_ (_23794_, _22914_, _01737_);
  or _46875_ (_23795_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _46876_ (_23796_, _23795_, _25365_);
  and _46877_ (_06387_, _23796_, _23794_);
  or _46878_ (_23797_, _22914_, _01184_);
  or _46879_ (_23798_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _46880_ (_23799_, _23798_, _25365_);
  and _46881_ (_06388_, _23799_, _23797_);
  or _46882_ (_23800_, _22914_, _02451_);
  or _46883_ (_23801_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _46884_ (_23802_, _23801_, _25365_);
  and _46885_ (_06389_, _23802_, _23800_);
  nand _46886_ (_23803_, _22909_, _02481_);
  or _46887_ (_23804_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _46888_ (_23805_, _23804_, _25365_);
  and _46889_ (_06390_, _23805_, _23803_);
  nand _46890_ (_23806_, _22909_, _02511_);
  or _46891_ (_23807_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _46892_ (_23808_, _23807_, _25365_);
  and _46893_ (_06391_, _23808_, _23806_);
  nand _46894_ (_23809_, _22909_, _02540_);
  or _46895_ (_23810_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _46896_ (_23811_, _23810_, _25365_);
  and _46897_ (_06392_, _23811_, _23809_);
  nand _46898_ (_23812_, _22909_, _02572_);
  or _46899_ (_23813_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _46900_ (_23814_, _23813_, _25365_);
  and _46901_ (_06393_, _23814_, _23812_);
  nand _46902_ (_23815_, _22909_, _02604_);
  or _46903_ (_23816_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _46904_ (_23817_, _23816_, _25365_);
  and _46905_ (_06394_, _23817_, _23815_);
  nand _46906_ (_23818_, _22909_, _02634_);
  or _46907_ (_23819_, _22909_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _46908_ (_23820_, _23819_, _25365_);
  and _46909_ (_06395_, _23820_, _23818_);
  nor _46910_ (_06419_, _05601_, rst);
  and _46911_ (_23821_, _05516_, _02159_);
  and _46912_ (_23822_, _23821_, _02783_);
  and _46913_ (_23823_, _23822_, _05518_);
  nand _46914_ (_23824_, _23823_, _02280_);
  or _46915_ (_23825_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _46916_ (_23826_, _23825_, _25365_);
  and _46917_ (_06420_, _23826_, _23824_);
  and _46918_ (_23827_, _23821_, _02982_);
  not _46919_ (_23828_, _23827_);
  nor _46920_ (_23829_, _23828_, _02280_);
  not _46921_ (_23830_, _05518_);
  and _46922_ (_23831_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _46923_ (_23832_, _23831_, _23830_);
  or _46924_ (_23833_, _23832_, _23829_);
  or _46925_ (_23834_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _46926_ (_23835_, _23834_, _25365_);
  and _46927_ (_06421_, _23835_, _23833_);
  and _46928_ (_23836_, _00860_, _00922_);
  and _46929_ (_23837_, _23821_, _23836_);
  and _46930_ (_23838_, _23837_, _05518_);
  not _46931_ (_23839_, _23838_);
  nor _46932_ (_23840_, _23839_, _02280_);
  nor _46933_ (_23841_, _23827_, _23822_);
  not _46934_ (_23842_, _23841_);
  nor _46935_ (_23843_, _23837_, _23842_);
  or _46936_ (_23844_, _23843_, _23830_);
  and _46937_ (_23845_, _23844_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nand _46938_ (_23846_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _46939_ (_23847_, _23846_, _23841_);
  or _46940_ (_23848_, _23847_, _23845_);
  or _46941_ (_23849_, _23848_, _23840_);
  and _46942_ (_06422_, _23849_, _25365_);
  and _46943_ (_23850_, _23821_, _04675_);
  and _46944_ (_23851_, _23850_, _05518_);
  not _46945_ (_23852_, _23851_);
  nor _46946_ (_23853_, _23852_, _02280_);
  and _46947_ (_23854_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _46948_ (_23855_, _23854_, _23853_);
  and _46949_ (_06423_, _23855_, _25365_);
  and _46950_ (_23856_, _05516_, _02680_);
  and _46951_ (_23857_, _23856_, _02783_);
  and _46952_ (_23858_, _23857_, _05518_);
  not _46953_ (_23859_, _23858_);
  nor _46954_ (_23860_, _23859_, _02280_);
  and _46955_ (_23861_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or _46956_ (_23862_, _23861_, _23860_);
  and _46957_ (_06424_, _23862_, _25365_);
  and _46958_ (_23863_, _23856_, _02982_);
  and _46959_ (_23864_, _23863_, _05518_);
  not _46960_ (_23865_, _23864_);
  nor _46961_ (_23866_, _23865_, _02280_);
  not _46962_ (_23867_, _23850_);
  nor _46963_ (_23868_, _23863_, _23857_);
  and _46964_ (_23869_, _23868_, _23867_);
  and _46965_ (_23870_, _23869_, _23843_);
  or _46966_ (_23871_, _23870_, _23830_);
  or _46967_ (_23872_, _23850_, _23837_);
  or _46968_ (_23873_, _23857_, _23872_);
  and _46969_ (_23874_, _23873_, _05518_);
  or _46970_ (_23875_, _23874_, _23842_);
  or _46971_ (_23876_, _23875_, _23871_);
  and _46972_ (_23877_, _23876_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or _46973_ (_23878_, _23877_, _23866_);
  and _46974_ (_06425_, _23878_, _25365_);
  and _46975_ (_23879_, _23856_, _23836_);
  and _46976_ (_23880_, _23879_, _05518_);
  not _46977_ (_23881_, _23880_);
  and _46978_ (_23882_, _23881_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _46979_ (_23883_, _23881_, _02280_);
  or _46980_ (_23884_, _23883_, _23882_);
  and _46981_ (_06426_, _23884_, _25365_);
  and _46982_ (_23885_, _23856_, _04675_);
  and _46983_ (_23886_, _23885_, _05557_);
  not _46984_ (_23887_, _23879_);
  and _46985_ (_23888_, _23887_, _23868_);
  not _46986_ (_23889_, _23888_);
  nor _46987_ (_23890_, _23885_, _23879_);
  and _46988_ (_23891_, _23890_, _23870_);
  nor _46989_ (_23892_, _23872_, _23842_);
  nand _46990_ (_23893_, _23892_, _05518_);
  or _46991_ (_23894_, _23893_, _23891_);
  or _46992_ (_23895_, _23894_, _23889_);
  and _46993_ (_23896_, _23895_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or _46994_ (_23897_, _23896_, _23886_);
  or _46995_ (_23898_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _46996_ (_23899_, _23898_, _25365_);
  and _46997_ (_06427_, _23899_, _23897_);
  nand _46998_ (_23900_, _23823_, _02259_);
  or _46999_ (_23901_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _47000_ (_23902_, _23901_, _25365_);
  and _47001_ (_06438_, _23902_, _23900_);
  not _47002_ (_23903_, _23823_);
  or _47003_ (_23904_, _23903_, _02251_);
  or _47004_ (_23905_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _47005_ (_23906_, _23905_, _25365_);
  and _47006_ (_06439_, _23906_, _23904_);
  or _47007_ (_23907_, _23903_, _02236_);
  or _47008_ (_23908_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _47009_ (_23909_, _23908_, _25365_);
  and _47010_ (_06440_, _23909_, _23907_);
  or _47011_ (_23910_, _23903_, _02220_);
  or _47012_ (_23911_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _47013_ (_23912_, _23911_, _25365_);
  and _47014_ (_06441_, _23912_, _23910_);
  nand _47015_ (_23913_, _23823_, _02204_);
  or _47016_ (_23914_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _47017_ (_23915_, _23914_, _25365_);
  and _47018_ (_06442_, _23915_, _23913_);
  nand _47019_ (_23916_, _23823_, _02190_);
  or _47020_ (_23917_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _47021_ (_23918_, _23917_, _25365_);
  and _47022_ (_06443_, _23918_, _23916_);
  nand _47023_ (_23919_, _23823_, _02177_);
  or _47024_ (_23920_, _23823_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _47025_ (_23921_, _23920_, _25365_);
  and _47026_ (_06444_, _23921_, _23919_);
  and _47027_ (_23922_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _47028_ (_23923_, _23827_, _02260_);
  or _47029_ (_23924_, _23923_, _23830_);
  or _47030_ (_23925_, _23924_, _23922_);
  or _47031_ (_23926_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _47032_ (_23927_, _23926_, _25365_);
  and _47033_ (_06445_, _23927_, _23925_);
  and _47034_ (_23928_, _23827_, _02251_);
  and _47035_ (_23929_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _47036_ (_23930_, _23929_, _23830_);
  or _47037_ (_23931_, _23930_, _23928_);
  or _47038_ (_23932_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _47039_ (_23933_, _23932_, _25365_);
  and _47040_ (_06446_, _23933_, _23931_);
  and _47041_ (_23934_, _23827_, _02236_);
  and _47042_ (_23935_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _47043_ (_23936_, _23935_, _23830_);
  or _47044_ (_23937_, _23936_, _23934_);
  or _47045_ (_23938_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _47046_ (_23939_, _23938_, _25365_);
  and _47047_ (_06447_, _23939_, _23937_);
  and _47048_ (_23940_, _23827_, _02220_);
  and _47049_ (_23941_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _47050_ (_23942_, _23941_, _23830_);
  or _47051_ (_23943_, _23942_, _23940_);
  or _47052_ (_23944_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _47053_ (_23945_, _23944_, _25365_);
  and _47054_ (_06448_, _23945_, _23943_);
  nor _47055_ (_23946_, _23828_, _02204_);
  and _47056_ (_23947_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _47057_ (_23948_, _23947_, _23830_);
  or _47058_ (_23949_, _23948_, _23946_);
  or _47059_ (_23950_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _47060_ (_23951_, _23950_, _25365_);
  and _47061_ (_06449_, _23951_, _23949_);
  nor _47062_ (_23952_, _23828_, _02190_);
  and _47063_ (_23953_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _47064_ (_23954_, _23953_, _23830_);
  or _47065_ (_23955_, _23954_, _23952_);
  or _47066_ (_23956_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _47067_ (_23957_, _23956_, _25365_);
  and _47068_ (_06450_, _23957_, _23955_);
  nor _47069_ (_23958_, _23828_, _02177_);
  and _47070_ (_23959_, _23828_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _47071_ (_23960_, _23959_, _23830_);
  or _47072_ (_23961_, _23960_, _23958_);
  or _47073_ (_23962_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _47074_ (_23963_, _23962_, _25365_);
  and _47075_ (_06451_, _23963_, _23961_);
  and _47076_ (_23964_, _23844_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand _47077_ (_23965_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _47078_ (_23966_, _23965_, _23841_);
  and _47079_ (_23967_, _23838_, _02260_);
  or _47080_ (_23968_, _23967_, _23966_);
  or _47081_ (_23969_, _23968_, _23964_);
  and _47082_ (_06452_, _23969_, _25365_);
  and _47083_ (_23970_, _23838_, _02251_);
  and _47084_ (_23971_, _23844_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nand _47085_ (_23972_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _47086_ (_23973_, _23972_, _23841_);
  or _47087_ (_23974_, _23973_, _23971_);
  or _47088_ (_23975_, _23974_, _23970_);
  and _47089_ (_06453_, _23975_, _25365_);
  or _47090_ (_23976_, _23839_, _02236_);
  or _47091_ (_23977_, _23838_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _47092_ (_23978_, _23977_, _25365_);
  and _47093_ (_06454_, _23978_, _23976_);
  and _47094_ (_23979_, _23838_, _02220_);
  and _47095_ (_23980_, _23839_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _47096_ (_23981_, _23980_, _23979_);
  and _47097_ (_06455_, _23981_, _25365_);
  nand _47098_ (_23982_, _23838_, _02204_);
  or _47099_ (_23983_, _23838_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _47100_ (_23984_, _23983_, _25365_);
  and _47101_ (_06456_, _23984_, _23982_);
  nor _47102_ (_23985_, _23839_, _02190_);
  and _47103_ (_23986_, _23839_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _47104_ (_23987_, _23986_, _23985_);
  and _47105_ (_06457_, _23987_, _25365_);
  nor _47106_ (_23988_, _23839_, _02177_);
  and _47107_ (_23989_, _23839_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _47108_ (_23990_, _23989_, _23988_);
  and _47109_ (_06458_, _23990_, _25365_);
  and _47110_ (_23991_, _23851_, _02260_);
  and _47111_ (_23992_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _47112_ (_23993_, _23992_, _23991_);
  and _47113_ (_06459_, _23993_, _25365_);
  and _47114_ (_23994_, _23851_, _02251_);
  and _47115_ (_23995_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _47116_ (_23996_, _23995_, _23994_);
  and _47117_ (_06460_, _23996_, _25365_);
  and _47118_ (_23997_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _47119_ (_23998_, _23851_, _02236_);
  or _47120_ (_23999_, _23998_, _23997_);
  and _47121_ (_06461_, _23999_, _25365_);
  and _47122_ (_24000_, _23851_, _02220_);
  and _47123_ (_24001_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _47124_ (_24002_, _24001_, _24000_);
  and _47125_ (_06462_, _24002_, _25365_);
  and _47126_ (_24003_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _47127_ (_24004_, _23852_, _02204_);
  or _47128_ (_24005_, _24004_, _24003_);
  and _47129_ (_06463_, _24005_, _25365_);
  nor _47130_ (_24006_, _23852_, _02190_);
  and _47131_ (_24007_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _47132_ (_24008_, _24007_, _24006_);
  and _47133_ (_06464_, _24008_, _25365_);
  nor _47134_ (_24009_, _23852_, _02177_);
  and _47135_ (_24010_, _23852_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _47136_ (_24011_, _24010_, _24009_);
  and _47137_ (_06465_, _24011_, _25365_);
  and _47138_ (_24012_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _47139_ (_24013_, _23858_, _02260_);
  or _47140_ (_24014_, _24013_, _24012_);
  and _47141_ (_06466_, _24014_, _25365_);
  and _47142_ (_24015_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _47143_ (_24016_, _23858_, _02251_);
  or _47144_ (_24017_, _24016_, _24015_);
  and _47145_ (_06467_, _24017_, _25365_);
  and _47146_ (_24018_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _47147_ (_24019_, _23858_, _02236_);
  or _47148_ (_24020_, _24019_, _24018_);
  and _47149_ (_06468_, _24020_, _25365_);
  and _47150_ (_24021_, _23858_, _02220_);
  and _47151_ (_24022_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or _47152_ (_24023_, _24022_, _24021_);
  and _47153_ (_06469_, _24023_, _25365_);
  nor _47154_ (_24024_, _23859_, _02204_);
  and _47155_ (_24025_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or _47156_ (_24026_, _24025_, _24024_);
  and _47157_ (_06470_, _24026_, _25365_);
  nor _47158_ (_24027_, _23859_, _02190_);
  and _47159_ (_24028_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _47160_ (_24029_, _24028_, _24027_);
  and _47161_ (_06471_, _24029_, _25365_);
  nor _47162_ (_24030_, _23859_, _02177_);
  and _47163_ (_24031_, _23859_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or _47164_ (_24032_, _24031_, _24030_);
  and _47165_ (_06472_, _24032_, _25365_);
  and _47166_ (_24033_, _23864_, _02260_);
  and _47167_ (_24034_, _23865_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  or _47168_ (_24035_, _24034_, _24033_);
  and _47169_ (_06473_, _24035_, _25365_);
  and _47170_ (_24036_, _23865_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _47171_ (_24037_, _23864_, _02251_);
  or _47172_ (_24038_, _24037_, _24036_);
  and _47173_ (_06474_, _24038_, _25365_);
  and _47174_ (_24039_, _23864_, _02236_);
  and _47175_ (_24040_, _23865_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or _47176_ (_24041_, _24040_, _24039_);
  and _47177_ (_06475_, _24041_, _25365_);
  and _47178_ (_24042_, _23864_, _02220_);
  and _47179_ (_24043_, _23876_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or _47180_ (_24044_, _24043_, _24042_);
  and _47181_ (_06476_, _24044_, _25365_);
  nor _47182_ (_24045_, _23865_, _02204_);
  and _47183_ (_24046_, _23876_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or _47184_ (_24047_, _24046_, _24045_);
  and _47185_ (_06477_, _24047_, _25365_);
  nor _47186_ (_24048_, _23865_, _02190_);
  and _47187_ (_24049_, _23865_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or _47188_ (_24050_, _24049_, _24048_);
  and _47189_ (_06478_, _24050_, _25365_);
  nor _47190_ (_24051_, _23865_, _02177_);
  and _47191_ (_24052_, _23876_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _47192_ (_24053_, _24052_, _24051_);
  and _47193_ (_06479_, _24053_, _25365_);
  and _47194_ (_24054_, _23880_, _02260_);
  and _47195_ (_24055_, _23881_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or _47196_ (_24056_, _24055_, _24054_);
  and _47197_ (_06480_, _24056_, _25365_);
  nand _47198_ (_24057_, _23881_, _23871_);
  nand _47199_ (_24058_, _24057_, _23843_);
  and _47200_ (_24059_, _24058_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _47201_ (_24060_, _23880_, _02251_);
  nand _47202_ (_24061_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _47203_ (_24062_, _24061_, _23869_);
  or _47204_ (_24063_, _24062_, _24060_);
  or _47205_ (_24064_, _24063_, _24059_);
  and _47206_ (_06481_, _24064_, _25365_);
  and _47207_ (_24065_, _23880_, _02236_);
  and _47208_ (_24066_, _23881_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _47209_ (_24067_, _24066_, _24065_);
  and _47210_ (_06482_, _24067_, _25365_);
  and _47211_ (_24068_, _23880_, _02220_);
  and _47212_ (_24069_, _23881_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or _47213_ (_24070_, _24069_, _24068_);
  and _47214_ (_06483_, _24070_, _25365_);
  nor _47215_ (_24071_, _23881_, _02204_);
  and _47216_ (_24072_, _23881_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or _47217_ (_24073_, _24072_, _24071_);
  and _47218_ (_06484_, _24073_, _25365_);
  nor _47219_ (_24074_, _23881_, _02190_);
  and _47220_ (_24075_, _23881_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _47221_ (_24076_, _24075_, _24074_);
  and _47222_ (_06486_, _24076_, _25365_);
  nor _47223_ (_24077_, _23881_, _02177_);
  and _47224_ (_24078_, _23881_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _47225_ (_24079_, _24078_, _24077_);
  and _47226_ (_06487_, _24079_, _25365_);
  and _47227_ (_24080_, _23894_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _47228_ (_24081_, _23885_, _05518_);
  and _47229_ (_24082_, _24081_, _02260_);
  nand _47230_ (_24083_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _47231_ (_24084_, _24083_, _23888_);
  or _47232_ (_24085_, _24084_, _24082_);
  or _47233_ (_24086_, _24085_, _24080_);
  and _47234_ (_06488_, _24086_, _25365_);
  and _47235_ (_24087_, _23895_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _47236_ (_24088_, _24081_, _02251_);
  or _47237_ (_24089_, _24088_, _24087_);
  and _47238_ (_06489_, _24089_, _25365_);
  and _47239_ (_24090_, _23894_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and _47240_ (_24091_, _24081_, _02236_);
  nand _47241_ (_24092_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _47242_ (_24093_, _24092_, _23888_);
  or _47243_ (_24094_, _24093_, _24091_);
  or _47244_ (_24095_, _24094_, _24090_);
  and _47245_ (_06490_, _24095_, _25365_);
  and _47246_ (_24096_, _23894_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _47247_ (_24097_, _24081_, _02220_);
  nand _47248_ (_24098_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _47249_ (_24099_, _24098_, _23888_);
  or _47250_ (_24100_, _24099_, _24097_);
  or _47251_ (_24101_, _24100_, _24096_);
  and _47252_ (_06491_, _24101_, _25365_);
  and _47253_ (_24102_, _23895_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _47254_ (_24103_, _24081_, _05765_);
  or _47255_ (_24104_, _24103_, _24102_);
  and _47256_ (_06492_, _24104_, _25365_);
  and _47257_ (_24105_, _23894_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _47258_ (_24106_, _24081_, _03604_);
  nand _47259_ (_24107_, _05518_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _47260_ (_24108_, _24107_, _23888_);
  or _47261_ (_24109_, _24108_, _24106_);
  or _47262_ (_24110_, _24109_, _24105_);
  and _47263_ (_06493_, _24110_, _25365_);
  and _47264_ (_24111_, _24081_, _03628_);
  nor _47265_ (_24112_, _23888_, _23830_);
  or _47266_ (_24113_, _24112_, _23894_);
  and _47267_ (_24114_, _24113_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or _47268_ (_24115_, _24114_, _24111_);
  and _47269_ (_06494_, _24115_, _25365_);
  not _47270_ (_24116_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _47271_ (_24117_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and _47272_ (_24118_, _24117_, _24116_);
  and _47273_ (_24119_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _25365_);
  and _47274_ (_06501_, _24119_, _24118_);
  nor _47275_ (_24120_, _24118_, rst);
  nand _47276_ (_24121_, _24117_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _47277_ (_24122_, _24117_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _47278_ (_24123_, _24122_, _24121_);
  and _47279_ (_06502_, _24123_, _24120_);
  nor _47280_ (_24124_, _05867_, _05821_);
  and _47281_ (_24125_, _05775_, _06020_);
  and _47282_ (_24126_, _24125_, _24124_);
  and _47283_ (_24127_, _24126_, _05653_);
  and _47284_ (_24128_, _24127_, _02782_);
  nor _47285_ (_24129_, _24128_, _22374_);
  not _47286_ (_24130_, _05720_);
  nor _47287_ (_24131_, _24130_, _05994_);
  and _47288_ (_24132_, _24131_, _03628_);
  or _47289_ (_24133_, _24132_, _05918_);
  and _47290_ (_24134_, _05720_, _05994_);
  and _47291_ (_24135_, _24134_, _05765_);
  and _47292_ (_24136_, _24130_, _05994_);
  and _47293_ (_24137_, _24136_, _03604_);
  nor _47294_ (_24138_, _05720_, _05994_);
  and _47295_ (_24139_, _24138_, _05557_);
  or _47296_ (_24140_, _24139_, _24137_);
  or _47297_ (_24141_, _24140_, _24135_);
  or _47298_ (_24142_, _24141_, _24133_);
  not _47299_ (_24143_, _05918_);
  and _47300_ (_24144_, _24131_, _02236_);
  or _47301_ (_24145_, _24144_, _24143_);
  and _47302_ (_24146_, _24134_, _02260_);
  and _47303_ (_24147_, _24136_, _02251_);
  and _47304_ (_24148_, _24138_, _02220_);
  or _47305_ (_24149_, _24148_, _24147_);
  or _47306_ (_24150_, _24149_, _24146_);
  or _47307_ (_24151_, _24150_, _24145_);
  nand _47308_ (_24152_, _24151_, _24142_);
  nor _47309_ (_24153_, _24152_, _24129_);
  not _47310_ (_24154_, _05867_);
  and _47311_ (_24155_, _24154_, _05821_);
  nor _47312_ (_24156_, _05775_, _05584_);
  and _47313_ (_24157_, _24156_, _05653_);
  and _47314_ (_24158_, _24157_, _24155_);
  nand _47315_ (_24159_, _02847_, _02845_);
  nand _47316_ (_24160_, _02863_, _24159_);
  or _47317_ (_24161_, _02863_, _24159_);
  nand _47318_ (_24162_, _24161_, _24160_);
  not _47319_ (_24163_, _02835_);
  nand _47320_ (_24164_, _24163_, _02822_);
  or _47321_ (_24165_, _24163_, _02822_);
  nand _47322_ (_24166_, _24165_, _24164_);
  nand _47323_ (_24167_, _24166_, _24162_);
  or _47324_ (_24168_, _24166_, _24162_);
  nand _47325_ (_24169_, _24168_, _24167_);
  or _47326_ (_24170_, _02889_, _02876_);
  nand _47327_ (_24171_, _02889_, _02876_);
  nand _47328_ (_24172_, _24171_, _24170_);
  nand _47329_ (_24173_, _02901_, _02899_);
  nand _47330_ (_24174_, _24173_, _02810_);
  or _47331_ (_24175_, _24173_, _02810_);
  and _47332_ (_24176_, _24175_, _24174_);
  nand _47333_ (_24177_, _24176_, _24172_);
  or _47334_ (_24178_, _24176_, _24172_);
  nand _47335_ (_24179_, _24178_, _24177_);
  nand _47336_ (_24180_, _24179_, _24169_);
  or _47337_ (_24181_, _24179_, _24169_);
  nand _47338_ (_24182_, _24181_, _24180_);
  nand _47339_ (_24183_, _24182_, _05918_);
  or _47340_ (_24184_, _05918_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _47341_ (_24185_, _24184_, _24134_);
  and _47342_ (_24186_, _24185_, _24183_);
  and _47343_ (_24187_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _47344_ (_24188_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _47345_ (_24189_, _24188_, _24187_);
  and _47346_ (_24190_, _24189_, _24143_);
  nor _47347_ (_24191_, _05918_, _02670_);
  and _47348_ (_24192_, _05918_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _47349_ (_24193_, _24192_, _24191_);
  and _47350_ (_24194_, _24193_, _24138_);
  and _47351_ (_24195_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _47352_ (_24196_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _47353_ (_24197_, _24196_, _24195_);
  and _47354_ (_24198_, _24197_, _05918_);
  or _47355_ (_24199_, _24198_, _24194_);
  or _47356_ (_24200_, _24199_, _24190_);
  or _47357_ (_24201_, _24200_, _24186_);
  and _47358_ (_24202_, _24201_, _24158_);
  nor _47359_ (_24203_, _24154_, _05821_);
  nor _47360_ (_24204_, _21795_, _02016_);
  and _47361_ (_24205_, _24204_, _21851_);
  and _47362_ (_24206_, _02125_, _02006_);
  or _47363_ (_24207_, _24206_, _02069_);
  nor _47364_ (_24208_, _21978_, _24207_);
  and _47365_ (_24209_, _02118_, _01993_);
  or _47366_ (_24210_, _24209_, _02023_);
  nor _47367_ (_24211_, _24210_, _02104_);
  and _47368_ (_24212_, _02046_, _01948_);
  or _47369_ (_24213_, _24212_, _21796_);
  or _47370_ (_24214_, _24213_, _21869_);
  nor _47371_ (_24215_, _24214_, _21753_);
  and _47372_ (_24216_, _24215_, _24211_);
  and _47373_ (_24217_, _24216_, _24208_);
  and _47374_ (_24218_, _24217_, _24205_);
  and _47375_ (_24219_, _24218_, _02062_);
  nor _47376_ (_24220_, _24219_, _02140_);
  or _47377_ (_24221_, _24220_, p3_in[2]);
  not _47378_ (_24222_, _24220_);
  or _47379_ (_24223_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _47380_ (_24224_, _24223_, _24221_);
  and _47381_ (_24225_, _24224_, _24131_);
  nor _47382_ (_24226_, _24220_, p3_in[0]);
  and _47383_ (_24227_, _24220_, _03259_);
  nor _47384_ (_24228_, _24227_, _24226_);
  and _47385_ (_24229_, _24228_, _24134_);
  or _47386_ (_24230_, _24229_, _24225_);
  or _47387_ (_24231_, _24220_, p3_in[3]);
  or _47388_ (_24232_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _47389_ (_24233_, _24232_, _24231_);
  and _47390_ (_24234_, _24233_, _24138_);
  nor _47391_ (_24235_, _24220_, p3_in[1]);
  and _47392_ (_24236_, _24220_, _03272_);
  nor _47393_ (_24237_, _24236_, _24235_);
  and _47394_ (_24238_, _24237_, _24136_);
  or _47395_ (_24239_, _24238_, _24234_);
  or _47396_ (_24240_, _24239_, _24230_);
  and _47397_ (_24241_, _24240_, _05918_);
  nor _47398_ (_24242_, _24220_, p3_in[6]);
  and _47399_ (_24243_, _24220_, _03334_);
  nor _47400_ (_24244_, _24243_, _24242_);
  and _47401_ (_24245_, _24244_, _24131_);
  or _47402_ (_24246_, _24220_, p3_in[4]);
  or _47403_ (_24247_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47404_ (_24248_, _24247_, _24246_);
  and _47405_ (_24249_, _24248_, _24134_);
  or _47406_ (_24250_, _24249_, _24245_);
  or _47407_ (_24251_, _24220_, p3_in[7]);
  or _47408_ (_24252_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _47409_ (_24253_, _24252_, _24251_);
  and _47410_ (_24254_, _24253_, _24138_);
  or _47411_ (_24255_, _24220_, p3_in[5]);
  or _47412_ (_24256_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _47413_ (_24257_, _24256_, _24255_);
  and _47414_ (_24258_, _24257_, _24136_);
  or _47415_ (_24259_, _24258_, _24254_);
  or _47416_ (_24260_, _24259_, _24250_);
  and _47417_ (_24261_, _24260_, _24143_);
  or _47418_ (_24262_, _24261_, _24241_);
  and _47419_ (_24263_, _24262_, _24203_);
  and _47420_ (_24264_, _05867_, _05821_);
  nor _47421_ (_24265_, _24220_, p1_in[1]);
  and _47422_ (_24266_, _24220_, _03096_);
  nor _47423_ (_24267_, _24266_, _24265_);
  and _47424_ (_24268_, _24267_, _24136_);
  nor _47425_ (_24269_, _24220_, p1_in[0]);
  and _47426_ (_24270_, _24220_, _03081_);
  nor _47427_ (_24271_, _24270_, _24269_);
  and _47428_ (_24272_, _24271_, _24134_);
  or _47429_ (_24273_, _24272_, _24268_);
  or _47430_ (_24274_, _24220_, p1_in[2]);
  or _47431_ (_24275_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _47432_ (_24276_, _24275_, _24274_);
  and _47433_ (_24277_, _24276_, _24131_);
  or _47434_ (_24278_, _24220_, p1_in[3]);
  or _47435_ (_24279_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _47436_ (_24280_, _24279_, _24278_);
  and _47437_ (_24281_, _24280_, _24138_);
  or _47438_ (_24282_, _24281_, _24277_);
  or _47439_ (_24283_, _24282_, _24273_);
  and _47440_ (_24284_, _24283_, _05918_);
  or _47441_ (_24285_, _24220_, p1_in[5]);
  or _47442_ (_24286_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _47443_ (_24287_, _24286_, _24285_);
  and _47444_ (_24288_, _24287_, _24136_);
  or _47445_ (_24289_, _24220_, p1_in[4]);
  or _47446_ (_24290_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47447_ (_24291_, _24290_, _24289_);
  and _47448_ (_24292_, _24291_, _24134_);
  or _47449_ (_24293_, _24292_, _24288_);
  nor _47450_ (_24294_, _24220_, p1_in[6]);
  and _47451_ (_24295_, _24220_, _03162_);
  nor _47452_ (_24296_, _24295_, _24294_);
  and _47453_ (_24297_, _24296_, _24131_);
  or _47454_ (_24298_, _24220_, p1_in[7]);
  or _47455_ (_24299_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _47456_ (_24300_, _24299_, _24298_);
  and _47457_ (_24301_, _24300_, _24138_);
  or _47458_ (_24302_, _24301_, _24297_);
  or _47459_ (_24303_, _24302_, _24293_);
  and _47460_ (_24304_, _24303_, _24143_);
  or _47461_ (_24305_, _24304_, _24284_);
  and _47462_ (_24306_, _24305_, _24264_);
  and _47463_ (_24307_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _47464_ (_24308_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _47465_ (_24309_, _24308_, _24307_);
  and _47466_ (_24310_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _47467_ (_24311_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _47468_ (_24312_, _24311_, _24310_);
  or _47469_ (_24313_, _24312_, _24309_);
  and _47470_ (_24314_, _24313_, _24143_);
  and _47471_ (_24315_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _47472_ (_24316_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _47473_ (_24317_, _24316_, _24315_);
  and _47474_ (_24318_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _47475_ (_24319_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _47476_ (_24320_, _24319_, _24318_);
  or _47477_ (_24321_, _24320_, _24317_);
  and _47478_ (_24322_, _24321_, _05918_);
  or _47479_ (_24323_, _24322_, _24314_);
  and _47480_ (_24324_, _24323_, _24124_);
  or _47481_ (_24325_, _24324_, _24306_);
  or _47482_ (_24326_, _24325_, _24263_);
  and _47483_ (_24327_, _24326_, _24157_);
  not _47484_ (_24328_, _05653_);
  and _47485_ (_24329_, _24125_, _24328_);
  and _47486_ (_24330_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _47487_ (_24331_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _47488_ (_24332_, _24331_, _24330_);
  and _47489_ (_24333_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47490_ (_24334_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _47491_ (_24335_, _24334_, _24333_);
  or _47492_ (_24336_, _24335_, _24332_);
  and _47493_ (_24337_, _24336_, _24203_);
  and _47494_ (_24338_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _47495_ (_24339_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _47496_ (_24340_, _24339_, _24338_);
  and _47497_ (_24341_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _47498_ (_24342_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _47499_ (_24343_, _24342_, _24341_);
  or _47500_ (_24344_, _24343_, _24340_);
  and _47501_ (_24345_, _24344_, _24264_);
  or _47502_ (_24346_, _24345_, _24337_);
  and _47503_ (_24347_, _24346_, _05918_);
  and _47504_ (_24348_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _47505_ (_24349_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _47506_ (_24350_, _24349_, _24348_);
  and _47507_ (_24351_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _47508_ (_24352_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _47509_ (_24353_, _24352_, _24351_);
  or _47510_ (_24354_, _24353_, _24350_);
  and _47511_ (_24355_, _24354_, _24264_);
  and _47512_ (_24356_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _47513_ (_24357_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _47514_ (_24358_, _24357_, _24356_);
  and _47515_ (_24359_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _47516_ (_24360_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _47517_ (_24361_, _24360_, _24359_);
  or _47518_ (_24362_, _24361_, _24358_);
  and _47519_ (_24363_, _24362_, _24203_);
  or _47520_ (_24364_, _24363_, _24355_);
  and _47521_ (_24365_, _24364_, _24143_);
  or _47522_ (_24366_, _24365_, _24347_);
  and _47523_ (_24367_, _24366_, _24329_);
  and _47524_ (_24368_, _24264_, _24125_);
  and _47525_ (_24369_, _24368_, _05653_);
  or _47526_ (_24370_, _24220_, p0_in[5]);
  or _47527_ (_24371_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _47528_ (_24372_, _24371_, _24370_);
  and _47529_ (_24373_, _24372_, _24136_);
  or _47530_ (_24374_, _24220_, p0_in[7]);
  or _47531_ (_24375_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _47532_ (_24376_, _24375_, _24374_);
  and _47533_ (_24377_, _24376_, _24138_);
  or _47534_ (_24378_, _24377_, _24373_);
  nor _47535_ (_24379_, _24220_, p0_in[6]);
  and _47536_ (_24380_, _24220_, _03067_);
  nor _47537_ (_24381_, _24380_, _24379_);
  and _47538_ (_24382_, _24381_, _24131_);
  or _47539_ (_24383_, _24220_, p0_in[4]);
  or _47540_ (_24384_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _47541_ (_24385_, _24384_, _24383_);
  and _47542_ (_24386_, _24385_, _24134_);
  or _47543_ (_24387_, _24386_, _24382_);
  or _47544_ (_24388_, _24387_, _24378_);
  and _47545_ (_24389_, _24388_, _24143_);
  nor _47546_ (_24390_, _24220_, p0_in[1]);
  and _47547_ (_24391_, _24220_, _02994_);
  nor _47548_ (_24392_, _24391_, _24390_);
  and _47549_ (_24393_, _24392_, _24136_);
  or _47550_ (_24394_, _24220_, p0_in[3]);
  or _47551_ (_24395_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _47552_ (_24396_, _24395_, _24394_);
  and _47553_ (_24397_, _24396_, _24138_);
  or _47554_ (_24398_, _24397_, _24393_);
  or _47555_ (_24399_, _24220_, p0_in[2]);
  or _47556_ (_24400_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _47557_ (_24401_, _24400_, _24399_);
  and _47558_ (_24402_, _24401_, _24131_);
  nor _47559_ (_24403_, _24220_, p0_in[0]);
  and _47560_ (_24404_, _24220_, _02977_);
  nor _47561_ (_24405_, _24404_, _24403_);
  and _47562_ (_24406_, _24405_, _24134_);
  or _47563_ (_24407_, _24406_, _24402_);
  or _47564_ (_24408_, _24407_, _24398_);
  and _47565_ (_24409_, _24408_, _05918_);
  or _47566_ (_24410_, _24409_, _24389_);
  and _47567_ (_24411_, _24410_, _24369_);
  and _47568_ (_24412_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _47569_ (_24413_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _47570_ (_24414_, _24413_, _24412_);
  and _47571_ (_24415_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _47572_ (_24416_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _47573_ (_24417_, _24416_, _24415_);
  or _47574_ (_24418_, _24417_, _24414_);
  and _47575_ (_24419_, _24418_, _05918_);
  and _47576_ (_24420_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _47577_ (_24421_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _47578_ (_24422_, _24421_, _24420_);
  and _47579_ (_24423_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _47580_ (_24424_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _47581_ (_24425_, _24424_, _24423_);
  or _47582_ (_24426_, _24425_, _24422_);
  and _47583_ (_24427_, _24426_, _24143_);
  or _47584_ (_24428_, _24427_, _24419_);
  and _47585_ (_24429_, _24428_, _24127_);
  or _47586_ (_24430_, _24429_, _24411_);
  and _47587_ (_24431_, _22389_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _47588_ (_24432_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _47589_ (_24433_, _24432_, _05918_);
  and _47590_ (_24434_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _47591_ (_24435_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _47592_ (_24436_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _47593_ (_24437_, _24436_, _24435_);
  or _47594_ (_24438_, _24437_, _24434_);
  or _47595_ (_24439_, _24438_, _24433_);
  and _47596_ (_24440_, _24156_, _24328_);
  and _47597_ (_24441_, _24440_, _24203_);
  and _47598_ (_24442_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _47599_ (_24443_, _24442_, _24143_);
  and _47600_ (_24444_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _47601_ (_24445_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47602_ (_24446_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _47603_ (_24447_, _24446_, _24445_);
  or _47604_ (_24448_, _24447_, _24444_);
  or _47605_ (_24449_, _24448_, _24443_);
  and _47606_ (_24450_, _24449_, _24441_);
  and _47607_ (_24451_, _24450_, _24439_);
  or _47608_ (_24452_, _24451_, _24431_);
  or _47609_ (_24453_, _24452_, _24430_);
  or _47610_ (_24454_, _24220_, p2_in[5]);
  or _47611_ (_24455_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _47612_ (_24456_, _24455_, _24454_);
  and _47613_ (_24457_, _24456_, _24136_);
  or _47614_ (_24458_, _24457_, _05918_);
  or _47615_ (_24459_, _24220_, p2_in[4]);
  or _47616_ (_24460_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _47617_ (_24461_, _24460_, _24459_);
  and _47618_ (_24462_, _24461_, _24134_);
  or _47619_ (_24463_, _24220_, p2_in[7]);
  or _47620_ (_24464_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _47621_ (_24465_, _24464_, _24463_);
  and _47622_ (_24466_, _24465_, _24138_);
  nor _47623_ (_24467_, _24220_, p2_in[6]);
  and _47624_ (_24468_, _24220_, _03246_);
  nor _47625_ (_24469_, _24468_, _24467_);
  and _47626_ (_24470_, _24469_, _24131_);
  or _47627_ (_24471_, _24470_, _24466_);
  or _47628_ (_24472_, _24471_, _24462_);
  or _47629_ (_24473_, _24472_, _24458_);
  and _47630_ (_24474_, _24203_, _24125_);
  and _47631_ (_24475_, _24474_, _05653_);
  nor _47632_ (_24476_, _24220_, p2_in[1]);
  and _47633_ (_24477_, _24220_, _03185_);
  nor _47634_ (_24478_, _24477_, _24476_);
  and _47635_ (_24479_, _24478_, _24136_);
  or _47636_ (_24480_, _24479_, _24143_);
  nor _47637_ (_24481_, _24220_, p2_in[0]);
  and _47638_ (_24482_, _24220_, _03172_);
  nor _47639_ (_24483_, _24482_, _24481_);
  and _47640_ (_24484_, _24483_, _24134_);
  or _47641_ (_24485_, _24220_, p2_in[3]);
  or _47642_ (_24486_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _47643_ (_24487_, _24486_, _24485_);
  and _47644_ (_24488_, _24487_, _24138_);
  or _47645_ (_24489_, _24220_, p2_in[2]);
  or _47646_ (_24490_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _47647_ (_24491_, _24490_, _24489_);
  and _47648_ (_24492_, _24491_, _24131_);
  or _47649_ (_24493_, _24492_, _24488_);
  or _47650_ (_24494_, _24493_, _24484_);
  or _47651_ (_24495_, _24494_, _24480_);
  and _47652_ (_24496_, _24495_, _24475_);
  and _47653_ (_24497_, _24496_, _24473_);
  and _47654_ (_24498_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _47655_ (_24499_, _24498_, _05918_);
  and _47656_ (_24500_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _47657_ (_24501_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _47658_ (_24502_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _47659_ (_24503_, _24502_, _24501_);
  or _47660_ (_24504_, _24503_, _24500_);
  or _47661_ (_24505_, _24504_, _24499_);
  and _47662_ (_24506_, _24440_, _24264_);
  and _47663_ (_24507_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _47664_ (_24508_, _24507_, _24143_);
  and _47665_ (_24509_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _47666_ (_24510_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _47667_ (_24511_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _47668_ (_24512_, _24511_, _24510_);
  or _47669_ (_24513_, _24512_, _24509_);
  or _47670_ (_24514_, _24513_, _24508_);
  and _47671_ (_24515_, _24514_, _24506_);
  and _47672_ (_24516_, _24515_, _24505_);
  or _47673_ (_24517_, _24516_, _24497_);
  and _47674_ (_24518_, _24329_, _24155_);
  and _47675_ (_24519_, _05867_, _06020_);
  nand _47676_ (_24520_, _24519_, _24328_);
  nand _47677_ (_24521_, _24520_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _47678_ (_24522_, _24521_, _24518_);
  nor _47679_ (_24523_, _24369_, _24127_);
  nor _47680_ (_24524_, _24475_, _24157_);
  and _47681_ (_24525_, _24524_, _24523_);
  and _47682_ (_24526_, _24525_, _24522_);
  and _47683_ (_24527_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _47684_ (_24528_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _47685_ (_24529_, _24528_, _24527_);
  and _47686_ (_24530_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _47687_ (_24531_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _47688_ (_24532_, _24531_, _24530_);
  or _47689_ (_24533_, _24532_, _24529_);
  and _47690_ (_24534_, _24533_, _24143_);
  and _47691_ (_24535_, _24131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _47692_ (_24536_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _47693_ (_24537_, _24536_, _24535_);
  and _47694_ (_24538_, _24136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _47695_ (_24539_, _24138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _47696_ (_24540_, _24539_, _24538_);
  or _47697_ (_24541_, _24540_, _24537_);
  and _47698_ (_24542_, _24541_, _05918_);
  or _47699_ (_24543_, _24542_, _24534_);
  and _47700_ (_24544_, _24543_, _24518_);
  or _47701_ (_24545_, _24544_, _24526_);
  or _47702_ (_24546_, _24545_, _24517_);
  or _47703_ (_24547_, _24546_, _24453_);
  or _47704_ (_24548_, _24547_, _24367_);
  or _47705_ (_24549_, _24548_, _24327_);
  or _47706_ (_24550_, _24549_, _24202_);
  nand _47707_ (_24551_, _24431_, _01289_);
  and _47708_ (_24552_, _24551_, _24129_);
  and _47709_ (_24553_, _24552_, _24550_);
  or _47710_ (_24554_, _24553_, _24153_);
  and _47711_ (_06503_, _24554_, _25365_);
  and _47712_ (_24555_, _05653_, _05918_);
  and _47713_ (_24556_, _24555_, _24134_);
  and _47714_ (_24557_, _24556_, _24126_);
  and _47715_ (_24558_, _24557_, _02782_);
  not _47716_ (_24559_, _02796_);
  and _47717_ (_24560_, _24138_, _24143_);
  nor _47718_ (_24561_, _24560_, _24559_);
  and _47719_ (_24562_, _24561_, _22372_);
  nor _47720_ (_24563_, _24562_, _24558_);
  and _47721_ (_24564_, _24563_, _22392_);
  and _47722_ (_24565_, _24555_, _24138_);
  and _47723_ (_24566_, _24565_, _24368_);
  nand _47724_ (_24567_, _24566_, _02328_);
  and _47725_ (_24568_, _24557_, _02792_);
  not _47726_ (_24569_, _05775_);
  and _47727_ (_24570_, _24569_, _05821_);
  nor _47728_ (_24571_, _05867_, _05584_);
  and _47729_ (_24572_, _24556_, _24571_);
  and _47730_ (_24573_, _24572_, _24570_);
  and _47731_ (_24574_, _24573_, _02675_);
  nor _47732_ (_24575_, _24574_, _24568_);
  and _47733_ (_24576_, _24575_, _24567_);
  nor _47734_ (_24577_, _24576_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _47735_ (_24578_, _24577_);
  and _47736_ (_24579_, _24578_, _24564_);
  and _47737_ (_24580_, _24555_, _24131_);
  and _47738_ (_24581_, _24580_, _24368_);
  and _47739_ (_24582_, _24581_, _02328_);
  or _47740_ (_24583_, _24582_, rst);
  nor _47741_ (_06504_, _24583_, _24579_);
  not _47742_ (_24584_, _24579_);
  nand _47743_ (_24585_, _24518_, _24134_);
  and _47744_ (_24586_, _24155_, _24125_);
  nor _47745_ (_24587_, _05653_, _05918_);
  and _47746_ (_24588_, _24587_, _24136_);
  and _47747_ (_24589_, _24588_, _24586_);
  and _47748_ (_24590_, _24328_, _05918_);
  and _47749_ (_24591_, _24590_, _24131_);
  and _47750_ (_24592_, _24591_, _24586_);
  nor _47751_ (_24593_, _24592_, _24589_);
  and _47752_ (_24594_, _24593_, _24585_);
  and _47753_ (_24595_, _24590_, _24134_);
  and _47754_ (_24596_, _24595_, _24368_);
  and _47755_ (_24597_, _24590_, _24138_);
  and _47756_ (_24598_, _24597_, _24586_);
  nor _47757_ (_24599_, _24598_, _24596_);
  and _47758_ (_24600_, _24595_, _24474_);
  nor _47759_ (_24601_, _05775_, _05821_);
  and _47760_ (_24602_, _24601_, _24519_);
  and _47761_ (_24603_, _24560_, _05653_);
  and _47762_ (_24604_, _24603_, _24602_);
  nor _47763_ (_24605_, _24604_, _24600_);
  and _47764_ (_24606_, _24605_, _24599_);
  and _47765_ (_24607_, _24606_, _24594_);
  and _47766_ (_24608_, _24590_, _24136_);
  and _47767_ (_24609_, _24608_, _24368_);
  and _47768_ (_24610_, _24597_, _24368_);
  nor _47769_ (_24611_, _24610_, _24609_);
  and _47770_ (_24612_, _24588_, _24368_);
  and _47771_ (_24613_, _24591_, _24368_);
  nor _47772_ (_24614_, _24613_, _24612_);
  and _47773_ (_24615_, _24614_, _24611_);
  and _47774_ (_24616_, _24587_, _24134_);
  and _47775_ (_24617_, _24616_, _24368_);
  and _47776_ (_24618_, _24603_, _24368_);
  nor _47777_ (_24619_, _24618_, _24617_);
  and _47778_ (_24620_, _24570_, _24519_);
  and _47779_ (_24621_, _24608_, _24620_);
  and _47780_ (_24622_, _24595_, _24620_);
  nor _47781_ (_24623_, _24622_, _24621_);
  and _47782_ (_24624_, _24623_, _24619_);
  and _47783_ (_24625_, _24624_, _24615_);
  and _47784_ (_24626_, _24625_, _24607_);
  and _47785_ (_24627_, _24556_, _24519_);
  nor _47786_ (_24628_, _24581_, _24566_);
  and _47787_ (_24629_, _24555_, _24136_);
  and _47788_ (_24630_, _24629_, _24368_);
  and _47789_ (_24631_, _24601_, _24572_);
  nor _47790_ (_24632_, _24631_, _24630_);
  nand _47791_ (_24633_, _24632_, _24628_);
  nor _47792_ (_24634_, _24633_, _24627_);
  nor _47793_ (_24635_, _24573_, _24557_);
  and _47794_ (_24636_, _24635_, _24634_);
  and _47795_ (_24637_, _24636_, _24626_);
  or _47796_ (_24638_, _24637_, _24584_);
  and _47797_ (_24639_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _47798_ (_24640_, _24616_, _24586_);
  and _47799_ (_24641_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _47800_ (_24642_, _24595_, _24586_);
  and _47801_ (_24643_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _47802_ (_24644_, _24643_, _24641_);
  and _47803_ (_24645_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _47804_ (_24646_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _47805_ (_24647_, _24646_, _24645_);
  or _47806_ (_24648_, _24647_, _24644_);
  and _47807_ (_24649_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _47808_ (_24650_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _47809_ (_24651_, _24650_, _24649_);
  and _47810_ (_24652_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47811_ (_24653_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _47812_ (_24654_, _24653_, _24652_);
  or _47813_ (_24655_, _24654_, _24651_);
  or _47814_ (_24656_, _24655_, _24648_);
  and _47815_ (_24657_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _47816_ (_24658_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _47817_ (_24659_, _24658_, _24657_);
  and _47818_ (_24660_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _47819_ (_24661_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _47820_ (_24662_, _24661_, _24660_);
  or _47821_ (_24663_, _24662_, _24659_);
  and _47822_ (_24664_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _47823_ (_24665_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _47824_ (_24666_, _24665_, _24664_);
  and _47825_ (_24667_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _47826_ (_24668_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _47827_ (_24669_, _24668_, _24667_);
  or _47828_ (_24670_, _24669_, _24666_);
  or _47829_ (_24671_, _24670_, _24663_);
  or _47830_ (_24672_, _24671_, _24656_);
  and _47831_ (_24673_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _47832_ (_24674_, _24630_, _02282_);
  or _47833_ (_24675_, _24674_, _24673_);
  and _47834_ (_24676_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _47835_ (_24677_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _47836_ (_24678_, _24677_, _24676_);
  or _47837_ (_24679_, _24678_, _24675_);
  and _47838_ (_24680_, _24556_, _24368_);
  and _47839_ (_24681_, _24680_, _24376_);
  and _47840_ (_24682_, _24620_, _24556_);
  and _47841_ (_24683_, _24682_, _24300_);
  or _47842_ (_24684_, _24683_, _24681_);
  and _47843_ (_24685_, _24556_, _24474_);
  and _47844_ (_24686_, _24685_, _24465_);
  and _47845_ (_24687_, _24602_, _24556_);
  and _47846_ (_24688_, _24687_, _24253_);
  or _47847_ (_24689_, _24688_, _24686_);
  or _47848_ (_24690_, _24689_, _24684_);
  or _47849_ (_24691_, _24690_, _24679_);
  and _47850_ (_24692_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _47851_ (_24693_, _24573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _47852_ (_24694_, _24693_, _24692_);
  or _47853_ (_24695_, _24694_, _24691_);
  or _47854_ (_24696_, _24695_, _24672_);
  and _47855_ (_24697_, _24696_, _24579_);
  or _47856_ (_24698_, _24697_, _24582_);
  or _47857_ (_24699_, _24698_, _24639_);
  not _47858_ (_24700_, _24582_);
  or _47859_ (_24701_, _24700_, _01184_);
  and _47860_ (_24702_, _24701_, _25365_);
  and _47861_ (_06505_, _24702_, _24699_);
  nor _47862_ (_06515_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _47863_ (_24703_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor _47864_ (_24704_, _24117_, rst);
  and _47865_ (_06516_, _24704_, _24703_);
  nor _47866_ (_24705_, _24117_, _24116_);
  or _47867_ (_24706_, _24705_, _24118_);
  and _47868_ (_24707_, _24121_, _25365_);
  and _47869_ (_06517_, _24707_, _24706_);
  nand _47870_ (_24708_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _47871_ (_24709_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _47872_ (_24710_, _24709_, _24708_);
  nand _47873_ (_24711_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _47874_ (_24712_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _47875_ (_24713_, _24712_, _24711_);
  and _47876_ (_24714_, _24713_, _24710_);
  nand _47877_ (_24715_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _47878_ (_24716_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _47879_ (_24717_, _24716_, _24715_);
  nand _47880_ (_24718_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _47881_ (_24719_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47882_ (_24720_, _24719_, _24718_);
  and _47883_ (_24721_, _24720_, _24717_);
  and _47884_ (_24722_, _24721_, _24714_);
  nand _47885_ (_24723_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand _47886_ (_24724_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47887_ (_24725_, _24724_, _24723_);
  nand _47888_ (_24726_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _47889_ (_24727_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47890_ (_24728_, _24727_, _24726_);
  and _47891_ (_24729_, _24728_, _24725_);
  nand _47892_ (_24730_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _47893_ (_24731_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _47894_ (_24732_, _24731_, _24730_);
  nand _47895_ (_24733_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47896_ (_24734_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _47897_ (_24735_, _24734_, _24733_);
  and _47898_ (_24736_, _24735_, _24732_);
  and _47899_ (_24737_, _24736_, _24729_);
  and _47900_ (_24738_, _24737_, _24722_);
  nand _47901_ (_24739_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand _47902_ (_24740_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _47903_ (_24741_, _24740_, _24739_);
  nand _47904_ (_24742_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _47905_ (_24743_, _24630_);
  or _47906_ (_24744_, _24743_, _02290_);
  and _47907_ (_24745_, _24744_, _24742_);
  and _47908_ (_24746_, _24745_, _24741_);
  nand _47909_ (_24747_, _24685_, _24483_);
  nand _47910_ (_24748_, _24687_, _24228_);
  and _47911_ (_24749_, _24748_, _24747_);
  nand _47912_ (_24750_, _24682_, _24271_);
  nand _47913_ (_24751_, _24680_, _24405_);
  and _47914_ (_24752_, _24751_, _24750_);
  and _47915_ (_24753_, _24752_, _24749_);
  and _47916_ (_24754_, _24753_, _24746_);
  not _47917_ (_24755_, _24573_);
  or _47918_ (_24756_, _24755_, _24182_);
  nand _47919_ (_24757_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _47920_ (_24758_, _24757_, _24756_);
  and _47921_ (_24759_, _24758_, _24754_);
  and _47922_ (_24760_, _24759_, _24738_);
  nor _47923_ (_24761_, _24760_, _24584_);
  nand _47924_ (_24762_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _47925_ (_24763_, _24762_, _24700_);
  or _47926_ (_24764_, _24763_, _24761_);
  or _47927_ (_24765_, _24700_, _01337_);
  and _47928_ (_24766_, _24765_, _25365_);
  and _47929_ (_06518_, _24766_, _24764_);
  and _47930_ (_24767_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _47931_ (_24768_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _47932_ (_24769_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _47933_ (_24770_, _24769_, _24768_);
  nand _47934_ (_24771_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand _47935_ (_24772_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _47936_ (_24773_, _24772_, _24771_);
  and _47937_ (_24774_, _24773_, _24770_);
  nand _47938_ (_24775_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nand _47939_ (_24776_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _47940_ (_24777_, _24776_, _24775_);
  nand _47941_ (_24778_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nand _47942_ (_24779_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47943_ (_24780_, _24779_, _24778_);
  and _47944_ (_24781_, _24780_, _24777_);
  and _47945_ (_24782_, _24781_, _24774_);
  nand _47946_ (_24783_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _47947_ (_24784_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47948_ (_24785_, _24784_, _24783_);
  nand _47949_ (_24786_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nand _47950_ (_24787_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _47951_ (_24788_, _24787_, _24786_);
  and _47952_ (_24789_, _24788_, _24785_);
  nand _47953_ (_24790_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  nand _47954_ (_24791_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _47955_ (_24792_, _24791_, _24790_);
  nand _47956_ (_24793_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _47957_ (_24794_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _47958_ (_24795_, _24794_, _24793_);
  and _47959_ (_24796_, _24795_, _24792_);
  and _47960_ (_24797_, _24796_, _24789_);
  and _47961_ (_24798_, _24797_, _24782_);
  nand _47962_ (_24799_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _47963_ (_24800_, _24743_, _02296_);
  and _47964_ (_24801_, _24800_, _24799_);
  nand _47965_ (_24802_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand _47966_ (_24803_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _47967_ (_24804_, _24803_, _24802_);
  and _47968_ (_24805_, _24804_, _24801_);
  nand _47969_ (_24806_, _24685_, _24478_);
  nand _47970_ (_24807_, _24687_, _24237_);
  and _47971_ (_24808_, _24807_, _24806_);
  nand _47972_ (_24809_, _24682_, _24267_);
  nand _47973_ (_24810_, _24680_, _24392_);
  and _47974_ (_24811_, _24810_, _24809_);
  and _47975_ (_24812_, _24811_, _24808_);
  and _47976_ (_24813_, _24812_, _24805_);
  nand _47977_ (_24814_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand _47978_ (_24815_, _24573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _47979_ (_24816_, _24815_, _24814_);
  and _47980_ (_24817_, _24816_, _24813_);
  and _47981_ (_24818_, _24817_, _24798_);
  nor _47982_ (_24819_, _24564_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or _47983_ (_24820_, _24819_, _24577_);
  nor _47984_ (_24821_, _24820_, _24818_);
  or _47985_ (_24822_, _24821_, _24582_);
  or _47986_ (_24823_, _24822_, _24767_);
  or _47987_ (_24824_, _24700_, _01397_);
  and _47988_ (_24825_, _24824_, _25365_);
  and _47989_ (_06519_, _24825_, _24823_);
  and _47990_ (_24826_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _47991_ (_24827_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _47992_ (_24828_, _24827_, _24826_);
  and _47993_ (_24829_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _47994_ (_24830_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _47995_ (_24831_, _24830_, _24829_);
  or _47996_ (_24832_, _24831_, _24828_);
  and _47997_ (_24833_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _47998_ (_24834_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _47999_ (_24835_, _24834_, _24833_);
  and _48000_ (_24836_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _48001_ (_24837_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _48002_ (_24838_, _24837_, _24836_);
  or _48003_ (_24839_, _24838_, _24835_);
  or _48004_ (_24840_, _24839_, _24832_);
  and _48005_ (_24841_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _48006_ (_24842_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or _48007_ (_24843_, _24842_, _24841_);
  and _48008_ (_24844_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _48009_ (_24845_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _48010_ (_24846_, _24845_, _24844_);
  or _48011_ (_24847_, _24846_, _24843_);
  and _48012_ (_24848_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _48013_ (_24849_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _48014_ (_24850_, _24849_, _24848_);
  and _48015_ (_24851_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _48016_ (_24852_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _48017_ (_24853_, _24852_, _24851_);
  or _48018_ (_24854_, _24853_, _24850_);
  or _48019_ (_24855_, _24854_, _24847_);
  or _48020_ (_24856_, _24855_, _24840_);
  and _48021_ (_24857_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _48022_ (_24858_, _24630_, _05914_);
  or _48023_ (_24859_, _24858_, _24857_);
  and _48024_ (_24860_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _48025_ (_24861_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or _48026_ (_24862_, _24861_, _24860_);
  or _48027_ (_24863_, _24862_, _24859_);
  and _48028_ (_24864_, _24685_, _24491_);
  and _48029_ (_24865_, _24687_, _24224_);
  or _48030_ (_24866_, _24865_, _24864_);
  and _48031_ (_24867_, _24682_, _24276_);
  and _48032_ (_24868_, _24680_, _24401_);
  or _48033_ (_24869_, _24868_, _24867_);
  or _48034_ (_24870_, _24869_, _24866_);
  or _48035_ (_24871_, _24870_, _24863_);
  and _48036_ (_24872_, _24573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _48037_ (_24873_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _48038_ (_24874_, _24873_, _24872_);
  or _48039_ (_24875_, _24874_, _24871_);
  or _48040_ (_24876_, _24875_, _24856_);
  and _48041_ (_24877_, _24876_, _24579_);
  and _48042_ (_24878_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or _48043_ (_24879_, _24878_, _24877_);
  or _48044_ (_24880_, _24879_, _24582_);
  or _48045_ (_24881_, _24700_, _01457_);
  and _48046_ (_24882_, _24881_, _25365_);
  and _48047_ (_06520_, _24882_, _24880_);
  and _48048_ (_24883_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _48049_ (_24884_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _48050_ (_24885_, _24884_, _24883_);
  and _48051_ (_24886_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _48052_ (_24887_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _48053_ (_24888_, _24887_, _24886_);
  or _48054_ (_24889_, _24888_, _24885_);
  and _48055_ (_24890_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _48056_ (_24891_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _48057_ (_24892_, _24891_, _24890_);
  and _48058_ (_24893_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _48059_ (_24894_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _48060_ (_24895_, _24894_, _24893_);
  or _48061_ (_24896_, _24895_, _24892_);
  or _48062_ (_24897_, _24896_, _24889_);
  and _48063_ (_24898_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _48064_ (_24899_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _48065_ (_24900_, _24899_, _24898_);
  and _48066_ (_24901_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _48067_ (_24902_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _48068_ (_24903_, _24902_, _24901_);
  or _48069_ (_24904_, _24903_, _24900_);
  and _48070_ (_24905_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _48071_ (_24906_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _48072_ (_24907_, _24906_, _24905_);
  and _48073_ (_24908_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _48074_ (_24909_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _48075_ (_24910_, _24909_, _24908_);
  or _48076_ (_24911_, _24910_, _24907_);
  or _48077_ (_24912_, _24911_, _24904_);
  or _48078_ (_24913_, _24912_, _24897_);
  nor _48079_ (_24914_, _24743_, _02308_);
  and _48080_ (_24915_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _48081_ (_24916_, _24915_, _24914_);
  and _48082_ (_24917_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _48083_ (_24918_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or _48084_ (_24919_, _24918_, _24917_);
  or _48085_ (_24920_, _24919_, _24916_);
  and _48086_ (_24921_, _24685_, _24487_);
  and _48087_ (_24922_, _24687_, _24233_);
  or _48088_ (_24923_, _24922_, _24921_);
  and _48089_ (_24924_, _24682_, _24280_);
  and _48090_ (_24925_, _24680_, _24396_);
  or _48091_ (_24926_, _24925_, _24924_);
  or _48092_ (_24927_, _24926_, _24923_);
  or _48093_ (_24928_, _24927_, _24920_);
  and _48094_ (_24929_, _24573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _48095_ (_24930_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _48096_ (_24931_, _24930_, _24929_);
  or _48097_ (_24932_, _24931_, _24928_);
  or _48098_ (_24933_, _24932_, _24913_);
  and _48099_ (_24934_, _24933_, _24579_);
  and _48100_ (_24935_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or _48101_ (_24936_, _24935_, _24934_);
  or _48102_ (_24937_, _24936_, _24582_);
  or _48103_ (_24938_, _24700_, _01522_);
  and _48104_ (_24939_, _24938_, _25365_);
  and _48105_ (_06521_, _24939_, _24937_);
  and _48106_ (_24940_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _48107_ (_24941_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _48108_ (_24942_, _24941_, _24940_);
  and _48109_ (_24943_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _48110_ (_24944_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _48111_ (_24945_, _24944_, _24943_);
  or _48112_ (_24946_, _24945_, _24942_);
  and _48113_ (_24947_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _48114_ (_24948_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or _48115_ (_24949_, _24948_, _24947_);
  and _48116_ (_24950_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _48117_ (_24951_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _48118_ (_24952_, _24951_, _24950_);
  or _48119_ (_24953_, _24952_, _24949_);
  or _48120_ (_24954_, _24953_, _24946_);
  and _48121_ (_24955_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _48122_ (_24956_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _48123_ (_24957_, _24956_, _24955_);
  and _48124_ (_24958_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _48125_ (_24959_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _48126_ (_24960_, _24959_, _24958_);
  or _48127_ (_24961_, _24960_, _24957_);
  and _48128_ (_24962_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _48129_ (_24963_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _48130_ (_24964_, _24963_, _24962_);
  and _48131_ (_24965_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _48132_ (_24966_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _48133_ (_24967_, _24966_, _24965_);
  or _48134_ (_24968_, _24967_, _24964_);
  or _48135_ (_24969_, _24968_, _24961_);
  or _48136_ (_24970_, _24969_, _24954_);
  and _48137_ (_24971_, _24573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _48138_ (_24972_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _48139_ (_24973_, _24972_, _24971_);
  and _48140_ (_24974_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _48141_ (_24975_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _48142_ (_24976_, _24975_, _24974_);
  nor _48143_ (_24977_, _24743_, _02314_);
  and _48144_ (_24978_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _48145_ (_24979_, _24978_, _24977_);
  or _48146_ (_24980_, _24979_, _24976_);
  and _48147_ (_24981_, _24685_, _24461_);
  and _48148_ (_24982_, _24687_, _24248_);
  or _48149_ (_24983_, _24982_, _24981_);
  and _48150_ (_24984_, _24680_, _24385_);
  and _48151_ (_24985_, _24682_, _24291_);
  or _48152_ (_24986_, _24985_, _24984_);
  or _48153_ (_24987_, _24986_, _24983_);
  or _48154_ (_24988_, _24987_, _24980_);
  or _48155_ (_24989_, _24988_, _24973_);
  or _48156_ (_24990_, _24989_, _24970_);
  and _48157_ (_24991_, _24990_, _24579_);
  and _48158_ (_24992_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or _48159_ (_24993_, _24992_, _24991_);
  or _48160_ (_24994_, _24993_, _24582_);
  or _48161_ (_24995_, _24700_, _01589_);
  and _48162_ (_24996_, _24995_, _25365_);
  and _48163_ (_06522_, _24996_, _24994_);
  and _48164_ (_24997_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _48165_ (_24998_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _48166_ (_24999_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _48167_ (_25000_, _24999_, _24998_);
  and _48168_ (_25001_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48169_ (_25002_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _48170_ (_25003_, _25002_, _25001_);
  or _48171_ (_25004_, _25003_, _25000_);
  and _48172_ (_25005_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _48173_ (_25006_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or _48174_ (_25007_, _25006_, _25005_);
  and _48175_ (_25008_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _48176_ (_25009_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _48177_ (_25010_, _25009_, _25008_);
  or _48178_ (_25011_, _25010_, _25007_);
  or _48179_ (_25012_, _25011_, _25004_);
  and _48180_ (_25013_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _48181_ (_25014_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _48182_ (_25015_, _25014_, _25013_);
  and _48183_ (_25016_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _48184_ (_25017_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _48185_ (_25018_, _25017_, _25016_);
  or _48186_ (_25019_, _25018_, _25015_);
  and _48187_ (_25020_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _48188_ (_25021_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _48189_ (_25022_, _25021_, _25020_);
  and _48190_ (_25023_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _48191_ (_25024_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _48192_ (_25025_, _25024_, _25023_);
  or _48193_ (_25026_, _25025_, _25022_);
  or _48194_ (_25027_, _25026_, _25019_);
  or _48195_ (_25028_, _25027_, _25012_);
  and _48196_ (_25029_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor _48197_ (_25030_, _24743_, _02320_);
  or _48198_ (_25031_, _25030_, _25029_);
  and _48199_ (_25032_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _48200_ (_25033_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _48201_ (_25034_, _25033_, _25032_);
  or _48202_ (_25035_, _25034_, _25031_);
  and _48203_ (_25036_, _24685_, _24456_);
  and _48204_ (_25037_, _24687_, _24257_);
  or _48205_ (_25038_, _25037_, _25036_);
  and _48206_ (_25039_, _24680_, _24372_);
  and _48207_ (_25040_, _24682_, _24287_);
  or _48208_ (_25041_, _25040_, _25039_);
  or _48209_ (_25042_, _25041_, _25038_);
  or _48210_ (_25043_, _25042_, _25035_);
  and _48211_ (_25044_, _24573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _48212_ (_25045_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _48213_ (_25046_, _25045_, _25044_);
  or _48214_ (_25047_, _25046_, _25043_);
  nor _48215_ (_25048_, _25047_, _25028_);
  nor _48216_ (_25049_, _24564_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or _48217_ (_25050_, _25049_, _24577_);
  nor _48218_ (_25051_, _25050_, _25048_);
  or _48219_ (_25052_, _25051_, _24582_);
  or _48220_ (_25053_, _25052_, _24997_);
  or _48221_ (_25054_, _24700_, _01673_);
  and _48222_ (_25055_, _25054_, _25365_);
  and _48223_ (_06523_, _25055_, _25053_);
  and _48224_ (_25056_, _24638_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _48225_ (_25057_, _24642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _48226_ (_25058_, _24640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _48227_ (_25059_, _25058_, _25057_);
  nand _48228_ (_25060_, _24592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand _48229_ (_25061_, _24589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _48230_ (_25062_, _25061_, _25060_);
  and _48231_ (_25063_, _25062_, _25059_);
  nand _48232_ (_25064_, _24598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand _48233_ (_25065_, _24596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _48234_ (_25066_, _25065_, _25064_);
  nand _48235_ (_25067_, _24600_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  nand _48236_ (_25068_, _24604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _48237_ (_25069_, _25068_, _25067_);
  and _48238_ (_25070_, _25069_, _25066_);
  and _48239_ (_25071_, _25070_, _25063_);
  nand _48240_ (_25072_, _24609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nand _48241_ (_25073_, _24610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _48242_ (_25074_, _25073_, _25072_);
  nand _48243_ (_25075_, _24613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _48244_ (_25076_, _24612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _48245_ (_25077_, _25076_, _25075_);
  and _48246_ (_25078_, _25077_, _25074_);
  nand _48247_ (_25079_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _48248_ (_25080_, _24621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _48249_ (_25081_, _25080_, _25079_);
  nand _48250_ (_25082_, _24617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _48251_ (_25083_, _24618_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _48252_ (_25084_, _25083_, _25082_);
  and _48253_ (_25085_, _25084_, _25081_);
  and _48254_ (_25086_, _25085_, _25078_);
  and _48255_ (_25087_, _25086_, _25071_);
  or _48256_ (_25088_, _24743_, _02326_);
  nand _48257_ (_25089_, _24631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _48258_ (_25090_, _25089_, _25088_);
  nand _48259_ (_25091_, _24581_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand _48260_ (_25092_, _24566_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _48261_ (_25093_, _25092_, _25091_);
  and _48262_ (_25094_, _25093_, _25090_);
  nand _48263_ (_25095_, _24685_, _24469_);
  nand _48264_ (_25096_, _24687_, _24244_);
  and _48265_ (_25097_, _25096_, _25095_);
  nand _48266_ (_25098_, _24680_, _24381_);
  nand _48267_ (_25099_, _24682_, _24296_);
  and _48268_ (_25100_, _25099_, _25098_);
  and _48269_ (_25101_, _25100_, _25097_);
  and _48270_ (_25102_, _25101_, _25094_);
  nand _48271_ (_25103_, _24573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _48272_ (_25104_, _24557_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _48273_ (_25105_, _25104_, _25103_);
  and _48274_ (_25106_, _25105_, _25102_);
  and _48275_ (_25107_, _25106_, _25087_);
  nor _48276_ (_25108_, _24564_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or _48277_ (_25109_, _25108_, _24577_);
  nor _48278_ (_25110_, _25109_, _25107_);
  or _48279_ (_25111_, _25110_, _24582_);
  or _48280_ (_25112_, _25111_, _25056_);
  or _48281_ (_25113_, _24700_, _01737_);
  and _48282_ (_25114_, _25113_, _25365_);
  and _48283_ (_06524_, _25114_, _25112_);
  and _48284_ (_06533_, _06019_, _25365_);
  and _48285_ (_06534_, _09510_, _25365_);
  nor _48286_ (_06536_, _05918_, rst);
  and _48287_ (_06538_, _09334_, _25365_);
  and _48288_ (_06539_, _09453_, _25365_);
  and _48289_ (_06540_, _09463_, _25365_);
  and _48290_ (_06541_, _09472_, _25365_);
  and _48291_ (_06542_, _09482_, _25365_);
  and _48292_ (_06543_, _09492_, _25365_);
  and _48293_ (_06544_, _09502_, _25365_);
  nor _48294_ (_06545_, _05720_, rst);
  nor _48295_ (_06546_, _05994_, rst);
  and _48296_ (_06584_, \uc8051golden_1.B [7], _25365_);
  and _48297_ (_06585_, \uc8051golden_1.ACC [7], _25365_);
  and _48298_ (_06586_, \uc8051golden_1.PCON [7], _25365_);
  and _48299_ (_06587_, \uc8051golden_1.TMOD [7], _25365_);
  and _48300_ (_06588_, \uc8051golden_1.DPL [7], _25365_);
  and _48301_ (_06590_, \uc8051golden_1.DPH [7], _25365_);
  and _48302_ (_06591_, \uc8051golden_1.TL1 [7], _25365_);
  and _48303_ (_06592_, \uc8051golden_1.TL0 [7], _25365_);
  and _48304_ (_06593_, \uc8051golden_1.TCON [7], _25365_);
  and _48305_ (_06594_, \uc8051golden_1.TH1 [7], _25365_);
  and _48306_ (_06595_, \uc8051golden_1.TH0 [7], _25365_);
  not _48307_ (_25115_, \uc8051golden_1.PC [15]);
  and _48308_ (_25116_, \uc8051golden_1.PC [1], \uc8051golden_1.PC [0]);
  and _48309_ (_25117_, _25116_, \uc8051golden_1.PC [2]);
  and _48310_ (_25118_, _25117_, \uc8051golden_1.PC [3]);
  and _48311_ (_25119_, _25118_, \uc8051golden_1.PC [4]);
  and _48312_ (_25120_, _25119_, \uc8051golden_1.PC [5]);
  and _48313_ (_25121_, _25120_, \uc8051golden_1.PC [6]);
  and _48314_ (_25122_, _25121_, \uc8051golden_1.PC [7]);
  and _48315_ (_25123_, _25122_, \uc8051golden_1.PC [8]);
  and _48316_ (_25124_, _25123_, \uc8051golden_1.PC [9]);
  and _48317_ (_25125_, _25124_, \uc8051golden_1.PC [10]);
  and _48318_ (_25126_, _25125_, \uc8051golden_1.PC [11]);
  and _48319_ (_25127_, _25126_, \uc8051golden_1.PC [12]);
  and _48320_ (_25128_, _25127_, \uc8051golden_1.PC [13]);
  nand _48321_ (_25129_, _25128_, \uc8051golden_1.PC [14]);
  nand _48322_ (_25130_, _25129_, _25115_);
  or _48323_ (_25131_, _25129_, _25115_);
  and _48324_ (_25132_, _25131_, _25130_);
  or _48325_ (_25133_, _25132_, _22350_);
  or _48326_ (_25134_, _22345_, \uc8051golden_1.PC [15]);
  and _48327_ (_25135_, _25134_, _25365_);
  and _48328_ (_06596_, _25135_, _25133_);
  and _48329_ (_06597_, \uc8051golden_1.P2 [7], _25365_);
  and _48330_ (_06598_, \uc8051golden_1.P3 [7], _25365_);
  and _48331_ (_06599_, \uc8051golden_1.P0 [7], _25365_);
  and _48332_ (_06600_, \uc8051golden_1.P1 [7], _25365_);
  and _48333_ (_06601_, \uc8051golden_1.IP [7], _25365_);
  and _48334_ (_06602_, \uc8051golden_1.IE [7], _25365_);
  and _48335_ (_06603_, \uc8051golden_1.SCON [7], _25365_);
  and _48336_ (_06604_, \uc8051golden_1.SP [7], _25365_);
  and _48337_ (_06605_, \uc8051golden_1.SBUF [7], _25365_);
  and _48338_ (_06606_, \uc8051golden_1.PSW [7], _25365_);
  and _48339_ (_09277_, \uc8051golden_1.B [0], _25365_);
  and _48340_ (_09278_, \uc8051golden_1.B [1], _25365_);
  and _48341_ (_09279_, \uc8051golden_1.B [2], _25365_);
  and _48342_ (_09280_, \uc8051golden_1.B [3], _25365_);
  and _48343_ (_09281_, \uc8051golden_1.B [4], _25365_);
  and _48344_ (_09282_, \uc8051golden_1.B [5], _25365_);
  and _48345_ (_09283_, \uc8051golden_1.B [6], _25365_);
  and _48346_ (_09284_, \uc8051golden_1.ACC [0], _25365_);
  and _48347_ (_09285_, \uc8051golden_1.ACC [1], _25365_);
  and _48348_ (_09286_, \uc8051golden_1.ACC [2], _25365_);
  and _48349_ (_09287_, \uc8051golden_1.ACC [3], _25365_);
  and _48350_ (_09288_, \uc8051golden_1.ACC [4], _25365_);
  and _48351_ (_09289_, \uc8051golden_1.ACC [5], _25365_);
  and _48352_ (_09290_, \uc8051golden_1.ACC [6], _25365_);
  and _48353_ (_09291_, \uc8051golden_1.PCON [0], _25365_);
  and _48354_ (_09292_, \uc8051golden_1.PCON [1], _25365_);
  and _48355_ (_09293_, \uc8051golden_1.PCON [2], _25365_);
  and _48356_ (_09294_, \uc8051golden_1.PCON [3], _25365_);
  and _48357_ (_09295_, \uc8051golden_1.PCON [4], _25365_);
  and _48358_ (_09296_, \uc8051golden_1.PCON [5], _25365_);
  and _48359_ (_09297_, \uc8051golden_1.PCON [6], _25365_);
  and _48360_ (_09298_, \uc8051golden_1.TMOD [0], _25365_);
  and _48361_ (_09299_, \uc8051golden_1.TMOD [1], _25365_);
  and _48362_ (_09300_, \uc8051golden_1.TMOD [2], _25365_);
  and _48363_ (_09301_, \uc8051golden_1.TMOD [3], _25365_);
  and _48364_ (_09302_, \uc8051golden_1.TMOD [4], _25365_);
  and _48365_ (_09303_, \uc8051golden_1.TMOD [5], _25365_);
  and _48366_ (_09304_, \uc8051golden_1.TMOD [6], _25365_);
  and _48367_ (_09305_, \uc8051golden_1.DPL [0], _25365_);
  and _48368_ (_09306_, \uc8051golden_1.DPL [1], _25365_);
  and _48369_ (_09307_, \uc8051golden_1.DPL [2], _25365_);
  and _48370_ (_09309_, \uc8051golden_1.DPL [3], _25365_);
  and _48371_ (_09310_, \uc8051golden_1.DPL [4], _25365_);
  and _48372_ (_09311_, \uc8051golden_1.DPL [5], _25365_);
  and _48373_ (_09312_, \uc8051golden_1.DPL [6], _25365_);
  and _48374_ (_09313_, \uc8051golden_1.DPH [0], _25365_);
  and _48375_ (_09314_, \uc8051golden_1.DPH [1], _25365_);
  and _48376_ (_09315_, \uc8051golden_1.DPH [2], _25365_);
  and _48377_ (_09316_, \uc8051golden_1.DPH [3], _25365_);
  and _48378_ (_09317_, \uc8051golden_1.DPH [4], _25365_);
  and _48379_ (_09318_, \uc8051golden_1.DPH [5], _25365_);
  and _48380_ (_09319_, \uc8051golden_1.DPH [6], _25365_);
  and _48381_ (_09320_, \uc8051golden_1.TL1 [0], _25365_);
  and _48382_ (_09321_, \uc8051golden_1.TL1 [1], _25365_);
  and _48383_ (_09322_, \uc8051golden_1.TL1 [2], _25365_);
  and _48384_ (_09323_, \uc8051golden_1.TL1 [3], _25365_);
  and _48385_ (_09324_, \uc8051golden_1.TL1 [4], _25365_);
  and _48386_ (_09325_, \uc8051golden_1.TL1 [5], _25365_);
  and _48387_ (_09326_, \uc8051golden_1.TL1 [6], _25365_);
  and _48388_ (_09327_, \uc8051golden_1.TL0 [0], _25365_);
  and _48389_ (_09328_, \uc8051golden_1.TL0 [1], _25365_);
  and _48390_ (_09329_, \uc8051golden_1.TL0 [2], _25365_);
  and _48391_ (_09330_, \uc8051golden_1.TL0 [3], _25365_);
  and _48392_ (_09331_, \uc8051golden_1.TL0 [4], _25365_);
  and _48393_ (_09332_, \uc8051golden_1.TL0 [5], _25365_);
  and _48394_ (_09333_, \uc8051golden_1.TL0 [6], _25365_);
  and _48395_ (_09335_, \uc8051golden_1.TCON [0], _25365_);
  and _48396_ (_09336_, \uc8051golden_1.TCON [1], _25365_);
  and _48397_ (_09337_, \uc8051golden_1.TCON [2], _25365_);
  and _48398_ (_09338_, \uc8051golden_1.TCON [3], _25365_);
  and _48399_ (_09339_, \uc8051golden_1.TCON [4], _25365_);
  and _48400_ (_09340_, \uc8051golden_1.TCON [5], _25365_);
  and _48401_ (_09341_, \uc8051golden_1.TCON [6], _25365_);
  and _48402_ (_09342_, \uc8051golden_1.TH1 [0], _25365_);
  and _48403_ (_09343_, \uc8051golden_1.TH1 [1], _25365_);
  and _48404_ (_09344_, \uc8051golden_1.TH1 [2], _25365_);
  and _48405_ (_09345_, \uc8051golden_1.TH1 [3], _25365_);
  and _48406_ (_09346_, \uc8051golden_1.TH1 [4], _25365_);
  and _48407_ (_09347_, \uc8051golden_1.TH1 [5], _25365_);
  and _48408_ (_09348_, \uc8051golden_1.TH1 [6], _25365_);
  and _48409_ (_09349_, \uc8051golden_1.TH0 [0], _25365_);
  and _48410_ (_09350_, \uc8051golden_1.TH0 [1], _25365_);
  and _48411_ (_09351_, \uc8051golden_1.TH0 [2], _25365_);
  and _48412_ (_09352_, \uc8051golden_1.TH0 [3], _25365_);
  and _48413_ (_09353_, \uc8051golden_1.TH0 [4], _25365_);
  and _48414_ (_09354_, \uc8051golden_1.TH0 [5], _25365_);
  and _48415_ (_09355_, \uc8051golden_1.TH0 [6], _25365_);
  nand _48416_ (_25136_, _22345_, \uc8051golden_1.PC [0]);
  or _48417_ (_25137_, _22345_, \uc8051golden_1.PC [0]);
  and _48418_ (_25138_, _25137_, _25136_);
  and _48419_ (_09357_, _25138_, _25365_);
  or _48420_ (_25139_, _22345_, \uc8051golden_1.PC [1]);
  nor _48421_ (_25140_, \uc8051golden_1.PC [1], \uc8051golden_1.PC [0]);
  nor _48422_ (_25141_, _25140_, _25116_);
  or _48423_ (_25142_, _25141_, _22350_);
  and _48424_ (_25143_, _25142_, _25365_);
  and _48425_ (_09358_, _25143_, _25139_);
  or _48426_ (_25144_, _22345_, \uc8051golden_1.PC [2]);
  nor _48427_ (_25145_, _25116_, \uc8051golden_1.PC [2]);
  nor _48428_ (_25146_, _25145_, _25117_);
  or _48429_ (_25147_, _25146_, _22350_);
  and _48430_ (_25148_, _25147_, _25365_);
  and _48431_ (_09359_, _25148_, _25144_);
  nor _48432_ (_25149_, _25117_, \uc8051golden_1.PC [3]);
  nor _48433_ (_25150_, _25149_, _25118_);
  and _48434_ (_25151_, _25150_, _22345_);
  and _48435_ (_25152_, _22350_, \uc8051golden_1.PC [3]);
  or _48436_ (_25153_, _25152_, _25151_);
  and _48437_ (_09360_, _25153_, _25365_);
  nor _48438_ (_25154_, _25118_, \uc8051golden_1.PC [4]);
  nor _48439_ (_25155_, _25154_, _25119_);
  or _48440_ (_25156_, _25155_, _22350_);
  or _48441_ (_25157_, _22345_, \uc8051golden_1.PC [4]);
  and _48442_ (_25158_, _25157_, _25365_);
  and _48443_ (_09361_, _25158_, _25156_);
  nor _48444_ (_25159_, _25119_, \uc8051golden_1.PC [5]);
  nor _48445_ (_25160_, _25159_, _25120_);
  or _48446_ (_25161_, _25160_, _22350_);
  or _48447_ (_25162_, _22345_, \uc8051golden_1.PC [5]);
  and _48448_ (_25163_, _25162_, _25365_);
  and _48449_ (_09362_, _25163_, _25161_);
  nor _48450_ (_25164_, _25120_, \uc8051golden_1.PC [6]);
  nor _48451_ (_25165_, _25164_, _25121_);
  or _48452_ (_25166_, _25165_, _22350_);
  or _48453_ (_25167_, _22345_, \uc8051golden_1.PC [6]);
  and _48454_ (_25168_, _25167_, _25365_);
  and _48455_ (_09363_, _25168_, _25166_);
  nor _48456_ (_25169_, _25121_, \uc8051golden_1.PC [7]);
  nor _48457_ (_25170_, _25169_, _25122_);
  or _48458_ (_25171_, _25170_, _22350_);
  or _48459_ (_25172_, _22345_, \uc8051golden_1.PC [7]);
  and _48460_ (_25173_, _25172_, _25365_);
  and _48461_ (_09364_, _25173_, _25171_);
  nor _48462_ (_25174_, _25122_, \uc8051golden_1.PC [8]);
  nor _48463_ (_25175_, _25174_, _25123_);
  or _48464_ (_25176_, _25175_, _22350_);
  or _48465_ (_25177_, _22345_, \uc8051golden_1.PC [8]);
  and _48466_ (_25178_, _25177_, _25365_);
  and _48467_ (_09365_, _25178_, _25176_);
  nor _48468_ (_25179_, _25123_, \uc8051golden_1.PC [9]);
  nor _48469_ (_25180_, _25179_, _25124_);
  or _48470_ (_25181_, _25180_, _22350_);
  or _48471_ (_25182_, _22345_, \uc8051golden_1.PC [9]);
  and _48472_ (_25183_, _25182_, _25365_);
  and _48473_ (_09366_, _25183_, _25181_);
  nor _48474_ (_25184_, _25124_, \uc8051golden_1.PC [10]);
  nor _48475_ (_25185_, _25184_, _25125_);
  or _48476_ (_25186_, _25185_, _22350_);
  or _48477_ (_25187_, _22345_, \uc8051golden_1.PC [10]);
  and _48478_ (_25188_, _25187_, _25365_);
  and _48479_ (_09367_, _25188_, _25186_);
  nor _48480_ (_25189_, _25125_, \uc8051golden_1.PC [11]);
  nor _48481_ (_25190_, _25189_, _25126_);
  or _48482_ (_25191_, _25190_, _22350_);
  or _48483_ (_25192_, _22345_, \uc8051golden_1.PC [11]);
  and _48484_ (_25193_, _25192_, _25365_);
  and _48485_ (_09368_, _25193_, _25191_);
  nor _48486_ (_25194_, _25126_, \uc8051golden_1.PC [12]);
  nor _48487_ (_25195_, _25194_, _25127_);
  or _48488_ (_25196_, _25195_, _22350_);
  or _48489_ (_25197_, _22345_, \uc8051golden_1.PC [12]);
  and _48490_ (_25198_, _25197_, _25365_);
  and _48491_ (_09369_, _25198_, _25196_);
  nor _48492_ (_25199_, _25127_, \uc8051golden_1.PC [13]);
  nor _48493_ (_25200_, _25199_, _25128_);
  or _48494_ (_25201_, _25200_, _22350_);
  or _48495_ (_25202_, _22345_, \uc8051golden_1.PC [13]);
  and _48496_ (_25203_, _25202_, _25365_);
  and _48497_ (_09370_, _25203_, _25201_);
  or _48498_ (_25204_, _25128_, \uc8051golden_1.PC [14]);
  and _48499_ (_25205_, _25204_, _25129_);
  or _48500_ (_25206_, _25205_, _22350_);
  or _48501_ (_25207_, _22345_, \uc8051golden_1.PC [14]);
  and _48502_ (_25208_, _25207_, _25365_);
  and _48503_ (_09371_, _25208_, _25206_);
  and _48504_ (_09372_, \uc8051golden_1.P2 [0], _25365_);
  and _48505_ (_09373_, \uc8051golden_1.P2 [1], _25365_);
  and _48506_ (_09374_, \uc8051golden_1.P2 [2], _25365_);
  and _48507_ (_09375_, \uc8051golden_1.P2 [3], _25365_);
  and _48508_ (_09376_, \uc8051golden_1.P2 [4], _25365_);
  and _48509_ (_09377_, \uc8051golden_1.P2 [5], _25365_);
  and _48510_ (_09378_, \uc8051golden_1.P2 [6], _25365_);
  and _48511_ (_09379_, \uc8051golden_1.P3 [0], _25365_);
  and _48512_ (_09380_, \uc8051golden_1.P3 [1], _25365_);
  and _48513_ (_09381_, \uc8051golden_1.P3 [2], _25365_);
  and _48514_ (_09382_, \uc8051golden_1.P3 [3], _25365_);
  and _48515_ (_09383_, \uc8051golden_1.P3 [4], _25365_);
  and _48516_ (_09384_, \uc8051golden_1.P3 [5], _25365_);
  and _48517_ (_09385_, \uc8051golden_1.P3 [6], _25365_);
  and _48518_ (_09386_, \uc8051golden_1.P0 [0], _25365_);
  and _48519_ (_09387_, \uc8051golden_1.P0 [1], _25365_);
  and _48520_ (_09388_, \uc8051golden_1.P0 [2], _25365_);
  and _48521_ (_09389_, \uc8051golden_1.P0 [3], _25365_);
  and _48522_ (_09390_, \uc8051golden_1.P0 [4], _25365_);
  and _48523_ (_09391_, \uc8051golden_1.P0 [5], _25365_);
  and _48524_ (_09392_, \uc8051golden_1.P0 [6], _25365_);
  and _48525_ (_09393_, \uc8051golden_1.P1 [0], _25365_);
  and _48526_ (_09394_, \uc8051golden_1.P1 [1], _25365_);
  and _48527_ (_09395_, \uc8051golden_1.P1 [2], _25365_);
  and _48528_ (_09396_, \uc8051golden_1.P1 [3], _25365_);
  and _48529_ (_09397_, \uc8051golden_1.P1 [4], _25365_);
  and _48530_ (_09398_, \uc8051golden_1.P1 [5], _25365_);
  and _48531_ (_09399_, \uc8051golden_1.P1 [6], _25365_);
  and _48532_ (_09400_, \uc8051golden_1.IP [0], _25365_);
  and _48533_ (_09401_, \uc8051golden_1.IP [1], _25365_);
  and _48534_ (_09402_, \uc8051golden_1.IP [2], _25365_);
  and _48535_ (_09403_, \uc8051golden_1.IP [3], _25365_);
  and _48536_ (_09404_, \uc8051golden_1.IP [4], _25365_);
  and _48537_ (_09405_, \uc8051golden_1.IP [5], _25365_);
  and _48538_ (_09406_, \uc8051golden_1.IP [6], _25365_);
  and _48539_ (_09407_, \uc8051golden_1.IE [0], _25365_);
  and _48540_ (_09408_, \uc8051golden_1.IE [1], _25365_);
  and _48541_ (_09409_, \uc8051golden_1.IE [2], _25365_);
  and _48542_ (_09410_, \uc8051golden_1.IE [3], _25365_);
  and _48543_ (_09411_, \uc8051golden_1.IE [4], _25365_);
  and _48544_ (_09412_, \uc8051golden_1.IE [5], _25365_);
  and _48545_ (_09413_, \uc8051golden_1.IE [6], _25365_);
  and _48546_ (_09414_, \uc8051golden_1.SCON [0], _25365_);
  and _48547_ (_09415_, \uc8051golden_1.SCON [1], _25365_);
  and _48548_ (_09417_, \uc8051golden_1.SCON [2], _25365_);
  and _48549_ (_09418_, \uc8051golden_1.SCON [3], _25365_);
  and _48550_ (_09419_, \uc8051golden_1.SCON [4], _25365_);
  and _48551_ (_09420_, \uc8051golden_1.SCON [5], _25365_);
  and _48552_ (_09421_, \uc8051golden_1.SCON [6], _25365_);
  and _48553_ (_09422_, \uc8051golden_1.SP [0], _25365_);
  and _48554_ (_09423_, \uc8051golden_1.SP [1], _25365_);
  and _48555_ (_09424_, \uc8051golden_1.SP [2], _25365_);
  and _48556_ (_09425_, \uc8051golden_1.SP [3], _25365_);
  and _48557_ (_09426_, \uc8051golden_1.SP [4], _25365_);
  and _48558_ (_09427_, \uc8051golden_1.SP [5], _25365_);
  and _48559_ (_09428_, \uc8051golden_1.SP [6], _25365_);
  and _48560_ (_09429_, \uc8051golden_1.SBUF [0], _25365_);
  and _48561_ (_09430_, \uc8051golden_1.SBUF [1], _25365_);
  and _48562_ (_09431_, \uc8051golden_1.SBUF [2], _25365_);
  and _48563_ (_09432_, \uc8051golden_1.SBUF [3], _25365_);
  and _48564_ (_09433_, \uc8051golden_1.SBUF [4], _25365_);
  and _48565_ (_09434_, \uc8051golden_1.SBUF [5], _25365_);
  and _48566_ (_09435_, \uc8051golden_1.SBUF [6], _25365_);
  and _48567_ (_09436_, \uc8051golden_1.PSW [0], _25365_);
  and _48568_ (_09437_, \uc8051golden_1.PSW [1], _25365_);
  and _48569_ (_09438_, \uc8051golden_1.PSW [2], _25365_);
  and _48570_ (_09439_, \uc8051golden_1.PSW [3], _25365_);
  and _48571_ (_09440_, \uc8051golden_1.PSW [4], _25365_);
  and _48572_ (_09441_, \uc8051golden_1.PSW [5], _25365_);
  and _48573_ (_09442_, \uc8051golden_1.PSW [6], _25365_);
  nor _48574_ (_25209_, _25132_, _02402_);
  and _48575_ (_25210_, _25132_, _02402_);
  or _48576_ (_25211_, _25210_, _25209_);
  nor _48577_ (_25212_, _25205_, _02397_);
  and _48578_ (_25213_, _25205_, _02397_);
  or _48579_ (_25214_, _25213_, _25212_);
  nor _48580_ (_25215_, _25200_, _02366_);
  and _48581_ (_25216_, _25200_, _02366_);
  or _48582_ (_25217_, _25216_, _25215_);
  nor _48583_ (_25218_, _25195_, _02391_);
  and _48584_ (_25219_, _25195_, _02391_);
  or _48585_ (_25220_, _25219_, _25218_);
  nor _48586_ (_25221_, _25190_, _02370_);
  and _48587_ (_25222_, _25190_, _02370_);
  or _48588_ (_25223_, _25222_, _25221_);
  and _48589_ (_25224_, _25185_, _02385_);
  nor _48590_ (_25225_, _25185_, _02385_);
  or _48591_ (_25226_, _25225_, _25224_);
  nor _48592_ (_25227_, _25180_, _02380_);
  and _48593_ (_25228_, _25180_, _02380_);
  or _48594_ (_25229_, _25228_, _25227_);
  nor _48595_ (_25230_, _25170_, _00271_);
  and _48596_ (_25231_, _25170_, _00271_);
  or _48597_ (_25232_, _25231_, _25230_);
  nor _48598_ (_25233_, _25165_, _00241_);
  and _48599_ (_25234_, _25165_, _00241_);
  or _48600_ (_25235_, _25234_, _25233_);
  nor _48601_ (_25236_, _25160_, _00220_);
  and _48602_ (_25237_, _25160_, _00220_);
  or _48603_ (_25238_, _25237_, _25236_);
  and _48604_ (_25239_, _25150_, _00202_);
  nor _48605_ (_25240_, _25150_, _00202_);
  or _48606_ (_25241_, _25240_, _25239_);
  and _48607_ (_25242_, _25141_, _00299_);
  nor _48608_ (_25243_, \uc8051golden_1.PC [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _48609_ (_25244_, \uc8051golden_1.PC [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _48610_ (_25245_, _25244_, _25243_);
  nor _48611_ (_25246_, _25141_, _00299_);
  or _48612_ (_25247_, _25246_, _25245_);
  or _48613_ (_25248_, _25247_, _25242_);
  and _48614_ (_25249_, _25146_, _00317_);
  nor _48615_ (_25250_, _25146_, _00317_);
  or _48616_ (_25251_, _25250_, _25249_);
  or _48617_ (_25252_, _25251_, _25248_);
  or _48618_ (_25253_, _25252_, _25241_);
  nor _48619_ (_25254_, _25155_, _00031_);
  and _48620_ (_25255_, _25155_, _00031_);
  or _48621_ (_25256_, _25255_, _25254_);
  or _48622_ (_25257_, _25256_, _25253_);
  or _48623_ (_25258_, _25257_, _25238_);
  or _48624_ (_25259_, _25258_, _25235_);
  or _48625_ (_25260_, _25259_, _25232_);
  nor _48626_ (_25261_, _25175_, _02374_);
  and _48627_ (_25262_, _25175_, _02374_);
  or _48628_ (_25263_, _25262_, _25261_);
  or _48629_ (_25264_, _25263_, _25260_);
  or _48630_ (_25265_, _25264_, _25229_);
  or _48631_ (_25266_, _25265_, _25226_);
  or _48632_ (_25267_, _25266_, _25223_);
  or _48633_ (_25268_, _25267_, _25220_);
  or _48634_ (_25269_, _25268_, _25217_);
  or _48635_ (_25270_, _25269_, _25214_);
  or _48636_ (_25271_, _25270_, _25211_);
  and _48637_ (property_invalid_pc, _25271_, _22345_);
  buf _48638_ (_00488_, _25366_);
  buf _48639_ (_02668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7]);
  buf _48640_ (_14681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0]);
  buf _48641_ (_14683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1]);
  buf _48642_ (_14684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2]);
  buf _48643_ (_14685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3]);
  buf _48644_ (_14687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4]);
  buf _48645_ (_14688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5]);
  buf _48646_ (_14689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6]);
  buf _48647_ (_06116_, _06080_);
  buf _48648_ (_06117_, _06081_);
  buf _48649_ (_06128_, _06080_);
  buf _48650_ (_06129_, _06081_);
  buf _48651_ (_06242_, _06090_);
  buf _48652_ (_06243_, _06091_);
  buf _48653_ (_06244_, _06092_);
  buf _48654_ (_06245_, _06093_);
  buf _48655_ (_06246_, _06094_);
  buf _48656_ (_06247_, _06096_);
  buf _48657_ (_06248_, _06097_);
  buf _48658_ (_06249_, _06098_);
  buf _48659_ (_06250_, _06099_);
  buf _48660_ (_06251_, _06100_);
  buf _48661_ (_06252_, _06101_);
  buf _48662_ (_06253_, _06102_);
  buf _48663_ (_06254_, _06103_);
  buf _48664_ (_06255_, _06104_);
  buf _48665_ (_06303_, _06090_);
  buf _48666_ (_06304_, _06091_);
  buf _48667_ (_06305_, _06092_);
  buf _48668_ (_06306_, _06093_);
  buf _48669_ (_06307_, _06094_);
  buf _48670_ (_06308_, _06096_);
  buf _48671_ (_06309_, _06097_);
  buf _48672_ (_06310_, _06098_);
  buf _48673_ (_06311_, _06099_);
  buf _48674_ (_06312_, _06100_);
  buf _48675_ (_06313_, _06101_);
  buf _48676_ (_06314_, _06102_);
  buf _48677_ (_06315_, _06103_);
  buf _48678_ (_06316_, _06104_);
  buf _48679_ (_06506_, _06419_);
  buf _48680_ (_06535_, _06419_);
  buf _48681_ (_06583_, \uc8051golden_1.IRAM[255] [7]);
  buf _48682_ (_06726_, \uc8051golden_1.IRAM[0] [0]);
  buf _48683_ (_06727_, \uc8051golden_1.IRAM[0] [1]);
  buf _48684_ (_06728_, \uc8051golden_1.IRAM[0] [2]);
  buf _48685_ (_06729_, \uc8051golden_1.IRAM[0] [3]);
  buf _48686_ (_06730_, \uc8051golden_1.IRAM[0] [4]);
  buf _48687_ (_06731_, \uc8051golden_1.IRAM[0] [5]);
  buf _48688_ (_06732_, \uc8051golden_1.IRAM[0] [6]);
  buf _48689_ (_06733_, \uc8051golden_1.IRAM[0] [7]);
  buf _48690_ (_06734_, \uc8051golden_1.IRAM[1] [0]);
  buf _48691_ (_06735_, \uc8051golden_1.IRAM[1] [1]);
  buf _48692_ (_06736_, \uc8051golden_1.IRAM[1] [2]);
  buf _48693_ (_06737_, \uc8051golden_1.IRAM[1] [3]);
  buf _48694_ (_06738_, \uc8051golden_1.IRAM[1] [4]);
  buf _48695_ (_06739_, \uc8051golden_1.IRAM[1] [5]);
  buf _48696_ (_06740_, \uc8051golden_1.IRAM[1] [6]);
  buf _48697_ (_06741_, \uc8051golden_1.IRAM[1] [7]);
  buf _48698_ (_06742_, \uc8051golden_1.IRAM[2] [0]);
  buf _48699_ (_06743_, \uc8051golden_1.IRAM[2] [1]);
  buf _48700_ (_06744_, \uc8051golden_1.IRAM[2] [2]);
  buf _48701_ (_06746_, \uc8051golden_1.IRAM[2] [3]);
  buf _48702_ (_06747_, \uc8051golden_1.IRAM[2] [4]);
  buf _48703_ (_06748_, \uc8051golden_1.IRAM[2] [5]);
  buf _48704_ (_06749_, \uc8051golden_1.IRAM[2] [6]);
  buf _48705_ (_06750_, \uc8051golden_1.IRAM[2] [7]);
  buf _48706_ (_06751_, \uc8051golden_1.IRAM[3] [0]);
  buf _48707_ (_06752_, \uc8051golden_1.IRAM[3] [1]);
  buf _48708_ (_06753_, \uc8051golden_1.IRAM[3] [2]);
  buf _48709_ (_06754_, \uc8051golden_1.IRAM[3] [3]);
  buf _48710_ (_06755_, \uc8051golden_1.IRAM[3] [4]);
  buf _48711_ (_06756_, \uc8051golden_1.IRAM[3] [5]);
  buf _48712_ (_06757_, \uc8051golden_1.IRAM[3] [6]);
  buf _48713_ (_06758_, \uc8051golden_1.IRAM[3] [7]);
  buf _48714_ (_06759_, \uc8051golden_1.IRAM[4] [0]);
  buf _48715_ (_06760_, \uc8051golden_1.IRAM[4] [1]);
  buf _48716_ (_06761_, \uc8051golden_1.IRAM[4] [2]);
  buf _48717_ (_06762_, \uc8051golden_1.IRAM[4] [3]);
  buf _48718_ (_06763_, \uc8051golden_1.IRAM[4] [4]);
  buf _48719_ (_06764_, \uc8051golden_1.IRAM[4] [5]);
  buf _48720_ (_06765_, \uc8051golden_1.IRAM[4] [6]);
  buf _48721_ (_06766_, \uc8051golden_1.IRAM[4] [7]);
  buf _48722_ (_06767_, \uc8051golden_1.IRAM[5] [0]);
  buf _48723_ (_06768_, \uc8051golden_1.IRAM[5] [1]);
  buf _48724_ (_06769_, \uc8051golden_1.IRAM[5] [2]);
  buf _48725_ (_06770_, \uc8051golden_1.IRAM[5] [3]);
  buf _48726_ (_06771_, \uc8051golden_1.IRAM[5] [4]);
  buf _48727_ (_06772_, \uc8051golden_1.IRAM[5] [5]);
  buf _48728_ (_06773_, \uc8051golden_1.IRAM[5] [6]);
  buf _48729_ (_06774_, \uc8051golden_1.IRAM[5] [7]);
  buf _48730_ (_06775_, \uc8051golden_1.IRAM[6] [0]);
  buf _48731_ (_06776_, \uc8051golden_1.IRAM[6] [1]);
  buf _48732_ (_06778_, \uc8051golden_1.IRAM[6] [2]);
  buf _48733_ (_06779_, \uc8051golden_1.IRAM[6] [3]);
  buf _48734_ (_06780_, \uc8051golden_1.IRAM[6] [4]);
  buf _48735_ (_06781_, \uc8051golden_1.IRAM[6] [5]);
  buf _48736_ (_06782_, \uc8051golden_1.IRAM[6] [6]);
  buf _48737_ (_06783_, \uc8051golden_1.IRAM[6] [7]);
  buf _48738_ (_06784_, \uc8051golden_1.IRAM[7] [0]);
  buf _48739_ (_06785_, \uc8051golden_1.IRAM[7] [1]);
  buf _48740_ (_06786_, \uc8051golden_1.IRAM[7] [2]);
  buf _48741_ (_06787_, \uc8051golden_1.IRAM[7] [3]);
  buf _48742_ (_06788_, \uc8051golden_1.IRAM[7] [4]);
  buf _48743_ (_06789_, \uc8051golden_1.IRAM[7] [5]);
  buf _48744_ (_06790_, \uc8051golden_1.IRAM[7] [6]);
  buf _48745_ (_06791_, \uc8051golden_1.IRAM[7] [7]);
  buf _48746_ (_06792_, \uc8051golden_1.IRAM[8] [0]);
  buf _48747_ (_06793_, \uc8051golden_1.IRAM[8] [1]);
  buf _48748_ (_06794_, \uc8051golden_1.IRAM[8] [2]);
  buf _48749_ (_06795_, \uc8051golden_1.IRAM[8] [3]);
  buf _48750_ (_06796_, \uc8051golden_1.IRAM[8] [4]);
  buf _48751_ (_06797_, \uc8051golden_1.IRAM[8] [5]);
  buf _48752_ (_06798_, \uc8051golden_1.IRAM[8] [6]);
  buf _48753_ (_06799_, \uc8051golden_1.IRAM[8] [7]);
  buf _48754_ (_06800_, \uc8051golden_1.IRAM[9] [0]);
  buf _48755_ (_06801_, \uc8051golden_1.IRAM[9] [1]);
  buf _48756_ (_06802_, \uc8051golden_1.IRAM[9] [2]);
  buf _48757_ (_06803_, \uc8051golden_1.IRAM[9] [3]);
  buf _48758_ (_06804_, \uc8051golden_1.IRAM[9] [4]);
  buf _48759_ (_06805_, \uc8051golden_1.IRAM[9] [5]);
  buf _48760_ (_06806_, \uc8051golden_1.IRAM[9] [6]);
  buf _48761_ (_06807_, \uc8051golden_1.IRAM[9] [7]);
  buf _48762_ (_06808_, \uc8051golden_1.IRAM[10] [0]);
  buf _48763_ (_06810_, \uc8051golden_1.IRAM[10] [1]);
  buf _48764_ (_06811_, \uc8051golden_1.IRAM[10] [2]);
  buf _48765_ (_06812_, \uc8051golden_1.IRAM[10] [3]);
  buf _48766_ (_06813_, \uc8051golden_1.IRAM[10] [4]);
  buf _48767_ (_06814_, \uc8051golden_1.IRAM[10] [5]);
  buf _48768_ (_06815_, \uc8051golden_1.IRAM[10] [6]);
  buf _48769_ (_06816_, \uc8051golden_1.IRAM[10] [7]);
  buf _48770_ (_06817_, \uc8051golden_1.IRAM[11] [0]);
  buf _48771_ (_06818_, \uc8051golden_1.IRAM[11] [1]);
  buf _48772_ (_06819_, \uc8051golden_1.IRAM[11] [2]);
  buf _48773_ (_06820_, \uc8051golden_1.IRAM[11] [3]);
  buf _48774_ (_06821_, \uc8051golden_1.IRAM[11] [4]);
  buf _48775_ (_06822_, \uc8051golden_1.IRAM[11] [5]);
  buf _48776_ (_06823_, \uc8051golden_1.IRAM[11] [6]);
  buf _48777_ (_06824_, \uc8051golden_1.IRAM[11] [7]);
  buf _48778_ (_06825_, \uc8051golden_1.IRAM[12] [0]);
  buf _48779_ (_06826_, \uc8051golden_1.IRAM[12] [1]);
  buf _48780_ (_06827_, \uc8051golden_1.IRAM[12] [2]);
  buf _48781_ (_06828_, \uc8051golden_1.IRAM[12] [3]);
  buf _48782_ (_06829_, \uc8051golden_1.IRAM[12] [4]);
  buf _48783_ (_06830_, \uc8051golden_1.IRAM[12] [5]);
  buf _48784_ (_06831_, \uc8051golden_1.IRAM[12] [6]);
  buf _48785_ (_06832_, \uc8051golden_1.IRAM[12] [7]);
  buf _48786_ (_06833_, \uc8051golden_1.IRAM[13] [0]);
  buf _48787_ (_06834_, \uc8051golden_1.IRAM[13] [1]);
  buf _48788_ (_06835_, \uc8051golden_1.IRAM[13] [2]);
  buf _48789_ (_06836_, \uc8051golden_1.IRAM[13] [3]);
  buf _48790_ (_06837_, \uc8051golden_1.IRAM[13] [4]);
  buf _48791_ (_06838_, \uc8051golden_1.IRAM[13] [5]);
  buf _48792_ (_06839_, \uc8051golden_1.IRAM[13] [6]);
  buf _48793_ (_06840_, \uc8051golden_1.IRAM[13] [7]);
  buf _48794_ (_06841_, \uc8051golden_1.IRAM[14] [0]);
  buf _48795_ (_06843_, \uc8051golden_1.IRAM[14] [1]);
  buf _48796_ (_06844_, \uc8051golden_1.IRAM[14] [2]);
  buf _48797_ (_06845_, \uc8051golden_1.IRAM[14] [3]);
  buf _48798_ (_06846_, \uc8051golden_1.IRAM[14] [4]);
  buf _48799_ (_06847_, \uc8051golden_1.IRAM[14] [5]);
  buf _48800_ (_06848_, \uc8051golden_1.IRAM[14] [6]);
  buf _48801_ (_06849_, \uc8051golden_1.IRAM[14] [7]);
  buf _48802_ (_06850_, \uc8051golden_1.IRAM[15] [0]);
  buf _48803_ (_06851_, \uc8051golden_1.IRAM[15] [1]);
  buf _48804_ (_06852_, \uc8051golden_1.IRAM[15] [2]);
  buf _48805_ (_06853_, \uc8051golden_1.IRAM[15] [3]);
  buf _48806_ (_06854_, \uc8051golden_1.IRAM[15] [4]);
  buf _48807_ (_06855_, \uc8051golden_1.IRAM[15] [5]);
  buf _48808_ (_06856_, \uc8051golden_1.IRAM[15] [6]);
  buf _48809_ (_06857_, \uc8051golden_1.IRAM[15] [7]);
  buf _48810_ (_06858_, \uc8051golden_1.IRAM[16] [0]);
  buf _48811_ (_06859_, \uc8051golden_1.IRAM[16] [1]);
  buf _48812_ (_06860_, \uc8051golden_1.IRAM[16] [2]);
  buf _48813_ (_06861_, \uc8051golden_1.IRAM[16] [3]);
  buf _48814_ (_06862_, \uc8051golden_1.IRAM[16] [4]);
  buf _48815_ (_06863_, \uc8051golden_1.IRAM[16] [5]);
  buf _48816_ (_06864_, \uc8051golden_1.IRAM[16] [6]);
  buf _48817_ (_06865_, \uc8051golden_1.IRAM[16] [7]);
  buf _48818_ (_06866_, \uc8051golden_1.IRAM[17] [0]);
  buf _48819_ (_06867_, \uc8051golden_1.IRAM[17] [1]);
  buf _48820_ (_06868_, \uc8051golden_1.IRAM[17] [2]);
  buf _48821_ (_06869_, \uc8051golden_1.IRAM[17] [3]);
  buf _48822_ (_06870_, \uc8051golden_1.IRAM[17] [4]);
  buf _48823_ (_06871_, \uc8051golden_1.IRAM[17] [5]);
  buf _48824_ (_06872_, \uc8051golden_1.IRAM[17] [6]);
  buf _48825_ (_06873_, \uc8051golden_1.IRAM[17] [7]);
  buf _48826_ (_06875_, \uc8051golden_1.IRAM[18] [0]);
  buf _48827_ (_06876_, \uc8051golden_1.IRAM[18] [1]);
  buf _48828_ (_06877_, \uc8051golden_1.IRAM[18] [2]);
  buf _48829_ (_06878_, \uc8051golden_1.IRAM[18] [3]);
  buf _48830_ (_06879_, \uc8051golden_1.IRAM[18] [4]);
  buf _48831_ (_06880_, \uc8051golden_1.IRAM[18] [5]);
  buf _48832_ (_06881_, \uc8051golden_1.IRAM[18] [6]);
  buf _48833_ (_06882_, \uc8051golden_1.IRAM[18] [7]);
  buf _48834_ (_06883_, \uc8051golden_1.IRAM[19] [0]);
  buf _48835_ (_06884_, \uc8051golden_1.IRAM[19] [1]);
  buf _48836_ (_06885_, \uc8051golden_1.IRAM[19] [2]);
  buf _48837_ (_06886_, \uc8051golden_1.IRAM[19] [3]);
  buf _48838_ (_06887_, \uc8051golden_1.IRAM[19] [4]);
  buf _48839_ (_06888_, \uc8051golden_1.IRAM[19] [5]);
  buf _48840_ (_06889_, \uc8051golden_1.IRAM[19] [6]);
  buf _48841_ (_06890_, \uc8051golden_1.IRAM[19] [7]);
  buf _48842_ (_06891_, \uc8051golden_1.IRAM[20] [0]);
  buf _48843_ (_06892_, \uc8051golden_1.IRAM[20] [1]);
  buf _48844_ (_06893_, \uc8051golden_1.IRAM[20] [2]);
  buf _48845_ (_06894_, \uc8051golden_1.IRAM[20] [3]);
  buf _48846_ (_06895_, \uc8051golden_1.IRAM[20] [4]);
  buf _48847_ (_06896_, \uc8051golden_1.IRAM[20] [5]);
  buf _48848_ (_06897_, \uc8051golden_1.IRAM[20] [6]);
  buf _48849_ (_06898_, \uc8051golden_1.IRAM[20] [7]);
  buf _48850_ (_06899_, \uc8051golden_1.IRAM[21] [0]);
  buf _48851_ (_06900_, \uc8051golden_1.IRAM[21] [1]);
  buf _48852_ (_06901_, \uc8051golden_1.IRAM[21] [2]);
  buf _48853_ (_06902_, \uc8051golden_1.IRAM[21] [3]);
  buf _48854_ (_06903_, \uc8051golden_1.IRAM[21] [4]);
  buf _48855_ (_06904_, \uc8051golden_1.IRAM[21] [5]);
  buf _48856_ (_06905_, \uc8051golden_1.IRAM[21] [6]);
  buf _48857_ (_06906_, \uc8051golden_1.IRAM[21] [7]);
  buf _48858_ (_06907_, \uc8051golden_1.IRAM[22] [0]);
  buf _48859_ (_06908_, \uc8051golden_1.IRAM[22] [1]);
  buf _48860_ (_06910_, \uc8051golden_1.IRAM[22] [2]);
  buf _48861_ (_06911_, \uc8051golden_1.IRAM[22] [3]);
  buf _48862_ (_06912_, \uc8051golden_1.IRAM[22] [4]);
  buf _48863_ (_06913_, \uc8051golden_1.IRAM[22] [5]);
  buf _48864_ (_06914_, \uc8051golden_1.IRAM[22] [6]);
  buf _48865_ (_06915_, \uc8051golden_1.IRAM[22] [7]);
  buf _48866_ (_06916_, \uc8051golden_1.IRAM[23] [0]);
  buf _48867_ (_06917_, \uc8051golden_1.IRAM[23] [1]);
  buf _48868_ (_06918_, \uc8051golden_1.IRAM[23] [2]);
  buf _48869_ (_06919_, \uc8051golden_1.IRAM[23] [3]);
  buf _48870_ (_06920_, \uc8051golden_1.IRAM[23] [4]);
  buf _48871_ (_06921_, \uc8051golden_1.IRAM[23] [5]);
  buf _48872_ (_06922_, \uc8051golden_1.IRAM[23] [6]);
  buf _48873_ (_06923_, \uc8051golden_1.IRAM[23] [7]);
  buf _48874_ (_06924_, \uc8051golden_1.IRAM[24] [0]);
  buf _48875_ (_06925_, \uc8051golden_1.IRAM[24] [1]);
  buf _48876_ (_06926_, \uc8051golden_1.IRAM[24] [2]);
  buf _48877_ (_06927_, \uc8051golden_1.IRAM[24] [3]);
  buf _48878_ (_06928_, \uc8051golden_1.IRAM[24] [4]);
  buf _48879_ (_06929_, \uc8051golden_1.IRAM[24] [5]);
  buf _48880_ (_06930_, \uc8051golden_1.IRAM[24] [6]);
  buf _48881_ (_06931_, \uc8051golden_1.IRAM[24] [7]);
  buf _48882_ (_06932_, \uc8051golden_1.IRAM[25] [0]);
  buf _48883_ (_06933_, \uc8051golden_1.IRAM[25] [1]);
  buf _48884_ (_06934_, \uc8051golden_1.IRAM[25] [2]);
  buf _48885_ (_06935_, \uc8051golden_1.IRAM[25] [3]);
  buf _48886_ (_06936_, \uc8051golden_1.IRAM[25] [4]);
  buf _48887_ (_06937_, \uc8051golden_1.IRAM[25] [5]);
  buf _48888_ (_06938_, \uc8051golden_1.IRAM[25] [6]);
  buf _48889_ (_06939_, \uc8051golden_1.IRAM[25] [7]);
  buf _48890_ (_06940_, \uc8051golden_1.IRAM[26] [0]);
  buf _48891_ (_06941_, \uc8051golden_1.IRAM[26] [1]);
  buf _48892_ (_06942_, \uc8051golden_1.IRAM[26] [2]);
  buf _48893_ (_06944_, \uc8051golden_1.IRAM[26] [3]);
  buf _48894_ (_06945_, \uc8051golden_1.IRAM[26] [4]);
  buf _48895_ (_06946_, \uc8051golden_1.IRAM[26] [5]);
  buf _48896_ (_06947_, \uc8051golden_1.IRAM[26] [6]);
  buf _48897_ (_06948_, \uc8051golden_1.IRAM[26] [7]);
  buf _48898_ (_06949_, \uc8051golden_1.IRAM[27] [0]);
  buf _48899_ (_06950_, \uc8051golden_1.IRAM[27] [1]);
  buf _48900_ (_06951_, \uc8051golden_1.IRAM[27] [2]);
  buf _48901_ (_06952_, \uc8051golden_1.IRAM[27] [3]);
  buf _48902_ (_06953_, \uc8051golden_1.IRAM[27] [4]);
  buf _48903_ (_06954_, \uc8051golden_1.IRAM[27] [5]);
  buf _48904_ (_06955_, \uc8051golden_1.IRAM[27] [6]);
  buf _48905_ (_06956_, \uc8051golden_1.IRAM[27] [7]);
  buf _48906_ (_06957_, \uc8051golden_1.IRAM[28] [0]);
  buf _48907_ (_06958_, \uc8051golden_1.IRAM[28] [1]);
  buf _48908_ (_06959_, \uc8051golden_1.IRAM[28] [2]);
  buf _48909_ (_06960_, \uc8051golden_1.IRAM[28] [3]);
  buf _48910_ (_06961_, \uc8051golden_1.IRAM[28] [4]);
  buf _48911_ (_06962_, \uc8051golden_1.IRAM[28] [5]);
  buf _48912_ (_06963_, \uc8051golden_1.IRAM[28] [6]);
  buf _48913_ (_06964_, \uc8051golden_1.IRAM[28] [7]);
  buf _48914_ (_06965_, \uc8051golden_1.IRAM[29] [0]);
  buf _48915_ (_06966_, \uc8051golden_1.IRAM[29] [1]);
  buf _48916_ (_06967_, \uc8051golden_1.IRAM[29] [2]);
  buf _48917_ (_06968_, \uc8051golden_1.IRAM[29] [3]);
  buf _48918_ (_06969_, \uc8051golden_1.IRAM[29] [4]);
  buf _48919_ (_06970_, \uc8051golden_1.IRAM[29] [5]);
  buf _48920_ (_06971_, \uc8051golden_1.IRAM[29] [6]);
  buf _48921_ (_06972_, \uc8051golden_1.IRAM[29] [7]);
  buf _48922_ (_06973_, \uc8051golden_1.IRAM[30] [0]);
  buf _48923_ (_06974_, \uc8051golden_1.IRAM[30] [1]);
  buf _48924_ (_06975_, \uc8051golden_1.IRAM[30] [2]);
  buf _48925_ (_06976_, \uc8051golden_1.IRAM[30] [3]);
  buf _48926_ (_06978_, \uc8051golden_1.IRAM[30] [4]);
  buf _48927_ (_06979_, \uc8051golden_1.IRAM[30] [5]);
  buf _48928_ (_06980_, \uc8051golden_1.IRAM[30] [6]);
  buf _48929_ (_06981_, \uc8051golden_1.IRAM[30] [7]);
  buf _48930_ (_06982_, \uc8051golden_1.IRAM[31] [0]);
  buf _48931_ (_06983_, \uc8051golden_1.IRAM[31] [1]);
  buf _48932_ (_06984_, \uc8051golden_1.IRAM[31] [2]);
  buf _48933_ (_06985_, \uc8051golden_1.IRAM[31] [3]);
  buf _48934_ (_06986_, \uc8051golden_1.IRAM[31] [4]);
  buf _48935_ (_06987_, \uc8051golden_1.IRAM[31] [5]);
  buf _48936_ (_06988_, \uc8051golden_1.IRAM[31] [6]);
  buf _48937_ (_06989_, \uc8051golden_1.IRAM[31] [7]);
  buf _48938_ (_06990_, \uc8051golden_1.IRAM[32] [0]);
  buf _48939_ (_06991_, \uc8051golden_1.IRAM[32] [1]);
  buf _48940_ (_06992_, \uc8051golden_1.IRAM[32] [2]);
  buf _48941_ (_06993_, \uc8051golden_1.IRAM[32] [3]);
  buf _48942_ (_06994_, \uc8051golden_1.IRAM[32] [4]);
  buf _48943_ (_06995_, \uc8051golden_1.IRAM[32] [5]);
  buf _48944_ (_06996_, \uc8051golden_1.IRAM[32] [6]);
  buf _48945_ (_06997_, \uc8051golden_1.IRAM[32] [7]);
  buf _48946_ (_06998_, \uc8051golden_1.IRAM[33] [0]);
  buf _48947_ (_06999_, \uc8051golden_1.IRAM[33] [1]);
  buf _48948_ (_07000_, \uc8051golden_1.IRAM[33] [2]);
  buf _48949_ (_07001_, \uc8051golden_1.IRAM[33] [3]);
  buf _48950_ (_07002_, \uc8051golden_1.IRAM[33] [4]);
  buf _48951_ (_07003_, \uc8051golden_1.IRAM[33] [5]);
  buf _48952_ (_07004_, \uc8051golden_1.IRAM[33] [6]);
  buf _48953_ (_07005_, \uc8051golden_1.IRAM[33] [7]);
  buf _48954_ (_07006_, \uc8051golden_1.IRAM[34] [0]);
  buf _48955_ (_07007_, \uc8051golden_1.IRAM[34] [1]);
  buf _48956_ (_07008_, \uc8051golden_1.IRAM[34] [2]);
  buf _48957_ (_07009_, \uc8051golden_1.IRAM[34] [3]);
  buf _48958_ (_07011_, \uc8051golden_1.IRAM[34] [4]);
  buf _48959_ (_07012_, \uc8051golden_1.IRAM[34] [5]);
  buf _48960_ (_07013_, \uc8051golden_1.IRAM[34] [6]);
  buf _48961_ (_07014_, \uc8051golden_1.IRAM[34] [7]);
  buf _48962_ (_07015_, \uc8051golden_1.IRAM[35] [0]);
  buf _48963_ (_07016_, \uc8051golden_1.IRAM[35] [1]);
  buf _48964_ (_07017_, \uc8051golden_1.IRAM[35] [2]);
  buf _48965_ (_07018_, \uc8051golden_1.IRAM[35] [3]);
  buf _48966_ (_07019_, \uc8051golden_1.IRAM[35] [4]);
  buf _48967_ (_07020_, \uc8051golden_1.IRAM[35] [5]);
  buf _48968_ (_07021_, \uc8051golden_1.IRAM[35] [6]);
  buf _48969_ (_07022_, \uc8051golden_1.IRAM[35] [7]);
  buf _48970_ (_07023_, \uc8051golden_1.IRAM[36] [0]);
  buf _48971_ (_07024_, \uc8051golden_1.IRAM[36] [1]);
  buf _48972_ (_07025_, \uc8051golden_1.IRAM[36] [2]);
  buf _48973_ (_07026_, \uc8051golden_1.IRAM[36] [3]);
  buf _48974_ (_07027_, \uc8051golden_1.IRAM[36] [4]);
  buf _48975_ (_07028_, \uc8051golden_1.IRAM[36] [5]);
  buf _48976_ (_07029_, \uc8051golden_1.IRAM[36] [6]);
  buf _48977_ (_07030_, \uc8051golden_1.IRAM[36] [7]);
  buf _48978_ (_07031_, \uc8051golden_1.IRAM[37] [0]);
  buf _48979_ (_07032_, \uc8051golden_1.IRAM[37] [1]);
  buf _48980_ (_07033_, \uc8051golden_1.IRAM[37] [2]);
  buf _48981_ (_07034_, \uc8051golden_1.IRAM[37] [3]);
  buf _48982_ (_07035_, \uc8051golden_1.IRAM[37] [4]);
  buf _48983_ (_07036_, \uc8051golden_1.IRAM[37] [5]);
  buf _48984_ (_07037_, \uc8051golden_1.IRAM[37] [6]);
  buf _48985_ (_07038_, \uc8051golden_1.IRAM[37] [7]);
  buf _48986_ (_07039_, \uc8051golden_1.IRAM[38] [0]);
  buf _48987_ (_07040_, \uc8051golden_1.IRAM[38] [1]);
  buf _48988_ (_07041_, \uc8051golden_1.IRAM[38] [2]);
  buf _48989_ (_07042_, \uc8051golden_1.IRAM[38] [3]);
  buf _48990_ (_07043_, \uc8051golden_1.IRAM[38] [4]);
  buf _48991_ (_07044_, \uc8051golden_1.IRAM[38] [5]);
  buf _48992_ (_07046_, \uc8051golden_1.IRAM[38] [6]);
  buf _48993_ (_07047_, \uc8051golden_1.IRAM[38] [7]);
  buf _48994_ (_07048_, \uc8051golden_1.IRAM[39] [0]);
  buf _48995_ (_07049_, \uc8051golden_1.IRAM[39] [1]);
  buf _48996_ (_07050_, \uc8051golden_1.IRAM[39] [2]);
  buf _48997_ (_07051_, \uc8051golden_1.IRAM[39] [3]);
  buf _48998_ (_07052_, \uc8051golden_1.IRAM[39] [4]);
  buf _48999_ (_07053_, \uc8051golden_1.IRAM[39] [5]);
  buf _49000_ (_07054_, \uc8051golden_1.IRAM[39] [6]);
  buf _49001_ (_07055_, \uc8051golden_1.IRAM[39] [7]);
  buf _49002_ (_07056_, \uc8051golden_1.IRAM[40] [0]);
  buf _49003_ (_07057_, \uc8051golden_1.IRAM[40] [1]);
  buf _49004_ (_07058_, \uc8051golden_1.IRAM[40] [2]);
  buf _49005_ (_07059_, \uc8051golden_1.IRAM[40] [3]);
  buf _49006_ (_07060_, \uc8051golden_1.IRAM[40] [4]);
  buf _49007_ (_07061_, \uc8051golden_1.IRAM[40] [5]);
  buf _49008_ (_07062_, \uc8051golden_1.IRAM[40] [6]);
  buf _49009_ (_07063_, \uc8051golden_1.IRAM[40] [7]);
  buf _49010_ (_07064_, \uc8051golden_1.IRAM[41] [0]);
  buf _49011_ (_07065_, \uc8051golden_1.IRAM[41] [1]);
  buf _49012_ (_07066_, \uc8051golden_1.IRAM[41] [2]);
  buf _49013_ (_07067_, \uc8051golden_1.IRAM[41] [3]);
  buf _49014_ (_07068_, \uc8051golden_1.IRAM[41] [4]);
  buf _49015_ (_07069_, \uc8051golden_1.IRAM[41] [5]);
  buf _49016_ (_07070_, \uc8051golden_1.IRAM[41] [6]);
  buf _49017_ (_07071_, \uc8051golden_1.IRAM[41] [7]);
  buf _49018_ (_07072_, \uc8051golden_1.IRAM[42] [0]);
  buf _49019_ (_07073_, \uc8051golden_1.IRAM[42] [1]);
  buf _49020_ (_07074_, \uc8051golden_1.IRAM[42] [2]);
  buf _49021_ (_07075_, \uc8051golden_1.IRAM[42] [3]);
  buf _49022_ (_07076_, \uc8051golden_1.IRAM[42] [4]);
  buf _49023_ (_07077_, \uc8051golden_1.IRAM[42] [5]);
  buf _49024_ (_07078_, \uc8051golden_1.IRAM[42] [6]);
  buf _49025_ (_07080_, \uc8051golden_1.IRAM[42] [7]);
  buf _49026_ (_07081_, \uc8051golden_1.IRAM[43] [0]);
  buf _49027_ (_07082_, \uc8051golden_1.IRAM[43] [1]);
  buf _49028_ (_07083_, \uc8051golden_1.IRAM[43] [2]);
  buf _49029_ (_07084_, \uc8051golden_1.IRAM[43] [3]);
  buf _49030_ (_07085_, \uc8051golden_1.IRAM[43] [4]);
  buf _49031_ (_07086_, \uc8051golden_1.IRAM[43] [5]);
  buf _49032_ (_07087_, \uc8051golden_1.IRAM[43] [6]);
  buf _49033_ (_07088_, \uc8051golden_1.IRAM[43] [7]);
  buf _49034_ (_07089_, \uc8051golden_1.IRAM[44] [0]);
  buf _49035_ (_07090_, \uc8051golden_1.IRAM[44] [1]);
  buf _49036_ (_07091_, \uc8051golden_1.IRAM[44] [2]);
  buf _49037_ (_07092_, \uc8051golden_1.IRAM[44] [3]);
  buf _49038_ (_07093_, \uc8051golden_1.IRAM[44] [4]);
  buf _49039_ (_07094_, \uc8051golden_1.IRAM[44] [5]);
  buf _49040_ (_07095_, \uc8051golden_1.IRAM[44] [6]);
  buf _49041_ (_07096_, \uc8051golden_1.IRAM[44] [7]);
  buf _49042_ (_07097_, \uc8051golden_1.IRAM[45] [0]);
  buf _49043_ (_07098_, \uc8051golden_1.IRAM[45] [1]);
  buf _49044_ (_07099_, \uc8051golden_1.IRAM[45] [2]);
  buf _49045_ (_07100_, \uc8051golden_1.IRAM[45] [3]);
  buf _49046_ (_07101_, \uc8051golden_1.IRAM[45] [4]);
  buf _49047_ (_07102_, \uc8051golden_1.IRAM[45] [5]);
  buf _49048_ (_07103_, \uc8051golden_1.IRAM[45] [6]);
  buf _49049_ (_07104_, \uc8051golden_1.IRAM[45] [7]);
  buf _49050_ (_07105_, \uc8051golden_1.IRAM[46] [0]);
  buf _49051_ (_07106_, \uc8051golden_1.IRAM[46] [1]);
  buf _49052_ (_07107_, \uc8051golden_1.IRAM[46] [2]);
  buf _49053_ (_07108_, \uc8051golden_1.IRAM[46] [3]);
  buf _49054_ (_07109_, \uc8051golden_1.IRAM[46] [4]);
  buf _49055_ (_07110_, \uc8051golden_1.IRAM[46] [5]);
  buf _49056_ (_07111_, \uc8051golden_1.IRAM[46] [6]);
  buf _49057_ (_07112_, \uc8051golden_1.IRAM[46] [7]);
  buf _49058_ (_07114_, \uc8051golden_1.IRAM[47] [0]);
  buf _49059_ (_07115_, \uc8051golden_1.IRAM[47] [1]);
  buf _49060_ (_07116_, \uc8051golden_1.IRAM[47] [2]);
  buf _49061_ (_07117_, \uc8051golden_1.IRAM[47] [3]);
  buf _49062_ (_07118_, \uc8051golden_1.IRAM[47] [4]);
  buf _49063_ (_07119_, \uc8051golden_1.IRAM[47] [5]);
  buf _49064_ (_07120_, \uc8051golden_1.IRAM[47] [6]);
  buf _49065_ (_07121_, \uc8051golden_1.IRAM[47] [7]);
  buf _49066_ (_07122_, \uc8051golden_1.IRAM[48] [0]);
  buf _49067_ (_07123_, \uc8051golden_1.IRAM[48] [1]);
  buf _49068_ (_07124_, \uc8051golden_1.IRAM[48] [2]);
  buf _49069_ (_07125_, \uc8051golden_1.IRAM[48] [3]);
  buf _49070_ (_07126_, \uc8051golden_1.IRAM[48] [4]);
  buf _49071_ (_07127_, \uc8051golden_1.IRAM[48] [5]);
  buf _49072_ (_07128_, \uc8051golden_1.IRAM[48] [6]);
  buf _49073_ (_07129_, \uc8051golden_1.IRAM[48] [7]);
  buf _49074_ (_07130_, \uc8051golden_1.IRAM[49] [0]);
  buf _49075_ (_07131_, \uc8051golden_1.IRAM[49] [1]);
  buf _49076_ (_07132_, \uc8051golden_1.IRAM[49] [2]);
  buf _49077_ (_07133_, \uc8051golden_1.IRAM[49] [3]);
  buf _49078_ (_07134_, \uc8051golden_1.IRAM[49] [4]);
  buf _49079_ (_07135_, \uc8051golden_1.IRAM[49] [5]);
  buf _49080_ (_07136_, \uc8051golden_1.IRAM[49] [6]);
  buf _49081_ (_07137_, \uc8051golden_1.IRAM[49] [7]);
  buf _49082_ (_07138_, \uc8051golden_1.IRAM[50] [0]);
  buf _49083_ (_07139_, \uc8051golden_1.IRAM[50] [1]);
  buf _49084_ (_07140_, \uc8051golden_1.IRAM[50] [2]);
  buf _49085_ (_07141_, \uc8051golden_1.IRAM[50] [3]);
  buf _49086_ (_07142_, \uc8051golden_1.IRAM[50] [4]);
  buf _49087_ (_07143_, \uc8051golden_1.IRAM[50] [5]);
  buf _49088_ (_07144_, \uc8051golden_1.IRAM[50] [6]);
  buf _49089_ (_07145_, \uc8051golden_1.IRAM[50] [7]);
  buf _49090_ (_07146_, \uc8051golden_1.IRAM[51] [0]);
  buf _49091_ (_07148_, \uc8051golden_1.IRAM[51] [1]);
  buf _49092_ (_07149_, \uc8051golden_1.IRAM[51] [2]);
  buf _49093_ (_07150_, \uc8051golden_1.IRAM[51] [3]);
  buf _49094_ (_07151_, \uc8051golden_1.IRAM[51] [4]);
  buf _49095_ (_07152_, \uc8051golden_1.IRAM[51] [5]);
  buf _49096_ (_07153_, \uc8051golden_1.IRAM[51] [6]);
  buf _49097_ (_07154_, \uc8051golden_1.IRAM[51] [7]);
  buf _49098_ (_07155_, \uc8051golden_1.IRAM[52] [0]);
  buf _49099_ (_07156_, \uc8051golden_1.IRAM[52] [1]);
  buf _49100_ (_07157_, \uc8051golden_1.IRAM[52] [2]);
  buf _49101_ (_07158_, \uc8051golden_1.IRAM[52] [3]);
  buf _49102_ (_07159_, \uc8051golden_1.IRAM[52] [4]);
  buf _49103_ (_07160_, \uc8051golden_1.IRAM[52] [5]);
  buf _49104_ (_07161_, \uc8051golden_1.IRAM[52] [6]);
  buf _49105_ (_07162_, \uc8051golden_1.IRAM[52] [7]);
  buf _49106_ (_07163_, \uc8051golden_1.IRAM[53] [0]);
  buf _49107_ (_07164_, \uc8051golden_1.IRAM[53] [1]);
  buf _49108_ (_07165_, \uc8051golden_1.IRAM[53] [2]);
  buf _49109_ (_07166_, \uc8051golden_1.IRAM[53] [3]);
  buf _49110_ (_07167_, \uc8051golden_1.IRAM[53] [4]);
  buf _49111_ (_07168_, \uc8051golden_1.IRAM[53] [5]);
  buf _49112_ (_07169_, \uc8051golden_1.IRAM[53] [6]);
  buf _49113_ (_07170_, \uc8051golden_1.IRAM[53] [7]);
  buf _49114_ (_07171_, \uc8051golden_1.IRAM[54] [0]);
  buf _49115_ (_07172_, \uc8051golden_1.IRAM[54] [1]);
  buf _49116_ (_07173_, \uc8051golden_1.IRAM[54] [2]);
  buf _49117_ (_07174_, \uc8051golden_1.IRAM[54] [3]);
  buf _49118_ (_07175_, \uc8051golden_1.IRAM[54] [4]);
  buf _49119_ (_07176_, \uc8051golden_1.IRAM[54] [5]);
  buf _49120_ (_07177_, \uc8051golden_1.IRAM[54] [6]);
  buf _49121_ (_07178_, \uc8051golden_1.IRAM[54] [7]);
  buf _49122_ (_07179_, \uc8051golden_1.IRAM[55] [0]);
  buf _49123_ (_07180_, \uc8051golden_1.IRAM[55] [1]);
  buf _49124_ (_07182_, \uc8051golden_1.IRAM[55] [2]);
  buf _49125_ (_07183_, \uc8051golden_1.IRAM[55] [3]);
  buf _49126_ (_07184_, \uc8051golden_1.IRAM[55] [4]);
  buf _49127_ (_07185_, \uc8051golden_1.IRAM[55] [5]);
  buf _49128_ (_07186_, \uc8051golden_1.IRAM[55] [6]);
  buf _49129_ (_07187_, \uc8051golden_1.IRAM[55] [7]);
  buf _49130_ (_07188_, \uc8051golden_1.IRAM[56] [0]);
  buf _49131_ (_07189_, \uc8051golden_1.IRAM[56] [1]);
  buf _49132_ (_07190_, \uc8051golden_1.IRAM[56] [2]);
  buf _49133_ (_07191_, \uc8051golden_1.IRAM[56] [3]);
  buf _49134_ (_07192_, \uc8051golden_1.IRAM[56] [4]);
  buf _49135_ (_07193_, \uc8051golden_1.IRAM[56] [5]);
  buf _49136_ (_07194_, \uc8051golden_1.IRAM[56] [6]);
  buf _49137_ (_07195_, \uc8051golden_1.IRAM[56] [7]);
  buf _49138_ (_07196_, \uc8051golden_1.IRAM[57] [0]);
  buf _49139_ (_07197_, \uc8051golden_1.IRAM[57] [1]);
  buf _49140_ (_07198_, \uc8051golden_1.IRAM[57] [2]);
  buf _49141_ (_07199_, \uc8051golden_1.IRAM[57] [3]);
  buf _49142_ (_07200_, \uc8051golden_1.IRAM[57] [4]);
  buf _49143_ (_07201_, \uc8051golden_1.IRAM[57] [5]);
  buf _49144_ (_07202_, \uc8051golden_1.IRAM[57] [6]);
  buf _49145_ (_07203_, \uc8051golden_1.IRAM[57] [7]);
  buf _49146_ (_07204_, \uc8051golden_1.IRAM[58] [0]);
  buf _49147_ (_07205_, \uc8051golden_1.IRAM[58] [1]);
  buf _49148_ (_07206_, \uc8051golden_1.IRAM[58] [2]);
  buf _49149_ (_07207_, \uc8051golden_1.IRAM[58] [3]);
  buf _49150_ (_07208_, \uc8051golden_1.IRAM[58] [4]);
  buf _49151_ (_07209_, \uc8051golden_1.IRAM[58] [5]);
  buf _49152_ (_07210_, \uc8051golden_1.IRAM[58] [6]);
  buf _49153_ (_07211_, \uc8051golden_1.IRAM[58] [7]);
  buf _49154_ (_07212_, \uc8051golden_1.IRAM[59] [0]);
  buf _49155_ (_07213_, \uc8051golden_1.IRAM[59] [1]);
  buf _49156_ (_07214_, \uc8051golden_1.IRAM[59] [2]);
  buf _49157_ (_07215_, \uc8051golden_1.IRAM[59] [3]);
  buf _49158_ (_07217_, \uc8051golden_1.IRAM[59] [4]);
  buf _49159_ (_07218_, \uc8051golden_1.IRAM[59] [5]);
  buf _49160_ (_07219_, \uc8051golden_1.IRAM[59] [6]);
  buf _49161_ (_07220_, \uc8051golden_1.IRAM[59] [7]);
  buf _49162_ (_07221_, \uc8051golden_1.IRAM[60] [0]);
  buf _49163_ (_07222_, \uc8051golden_1.IRAM[60] [1]);
  buf _49164_ (_07223_, \uc8051golden_1.IRAM[60] [2]);
  buf _49165_ (_07224_, \uc8051golden_1.IRAM[60] [3]);
  buf _49166_ (_07225_, \uc8051golden_1.IRAM[60] [4]);
  buf _49167_ (_07226_, \uc8051golden_1.IRAM[60] [5]);
  buf _49168_ (_07227_, \uc8051golden_1.IRAM[60] [6]);
  buf _49169_ (_07228_, \uc8051golden_1.IRAM[60] [7]);
  buf _49170_ (_07229_, \uc8051golden_1.IRAM[61] [0]);
  buf _49171_ (_07230_, \uc8051golden_1.IRAM[61] [1]);
  buf _49172_ (_07231_, \uc8051golden_1.IRAM[61] [2]);
  buf _49173_ (_07232_, \uc8051golden_1.IRAM[61] [3]);
  buf _49174_ (_07233_, \uc8051golden_1.IRAM[61] [4]);
  buf _49175_ (_07234_, \uc8051golden_1.IRAM[61] [5]);
  buf _49176_ (_07235_, \uc8051golden_1.IRAM[61] [6]);
  buf _49177_ (_07236_, \uc8051golden_1.IRAM[61] [7]);
  buf _49178_ (_07237_, \uc8051golden_1.IRAM[62] [0]);
  buf _49179_ (_07238_, \uc8051golden_1.IRAM[62] [1]);
  buf _49180_ (_07239_, \uc8051golden_1.IRAM[62] [2]);
  buf _49181_ (_07240_, \uc8051golden_1.IRAM[62] [3]);
  buf _49182_ (_07241_, \uc8051golden_1.IRAM[62] [4]);
  buf _49183_ (_07242_, \uc8051golden_1.IRAM[62] [5]);
  buf _49184_ (_07243_, \uc8051golden_1.IRAM[62] [6]);
  buf _49185_ (_07244_, \uc8051golden_1.IRAM[62] [7]);
  buf _49186_ (_07245_, \uc8051golden_1.IRAM[63] [0]);
  buf _49187_ (_07246_, \uc8051golden_1.IRAM[63] [1]);
  buf _49188_ (_07247_, \uc8051golden_1.IRAM[63] [2]);
  buf _49189_ (_07248_, \uc8051golden_1.IRAM[63] [3]);
  buf _49190_ (_07249_, \uc8051golden_1.IRAM[63] [4]);
  buf _49191_ (_07251_, \uc8051golden_1.IRAM[63] [5]);
  buf _49192_ (_07252_, \uc8051golden_1.IRAM[63] [6]);
  buf _49193_ (_07253_, \uc8051golden_1.IRAM[63] [7]);
  buf _49194_ (_07254_, \uc8051golden_1.IRAM[64] [0]);
  buf _49195_ (_07255_, \uc8051golden_1.IRAM[64] [1]);
  buf _49196_ (_07256_, \uc8051golden_1.IRAM[64] [2]);
  buf _49197_ (_07257_, \uc8051golden_1.IRAM[64] [3]);
  buf _49198_ (_07258_, \uc8051golden_1.IRAM[64] [4]);
  buf _49199_ (_07259_, \uc8051golden_1.IRAM[64] [5]);
  buf _49200_ (_07260_, \uc8051golden_1.IRAM[64] [6]);
  buf _49201_ (_07261_, \uc8051golden_1.IRAM[64] [7]);
  buf _49202_ (_07262_, \uc8051golden_1.IRAM[65] [0]);
  buf _49203_ (_07263_, \uc8051golden_1.IRAM[65] [1]);
  buf _49204_ (_07264_, \uc8051golden_1.IRAM[65] [2]);
  buf _49205_ (_07265_, \uc8051golden_1.IRAM[65] [3]);
  buf _49206_ (_07266_, \uc8051golden_1.IRAM[65] [4]);
  buf _49207_ (_07267_, \uc8051golden_1.IRAM[65] [5]);
  buf _49208_ (_07268_, \uc8051golden_1.IRAM[65] [6]);
  buf _49209_ (_07269_, \uc8051golden_1.IRAM[65] [7]);
  buf _49210_ (_07270_, \uc8051golden_1.IRAM[66] [0]);
  buf _49211_ (_07271_, \uc8051golden_1.IRAM[66] [1]);
  buf _49212_ (_07272_, \uc8051golden_1.IRAM[66] [2]);
  buf _49213_ (_07273_, \uc8051golden_1.IRAM[66] [3]);
  buf _49214_ (_07274_, \uc8051golden_1.IRAM[66] [4]);
  buf _49215_ (_07275_, \uc8051golden_1.IRAM[66] [5]);
  buf _49216_ (_07276_, \uc8051golden_1.IRAM[66] [6]);
  buf _49217_ (_07277_, \uc8051golden_1.IRAM[66] [7]);
  buf _49218_ (_07278_, \uc8051golden_1.IRAM[67] [0]);
  buf _49219_ (_07279_, \uc8051golden_1.IRAM[67] [1]);
  buf _49220_ (_07280_, \uc8051golden_1.IRAM[67] [2]);
  buf _49221_ (_07281_, \uc8051golden_1.IRAM[67] [3]);
  buf _49222_ (_07282_, \uc8051golden_1.IRAM[67] [4]);
  buf _49223_ (_07284_, \uc8051golden_1.IRAM[67] [5]);
  buf _49224_ (_07285_, \uc8051golden_1.IRAM[67] [6]);
  buf _49225_ (_07286_, \uc8051golden_1.IRAM[67] [7]);
  buf _49226_ (_07287_, \uc8051golden_1.IRAM[68] [0]);
  buf _49227_ (_07288_, \uc8051golden_1.IRAM[68] [1]);
  buf _49228_ (_07289_, \uc8051golden_1.IRAM[68] [2]);
  buf _49229_ (_07290_, \uc8051golden_1.IRAM[68] [3]);
  buf _49230_ (_07291_, \uc8051golden_1.IRAM[68] [4]);
  buf _49231_ (_07292_, \uc8051golden_1.IRAM[68] [5]);
  buf _49232_ (_07293_, \uc8051golden_1.IRAM[68] [6]);
  buf _49233_ (_07294_, \uc8051golden_1.IRAM[68] [7]);
  buf _49234_ (_07295_, \uc8051golden_1.IRAM[69] [0]);
  buf _49235_ (_07296_, \uc8051golden_1.IRAM[69] [1]);
  buf _49236_ (_07297_, \uc8051golden_1.IRAM[69] [2]);
  buf _49237_ (_07298_, \uc8051golden_1.IRAM[69] [3]);
  buf _49238_ (_07299_, \uc8051golden_1.IRAM[69] [4]);
  buf _49239_ (_07300_, \uc8051golden_1.IRAM[69] [5]);
  buf _49240_ (_07301_, \uc8051golden_1.IRAM[69] [6]);
  buf _49241_ (_07302_, \uc8051golden_1.IRAM[69] [7]);
  buf _49242_ (_07303_, \uc8051golden_1.IRAM[70] [0]);
  buf _49243_ (_07304_, \uc8051golden_1.IRAM[70] [1]);
  buf _49244_ (_07305_, \uc8051golden_1.IRAM[70] [2]);
  buf _49245_ (_07306_, \uc8051golden_1.IRAM[70] [3]);
  buf _49246_ (_07307_, \uc8051golden_1.IRAM[70] [4]);
  buf _49247_ (_07308_, \uc8051golden_1.IRAM[70] [5]);
  buf _49248_ (_07309_, \uc8051golden_1.IRAM[70] [6]);
  buf _49249_ (_07310_, \uc8051golden_1.IRAM[70] [7]);
  buf _49250_ (_07311_, \uc8051golden_1.IRAM[71] [0]);
  buf _49251_ (_07312_, \uc8051golden_1.IRAM[71] [1]);
  buf _49252_ (_07313_, \uc8051golden_1.IRAM[71] [2]);
  buf _49253_ (_07314_, \uc8051golden_1.IRAM[71] [3]);
  buf _49254_ (_07315_, \uc8051golden_1.IRAM[71] [4]);
  buf _49255_ (_07316_, \uc8051golden_1.IRAM[71] [5]);
  buf _49256_ (_07318_, \uc8051golden_1.IRAM[71] [6]);
  buf _49257_ (_07319_, \uc8051golden_1.IRAM[71] [7]);
  buf _49258_ (_07320_, \uc8051golden_1.IRAM[72] [0]);
  buf _49259_ (_07321_, \uc8051golden_1.IRAM[72] [1]);
  buf _49260_ (_07322_, \uc8051golden_1.IRAM[72] [2]);
  buf _49261_ (_07323_, \uc8051golden_1.IRAM[72] [3]);
  buf _49262_ (_07324_, \uc8051golden_1.IRAM[72] [4]);
  buf _49263_ (_07325_, \uc8051golden_1.IRAM[72] [5]);
  buf _49264_ (_07326_, \uc8051golden_1.IRAM[72] [6]);
  buf _49265_ (_07327_, \uc8051golden_1.IRAM[72] [7]);
  buf _49266_ (_07328_, \uc8051golden_1.IRAM[73] [0]);
  buf _49267_ (_07329_, \uc8051golden_1.IRAM[73] [1]);
  buf _49268_ (_07330_, \uc8051golden_1.IRAM[73] [2]);
  buf _49269_ (_07331_, \uc8051golden_1.IRAM[73] [3]);
  buf _49270_ (_07332_, \uc8051golden_1.IRAM[73] [4]);
  buf _49271_ (_07333_, \uc8051golden_1.IRAM[73] [5]);
  buf _49272_ (_07334_, \uc8051golden_1.IRAM[73] [6]);
  buf _49273_ (_07335_, \uc8051golden_1.IRAM[73] [7]);
  buf _49274_ (_07336_, \uc8051golden_1.IRAM[74] [0]);
  buf _49275_ (_07337_, \uc8051golden_1.IRAM[74] [1]);
  buf _49276_ (_07338_, \uc8051golden_1.IRAM[74] [2]);
  buf _49277_ (_07339_, \uc8051golden_1.IRAM[74] [3]);
  buf _49278_ (_07340_, \uc8051golden_1.IRAM[74] [4]);
  buf _49279_ (_07341_, \uc8051golden_1.IRAM[74] [5]);
  buf _49280_ (_07342_, \uc8051golden_1.IRAM[74] [6]);
  buf _49281_ (_07343_, \uc8051golden_1.IRAM[74] [7]);
  buf _49282_ (_07344_, \uc8051golden_1.IRAM[75] [0]);
  buf _49283_ (_07345_, \uc8051golden_1.IRAM[75] [1]);
  buf _49284_ (_07346_, \uc8051golden_1.IRAM[75] [2]);
  buf _49285_ (_07347_, \uc8051golden_1.IRAM[75] [3]);
  buf _49286_ (_07348_, \uc8051golden_1.IRAM[75] [4]);
  buf _49287_ (_07349_, \uc8051golden_1.IRAM[75] [5]);
  buf _49288_ (_07350_, \uc8051golden_1.IRAM[75] [6]);
  buf _49289_ (_07351_, \uc8051golden_1.IRAM[75] [7]);
  buf _49290_ (_07353_, \uc8051golden_1.IRAM[76] [0]);
  buf _49291_ (_07354_, \uc8051golden_1.IRAM[76] [1]);
  buf _49292_ (_07355_, \uc8051golden_1.IRAM[76] [2]);
  buf _49293_ (_07356_, \uc8051golden_1.IRAM[76] [3]);
  buf _49294_ (_07357_, \uc8051golden_1.IRAM[76] [4]);
  buf _49295_ (_07358_, \uc8051golden_1.IRAM[76] [5]);
  buf _49296_ (_07359_, \uc8051golden_1.IRAM[76] [6]);
  buf _49297_ (_07360_, \uc8051golden_1.IRAM[76] [7]);
  buf _49298_ (_07361_, \uc8051golden_1.IRAM[77] [0]);
  buf _49299_ (_07362_, \uc8051golden_1.IRAM[77] [1]);
  buf _49300_ (_07363_, \uc8051golden_1.IRAM[77] [2]);
  buf _49301_ (_07364_, \uc8051golden_1.IRAM[77] [3]);
  buf _49302_ (_07365_, \uc8051golden_1.IRAM[77] [4]);
  buf _49303_ (_07366_, \uc8051golden_1.IRAM[77] [5]);
  buf _49304_ (_07367_, \uc8051golden_1.IRAM[77] [6]);
  buf _49305_ (_07368_, \uc8051golden_1.IRAM[77] [7]);
  buf _49306_ (_07369_, \uc8051golden_1.IRAM[78] [0]);
  buf _49307_ (_07370_, \uc8051golden_1.IRAM[78] [1]);
  buf _49308_ (_07371_, \uc8051golden_1.IRAM[78] [2]);
  buf _49309_ (_07372_, \uc8051golden_1.IRAM[78] [3]);
  buf _49310_ (_07373_, \uc8051golden_1.IRAM[78] [4]);
  buf _49311_ (_07374_, \uc8051golden_1.IRAM[78] [5]);
  buf _49312_ (_07375_, \uc8051golden_1.IRAM[78] [6]);
  buf _49313_ (_07376_, \uc8051golden_1.IRAM[78] [7]);
  buf _49314_ (_07377_, \uc8051golden_1.IRAM[79] [0]);
  buf _49315_ (_07378_, \uc8051golden_1.IRAM[79] [1]);
  buf _49316_ (_07379_, \uc8051golden_1.IRAM[79] [2]);
  buf _49317_ (_07380_, \uc8051golden_1.IRAM[79] [3]);
  buf _49318_ (_07381_, \uc8051golden_1.IRAM[79] [4]);
  buf _49319_ (_07382_, \uc8051golden_1.IRAM[79] [5]);
  buf _49320_ (_07383_, \uc8051golden_1.IRAM[79] [6]);
  buf _49321_ (_07384_, \uc8051golden_1.IRAM[79] [7]);
  buf _49322_ (_07385_, \uc8051golden_1.IRAM[80] [0]);
  buf _49323_ (_07387_, \uc8051golden_1.IRAM[80] [1]);
  buf _49324_ (_07388_, \uc8051golden_1.IRAM[80] [2]);
  buf _49325_ (_07389_, \uc8051golden_1.IRAM[80] [3]);
  buf _49326_ (_07390_, \uc8051golden_1.IRAM[80] [4]);
  buf _49327_ (_07391_, \uc8051golden_1.IRAM[80] [5]);
  buf _49328_ (_07392_, \uc8051golden_1.IRAM[80] [6]);
  buf _49329_ (_07393_, \uc8051golden_1.IRAM[80] [7]);
  buf _49330_ (_07394_, \uc8051golden_1.IRAM[81] [0]);
  buf _49331_ (_07395_, \uc8051golden_1.IRAM[81] [1]);
  buf _49332_ (_07396_, \uc8051golden_1.IRAM[81] [2]);
  buf _49333_ (_07397_, \uc8051golden_1.IRAM[81] [3]);
  buf _49334_ (_07398_, \uc8051golden_1.IRAM[81] [4]);
  buf _49335_ (_07399_, \uc8051golden_1.IRAM[81] [5]);
  buf _49336_ (_07400_, \uc8051golden_1.IRAM[81] [6]);
  buf _49337_ (_07401_, \uc8051golden_1.IRAM[81] [7]);
  buf _49338_ (_07402_, \uc8051golden_1.IRAM[82] [0]);
  buf _49339_ (_07403_, \uc8051golden_1.IRAM[82] [1]);
  buf _49340_ (_07404_, \uc8051golden_1.IRAM[82] [2]);
  buf _49341_ (_07405_, \uc8051golden_1.IRAM[82] [3]);
  buf _49342_ (_07406_, \uc8051golden_1.IRAM[82] [4]);
  buf _49343_ (_07407_, \uc8051golden_1.IRAM[82] [5]);
  buf _49344_ (_07408_, \uc8051golden_1.IRAM[82] [6]);
  buf _49345_ (_07409_, \uc8051golden_1.IRAM[82] [7]);
  buf _49346_ (_07410_, \uc8051golden_1.IRAM[83] [0]);
  buf _49347_ (_07411_, \uc8051golden_1.IRAM[83] [1]);
  buf _49348_ (_07412_, \uc8051golden_1.IRAM[83] [2]);
  buf _49349_ (_07413_, \uc8051golden_1.IRAM[83] [3]);
  buf _49350_ (_07414_, \uc8051golden_1.IRAM[83] [4]);
  buf _49351_ (_07415_, \uc8051golden_1.IRAM[83] [5]);
  buf _49352_ (_07416_, \uc8051golden_1.IRAM[83] [6]);
  buf _49353_ (_07417_, \uc8051golden_1.IRAM[83] [7]);
  buf _49354_ (_07418_, \uc8051golden_1.IRAM[84] [0]);
  buf _49355_ (_07419_, \uc8051golden_1.IRAM[84] [1]);
  buf _49356_ (_07421_, \uc8051golden_1.IRAM[84] [2]);
  buf _49357_ (_07422_, \uc8051golden_1.IRAM[84] [3]);
  buf _49358_ (_07423_, \uc8051golden_1.IRAM[84] [4]);
  buf _49359_ (_07424_, \uc8051golden_1.IRAM[84] [5]);
  buf _49360_ (_07425_, \uc8051golden_1.IRAM[84] [6]);
  buf _49361_ (_07426_, \uc8051golden_1.IRAM[84] [7]);
  buf _49362_ (_07427_, \uc8051golden_1.IRAM[85] [0]);
  buf _49363_ (_07428_, \uc8051golden_1.IRAM[85] [1]);
  buf _49364_ (_07429_, \uc8051golden_1.IRAM[85] [2]);
  buf _49365_ (_07430_, \uc8051golden_1.IRAM[85] [3]);
  buf _49366_ (_07431_, \uc8051golden_1.IRAM[85] [4]);
  buf _49367_ (_07432_, \uc8051golden_1.IRAM[85] [5]);
  buf _49368_ (_07433_, \uc8051golden_1.IRAM[85] [6]);
  buf _49369_ (_07434_, \uc8051golden_1.IRAM[85] [7]);
  buf _49370_ (_07435_, \uc8051golden_1.IRAM[86] [0]);
  buf _49371_ (_07436_, \uc8051golden_1.IRAM[86] [1]);
  buf _49372_ (_07437_, \uc8051golden_1.IRAM[86] [2]);
  buf _49373_ (_07438_, \uc8051golden_1.IRAM[86] [3]);
  buf _49374_ (_07439_, \uc8051golden_1.IRAM[86] [4]);
  buf _49375_ (_07440_, \uc8051golden_1.IRAM[86] [5]);
  buf _49376_ (_07441_, \uc8051golden_1.IRAM[86] [6]);
  buf _49377_ (_07442_, \uc8051golden_1.IRAM[86] [7]);
  buf _49378_ (_07443_, \uc8051golden_1.IRAM[87] [0]);
  buf _49379_ (_07444_, \uc8051golden_1.IRAM[87] [1]);
  buf _49380_ (_07445_, \uc8051golden_1.IRAM[87] [2]);
  buf _49381_ (_07446_, \uc8051golden_1.IRAM[87] [3]);
  buf _49382_ (_07447_, \uc8051golden_1.IRAM[87] [4]);
  buf _49383_ (_07448_, \uc8051golden_1.IRAM[87] [5]);
  buf _49384_ (_07449_, \uc8051golden_1.IRAM[87] [6]);
  buf _49385_ (_07450_, \uc8051golden_1.IRAM[87] [7]);
  buf _49386_ (_07451_, \uc8051golden_1.IRAM[88] [0]);
  buf _49387_ (_07452_, \uc8051golden_1.IRAM[88] [1]);
  buf _49388_ (_07453_, \uc8051golden_1.IRAM[88] [2]);
  buf _49389_ (_07455_, \uc8051golden_1.IRAM[88] [3]);
  buf _49390_ (_07456_, \uc8051golden_1.IRAM[88] [4]);
  buf _49391_ (_07457_, \uc8051golden_1.IRAM[88] [5]);
  buf _49392_ (_07458_, \uc8051golden_1.IRAM[88] [6]);
  buf _49393_ (_07459_, \uc8051golden_1.IRAM[88] [7]);
  buf _49394_ (_07460_, \uc8051golden_1.IRAM[89] [0]);
  buf _49395_ (_07461_, \uc8051golden_1.IRAM[89] [1]);
  buf _49396_ (_07462_, \uc8051golden_1.IRAM[89] [2]);
  buf _49397_ (_07463_, \uc8051golden_1.IRAM[89] [3]);
  buf _49398_ (_07464_, \uc8051golden_1.IRAM[89] [4]);
  buf _49399_ (_07465_, \uc8051golden_1.IRAM[89] [5]);
  buf _49400_ (_07466_, \uc8051golden_1.IRAM[89] [6]);
  buf _49401_ (_07467_, \uc8051golden_1.IRAM[89] [7]);
  buf _49402_ (_07468_, \uc8051golden_1.IRAM[90] [0]);
  buf _49403_ (_07469_, \uc8051golden_1.IRAM[90] [1]);
  buf _49404_ (_07470_, \uc8051golden_1.IRAM[90] [2]);
  buf _49405_ (_07471_, \uc8051golden_1.IRAM[90] [3]);
  buf _49406_ (_07472_, \uc8051golden_1.IRAM[90] [4]);
  buf _49407_ (_07473_, \uc8051golden_1.IRAM[90] [5]);
  buf _49408_ (_07474_, \uc8051golden_1.IRAM[90] [6]);
  buf _49409_ (_07475_, \uc8051golden_1.IRAM[90] [7]);
  buf _49410_ (_07476_, \uc8051golden_1.IRAM[91] [0]);
  buf _49411_ (_07477_, \uc8051golden_1.IRAM[91] [1]);
  buf _49412_ (_07478_, \uc8051golden_1.IRAM[91] [2]);
  buf _49413_ (_07479_, \uc8051golden_1.IRAM[91] [3]);
  buf _49414_ (_07480_, \uc8051golden_1.IRAM[91] [4]);
  buf _49415_ (_07481_, \uc8051golden_1.IRAM[91] [5]);
  buf _49416_ (_07482_, \uc8051golden_1.IRAM[91] [6]);
  buf _49417_ (_07483_, \uc8051golden_1.IRAM[91] [7]);
  buf _49418_ (_07484_, \uc8051golden_1.IRAM[92] [0]);
  buf _49419_ (_07485_, \uc8051golden_1.IRAM[92] [1]);
  buf _49420_ (_07486_, \uc8051golden_1.IRAM[92] [2]);
  buf _49421_ (_07487_, \uc8051golden_1.IRAM[92] [3]);
  buf _49422_ (_07488_, \uc8051golden_1.IRAM[92] [4]);
  buf _49423_ (_07490_, \uc8051golden_1.IRAM[92] [5]);
  buf _49424_ (_07491_, \uc8051golden_1.IRAM[92] [6]);
  buf _49425_ (_07492_, \uc8051golden_1.IRAM[92] [7]);
  buf _49426_ (_07493_, \uc8051golden_1.IRAM[93] [0]);
  buf _49427_ (_07494_, \uc8051golden_1.IRAM[93] [1]);
  buf _49428_ (_07495_, \uc8051golden_1.IRAM[93] [2]);
  buf _49429_ (_07496_, \uc8051golden_1.IRAM[93] [3]);
  buf _49430_ (_07497_, \uc8051golden_1.IRAM[93] [4]);
  buf _49431_ (_07498_, \uc8051golden_1.IRAM[93] [5]);
  buf _49432_ (_07499_, \uc8051golden_1.IRAM[93] [6]);
  buf _49433_ (_07500_, \uc8051golden_1.IRAM[93] [7]);
  buf _49434_ (_07501_, \uc8051golden_1.IRAM[94] [0]);
  buf _49435_ (_07502_, \uc8051golden_1.IRAM[94] [1]);
  buf _49436_ (_07503_, \uc8051golden_1.IRAM[94] [2]);
  buf _49437_ (_07504_, \uc8051golden_1.IRAM[94] [3]);
  buf _49438_ (_07505_, \uc8051golden_1.IRAM[94] [4]);
  buf _49439_ (_07506_, \uc8051golden_1.IRAM[94] [5]);
  buf _49440_ (_07507_, \uc8051golden_1.IRAM[94] [6]);
  buf _49441_ (_07508_, \uc8051golden_1.IRAM[94] [7]);
  buf _49442_ (_07509_, \uc8051golden_1.IRAM[95] [0]);
  buf _49443_ (_07510_, \uc8051golden_1.IRAM[95] [1]);
  buf _49444_ (_07511_, \uc8051golden_1.IRAM[95] [2]);
  buf _49445_ (_07512_, \uc8051golden_1.IRAM[95] [3]);
  buf _49446_ (_07513_, \uc8051golden_1.IRAM[95] [4]);
  buf _49447_ (_07514_, \uc8051golden_1.IRAM[95] [5]);
  buf _49448_ (_07515_, \uc8051golden_1.IRAM[95] [6]);
  buf _49449_ (_07516_, \uc8051golden_1.IRAM[95] [7]);
  buf _49450_ (_07517_, \uc8051golden_1.IRAM[96] [0]);
  buf _49451_ (_07518_, \uc8051golden_1.IRAM[96] [1]);
  buf _49452_ (_07519_, \uc8051golden_1.IRAM[96] [2]);
  buf _49453_ (_07520_, \uc8051golden_1.IRAM[96] [3]);
  buf _49454_ (_07521_, \uc8051golden_1.IRAM[96] [4]);
  buf _49455_ (_07522_, \uc8051golden_1.IRAM[96] [5]);
  buf _49456_ (_07524_, \uc8051golden_1.IRAM[96] [6]);
  buf _49457_ (_07525_, \uc8051golden_1.IRAM[96] [7]);
  buf _49458_ (_07526_, \uc8051golden_1.IRAM[97] [0]);
  buf _49459_ (_07527_, \uc8051golden_1.IRAM[97] [1]);
  buf _49460_ (_07528_, \uc8051golden_1.IRAM[97] [2]);
  buf _49461_ (_07529_, \uc8051golden_1.IRAM[97] [3]);
  buf _49462_ (_07530_, \uc8051golden_1.IRAM[97] [4]);
  buf _49463_ (_07531_, \uc8051golden_1.IRAM[97] [5]);
  buf _49464_ (_07532_, \uc8051golden_1.IRAM[97] [6]);
  buf _49465_ (_07533_, \uc8051golden_1.IRAM[97] [7]);
  buf _49466_ (_07534_, \uc8051golden_1.IRAM[98] [0]);
  buf _49467_ (_07535_, \uc8051golden_1.IRAM[98] [1]);
  buf _49468_ (_07536_, \uc8051golden_1.IRAM[98] [2]);
  buf _49469_ (_07537_, \uc8051golden_1.IRAM[98] [3]);
  buf _49470_ (_07538_, \uc8051golden_1.IRAM[98] [4]);
  buf _49471_ (_07539_, \uc8051golden_1.IRAM[98] [5]);
  buf _49472_ (_07540_, \uc8051golden_1.IRAM[98] [6]);
  buf _49473_ (_07541_, \uc8051golden_1.IRAM[98] [7]);
  buf _49474_ (_07542_, \uc8051golden_1.IRAM[99] [0]);
  buf _49475_ (_07543_, \uc8051golden_1.IRAM[99] [1]);
  buf _49476_ (_07544_, \uc8051golden_1.IRAM[99] [2]);
  buf _49477_ (_07545_, \uc8051golden_1.IRAM[99] [3]);
  buf _49478_ (_07546_, \uc8051golden_1.IRAM[99] [4]);
  buf _49479_ (_07547_, \uc8051golden_1.IRAM[99] [5]);
  buf _49480_ (_07548_, \uc8051golden_1.IRAM[99] [6]);
  buf _49481_ (_07549_, \uc8051golden_1.IRAM[99] [7]);
  buf _49482_ (_07550_, \uc8051golden_1.IRAM[100] [0]);
  buf _49483_ (_07551_, \uc8051golden_1.IRAM[100] [1]);
  buf _49484_ (_07552_, \uc8051golden_1.IRAM[100] [2]);
  buf _49485_ (_07553_, \uc8051golden_1.IRAM[100] [3]);
  buf _49486_ (_07554_, \uc8051golden_1.IRAM[100] [4]);
  buf _49487_ (_07555_, \uc8051golden_1.IRAM[100] [5]);
  buf _49488_ (_07556_, \uc8051golden_1.IRAM[100] [6]);
  buf _49489_ (_07558_, \uc8051golden_1.IRAM[100] [7]);
  buf _49490_ (_07559_, \uc8051golden_1.IRAM[101] [0]);
  buf _49491_ (_07560_, \uc8051golden_1.IRAM[101] [1]);
  buf _49492_ (_07561_, \uc8051golden_1.IRAM[101] [2]);
  buf _49493_ (_07562_, \uc8051golden_1.IRAM[101] [3]);
  buf _49494_ (_07563_, \uc8051golden_1.IRAM[101] [4]);
  buf _49495_ (_07564_, \uc8051golden_1.IRAM[101] [5]);
  buf _49496_ (_07565_, \uc8051golden_1.IRAM[101] [6]);
  buf _49497_ (_07566_, \uc8051golden_1.IRAM[101] [7]);
  buf _49498_ (_07567_, \uc8051golden_1.IRAM[102] [0]);
  buf _49499_ (_07568_, \uc8051golden_1.IRAM[102] [1]);
  buf _49500_ (_07569_, \uc8051golden_1.IRAM[102] [2]);
  buf _49501_ (_07570_, \uc8051golden_1.IRAM[102] [3]);
  buf _49502_ (_07571_, \uc8051golden_1.IRAM[102] [4]);
  buf _49503_ (_07572_, \uc8051golden_1.IRAM[102] [5]);
  buf _49504_ (_07573_, \uc8051golden_1.IRAM[102] [6]);
  buf _49505_ (_07574_, \uc8051golden_1.IRAM[102] [7]);
  buf _49506_ (_07575_, \uc8051golden_1.IRAM[103] [0]);
  buf _49507_ (_07576_, \uc8051golden_1.IRAM[103] [1]);
  buf _49508_ (_07577_, \uc8051golden_1.IRAM[103] [2]);
  buf _49509_ (_07578_, \uc8051golden_1.IRAM[103] [3]);
  buf _49510_ (_07579_, \uc8051golden_1.IRAM[103] [4]);
  buf _49511_ (_07580_, \uc8051golden_1.IRAM[103] [5]);
  buf _49512_ (_07581_, \uc8051golden_1.IRAM[103] [6]);
  buf _49513_ (_07582_, \uc8051golden_1.IRAM[103] [7]);
  buf _49514_ (_07583_, \uc8051golden_1.IRAM[104] [0]);
  buf _49515_ (_07584_, \uc8051golden_1.IRAM[104] [1]);
  buf _49516_ (_07585_, \uc8051golden_1.IRAM[104] [2]);
  buf _49517_ (_07586_, \uc8051golden_1.IRAM[104] [3]);
  buf _49518_ (_07587_, \uc8051golden_1.IRAM[104] [4]);
  buf _49519_ (_07588_, \uc8051golden_1.IRAM[104] [5]);
  buf _49520_ (_07589_, \uc8051golden_1.IRAM[104] [6]);
  buf _49521_ (_07590_, \uc8051golden_1.IRAM[104] [7]);
  buf _49522_ (_07592_, \uc8051golden_1.IRAM[105] [0]);
  buf _49523_ (_07593_, \uc8051golden_1.IRAM[105] [1]);
  buf _49524_ (_07594_, \uc8051golden_1.IRAM[105] [2]);
  buf _49525_ (_07595_, \uc8051golden_1.IRAM[105] [3]);
  buf _49526_ (_07596_, \uc8051golden_1.IRAM[105] [4]);
  buf _49527_ (_07597_, \uc8051golden_1.IRAM[105] [5]);
  buf _49528_ (_07598_, \uc8051golden_1.IRAM[105] [6]);
  buf _49529_ (_07599_, \uc8051golden_1.IRAM[105] [7]);
  buf _49530_ (_07600_, \uc8051golden_1.IRAM[106] [0]);
  buf _49531_ (_07601_, \uc8051golden_1.IRAM[106] [1]);
  buf _49532_ (_07602_, \uc8051golden_1.IRAM[106] [2]);
  buf _49533_ (_07603_, \uc8051golden_1.IRAM[106] [3]);
  buf _49534_ (_07604_, \uc8051golden_1.IRAM[106] [4]);
  buf _49535_ (_07605_, \uc8051golden_1.IRAM[106] [5]);
  buf _49536_ (_07606_, \uc8051golden_1.IRAM[106] [6]);
  buf _49537_ (_07607_, \uc8051golden_1.IRAM[106] [7]);
  buf _49538_ (_07608_, \uc8051golden_1.IRAM[107] [0]);
  buf _49539_ (_07609_, \uc8051golden_1.IRAM[107] [1]);
  buf _49540_ (_07610_, \uc8051golden_1.IRAM[107] [2]);
  buf _49541_ (_07611_, \uc8051golden_1.IRAM[107] [3]);
  buf _49542_ (_07612_, \uc8051golden_1.IRAM[107] [4]);
  buf _49543_ (_07613_, \uc8051golden_1.IRAM[107] [5]);
  buf _49544_ (_07614_, \uc8051golden_1.IRAM[107] [6]);
  buf _49545_ (_07615_, \uc8051golden_1.IRAM[107] [7]);
  buf _49546_ (_07616_, \uc8051golden_1.IRAM[108] [0]);
  buf _49547_ (_07617_, \uc8051golden_1.IRAM[108] [1]);
  buf _49548_ (_07618_, \uc8051golden_1.IRAM[108] [2]);
  buf _49549_ (_07619_, \uc8051golden_1.IRAM[108] [3]);
  buf _49550_ (_07620_, \uc8051golden_1.IRAM[108] [4]);
  buf _49551_ (_07621_, \uc8051golden_1.IRAM[108] [5]);
  buf _49552_ (_07622_, \uc8051golden_1.IRAM[108] [6]);
  buf _49553_ (_07623_, \uc8051golden_1.IRAM[108] [7]);
  buf _49554_ (_07624_, \uc8051golden_1.IRAM[109] [0]);
  buf _49555_ (_07625_, \uc8051golden_1.IRAM[109] [1]);
  buf _49556_ (_07627_, \uc8051golden_1.IRAM[109] [2]);
  buf _49557_ (_07628_, \uc8051golden_1.IRAM[109] [3]);
  buf _49558_ (_07629_, \uc8051golden_1.IRAM[109] [4]);
  buf _49559_ (_07630_, \uc8051golden_1.IRAM[109] [5]);
  buf _49560_ (_07631_, \uc8051golden_1.IRAM[109] [6]);
  buf _49561_ (_07632_, \uc8051golden_1.IRAM[109] [7]);
  buf _49562_ (_07633_, \uc8051golden_1.IRAM[110] [0]);
  buf _49563_ (_07634_, \uc8051golden_1.IRAM[110] [1]);
  buf _49564_ (_07635_, \uc8051golden_1.IRAM[110] [2]);
  buf _49565_ (_07636_, \uc8051golden_1.IRAM[110] [3]);
  buf _49566_ (_07637_, \uc8051golden_1.IRAM[110] [4]);
  buf _49567_ (_07638_, \uc8051golden_1.IRAM[110] [5]);
  buf _49568_ (_07639_, \uc8051golden_1.IRAM[110] [6]);
  buf _49569_ (_07640_, \uc8051golden_1.IRAM[110] [7]);
  buf _49570_ (_07641_, \uc8051golden_1.IRAM[111] [0]);
  buf _49571_ (_07642_, \uc8051golden_1.IRAM[111] [1]);
  buf _49572_ (_07643_, \uc8051golden_1.IRAM[111] [2]);
  buf _49573_ (_07644_, \uc8051golden_1.IRAM[111] [3]);
  buf _49574_ (_07645_, \uc8051golden_1.IRAM[111] [4]);
  buf _49575_ (_07646_, \uc8051golden_1.IRAM[111] [5]);
  buf _49576_ (_07647_, \uc8051golden_1.IRAM[111] [6]);
  buf _49577_ (_07648_, \uc8051golden_1.IRAM[111] [7]);
  buf _49578_ (_07649_, \uc8051golden_1.IRAM[112] [0]);
  buf _49579_ (_07650_, \uc8051golden_1.IRAM[112] [1]);
  buf _49580_ (_07651_, \uc8051golden_1.IRAM[112] [2]);
  buf _49581_ (_07652_, \uc8051golden_1.IRAM[112] [3]);
  buf _49582_ (_07653_, \uc8051golden_1.IRAM[112] [4]);
  buf _49583_ (_07654_, \uc8051golden_1.IRAM[112] [5]);
  buf _49584_ (_07655_, \uc8051golden_1.IRAM[112] [6]);
  buf _49585_ (_07656_, \uc8051golden_1.IRAM[112] [7]);
  buf _49586_ (_07657_, \uc8051golden_1.IRAM[113] [0]);
  buf _49587_ (_07658_, \uc8051golden_1.IRAM[113] [1]);
  buf _49588_ (_07659_, \uc8051golden_1.IRAM[113] [2]);
  buf _49589_ (_07661_, \uc8051golden_1.IRAM[113] [3]);
  buf _49590_ (_07662_, \uc8051golden_1.IRAM[113] [4]);
  buf _49591_ (_07663_, \uc8051golden_1.IRAM[113] [5]);
  buf _49592_ (_07664_, \uc8051golden_1.IRAM[113] [6]);
  buf _49593_ (_07665_, \uc8051golden_1.IRAM[113] [7]);
  buf _49594_ (_07666_, \uc8051golden_1.IRAM[114] [0]);
  buf _49595_ (_07667_, \uc8051golden_1.IRAM[114] [1]);
  buf _49596_ (_07668_, \uc8051golden_1.IRAM[114] [2]);
  buf _49597_ (_07669_, \uc8051golden_1.IRAM[114] [3]);
  buf _49598_ (_07670_, \uc8051golden_1.IRAM[114] [4]);
  buf _49599_ (_07671_, \uc8051golden_1.IRAM[114] [5]);
  buf _49600_ (_07672_, \uc8051golden_1.IRAM[114] [6]);
  buf _49601_ (_07673_, \uc8051golden_1.IRAM[114] [7]);
  buf _49602_ (_07674_, \uc8051golden_1.IRAM[115] [0]);
  buf _49603_ (_07675_, \uc8051golden_1.IRAM[115] [1]);
  buf _49604_ (_07676_, \uc8051golden_1.IRAM[115] [2]);
  buf _49605_ (_07677_, \uc8051golden_1.IRAM[115] [3]);
  buf _49606_ (_07678_, \uc8051golden_1.IRAM[115] [4]);
  buf _49607_ (_07679_, \uc8051golden_1.IRAM[115] [5]);
  buf _49608_ (_07680_, \uc8051golden_1.IRAM[115] [6]);
  buf _49609_ (_07681_, \uc8051golden_1.IRAM[115] [7]);
  buf _49610_ (_07682_, \uc8051golden_1.IRAM[116] [0]);
  buf _49611_ (_07683_, \uc8051golden_1.IRAM[116] [1]);
  buf _49612_ (_07684_, \uc8051golden_1.IRAM[116] [2]);
  buf _49613_ (_07685_, \uc8051golden_1.IRAM[116] [3]);
  buf _49614_ (_07686_, \uc8051golden_1.IRAM[116] [4]);
  buf _49615_ (_07687_, \uc8051golden_1.IRAM[116] [5]);
  buf _49616_ (_07688_, \uc8051golden_1.IRAM[116] [6]);
  buf _49617_ (_07689_, \uc8051golden_1.IRAM[116] [7]);
  buf _49618_ (_07690_, \uc8051golden_1.IRAM[117] [0]);
  buf _49619_ (_07691_, \uc8051golden_1.IRAM[117] [1]);
  buf _49620_ (_07692_, \uc8051golden_1.IRAM[117] [2]);
  buf _49621_ (_07693_, \uc8051golden_1.IRAM[117] [3]);
  buf _49622_ (_07695_, \uc8051golden_1.IRAM[117] [4]);
  buf _49623_ (_07696_, \uc8051golden_1.IRAM[117] [5]);
  buf _49624_ (_07697_, \uc8051golden_1.IRAM[117] [6]);
  buf _49625_ (_07698_, \uc8051golden_1.IRAM[117] [7]);
  buf _49626_ (_07699_, \uc8051golden_1.IRAM[118] [0]);
  buf _49627_ (_07700_, \uc8051golden_1.IRAM[118] [1]);
  buf _49628_ (_07701_, \uc8051golden_1.IRAM[118] [2]);
  buf _49629_ (_07702_, \uc8051golden_1.IRAM[118] [3]);
  buf _49630_ (_07703_, \uc8051golden_1.IRAM[118] [4]);
  buf _49631_ (_07704_, \uc8051golden_1.IRAM[118] [5]);
  buf _49632_ (_07705_, \uc8051golden_1.IRAM[118] [6]);
  buf _49633_ (_07706_, \uc8051golden_1.IRAM[118] [7]);
  buf _49634_ (_07707_, \uc8051golden_1.IRAM[119] [0]);
  buf _49635_ (_07708_, \uc8051golden_1.IRAM[119] [1]);
  buf _49636_ (_07709_, \uc8051golden_1.IRAM[119] [2]);
  buf _49637_ (_07710_, \uc8051golden_1.IRAM[119] [3]);
  buf _49638_ (_07711_, \uc8051golden_1.IRAM[119] [4]);
  buf _49639_ (_07712_, \uc8051golden_1.IRAM[119] [5]);
  buf _49640_ (_07713_, \uc8051golden_1.IRAM[119] [6]);
  buf _49641_ (_07714_, \uc8051golden_1.IRAM[119] [7]);
  buf _49642_ (_07715_, \uc8051golden_1.IRAM[120] [0]);
  buf _49643_ (_07716_, \uc8051golden_1.IRAM[120] [1]);
  buf _49644_ (_07717_, \uc8051golden_1.IRAM[120] [2]);
  buf _49645_ (_07718_, \uc8051golden_1.IRAM[120] [3]);
  buf _49646_ (_07719_, \uc8051golden_1.IRAM[120] [4]);
  buf _49647_ (_07720_, \uc8051golden_1.IRAM[120] [5]);
  buf _49648_ (_07721_, \uc8051golden_1.IRAM[120] [6]);
  buf _49649_ (_07722_, \uc8051golden_1.IRAM[120] [7]);
  buf _49650_ (_07723_, \uc8051golden_1.IRAM[121] [0]);
  buf _49651_ (_07724_, \uc8051golden_1.IRAM[121] [1]);
  buf _49652_ (_07725_, \uc8051golden_1.IRAM[121] [2]);
  buf _49653_ (_07726_, \uc8051golden_1.IRAM[121] [3]);
  buf _49654_ (_07727_, \uc8051golden_1.IRAM[121] [4]);
  buf _49655_ (_07729_, \uc8051golden_1.IRAM[121] [5]);
  buf _49656_ (_07730_, \uc8051golden_1.IRAM[121] [6]);
  buf _49657_ (_07731_, \uc8051golden_1.IRAM[121] [7]);
  buf _49658_ (_07732_, \uc8051golden_1.IRAM[122] [0]);
  buf _49659_ (_07733_, \uc8051golden_1.IRAM[122] [1]);
  buf _49660_ (_07734_, \uc8051golden_1.IRAM[122] [2]);
  buf _49661_ (_07735_, \uc8051golden_1.IRAM[122] [3]);
  buf _49662_ (_07736_, \uc8051golden_1.IRAM[122] [4]);
  buf _49663_ (_07737_, \uc8051golden_1.IRAM[122] [5]);
  buf _49664_ (_07738_, \uc8051golden_1.IRAM[122] [6]);
  buf _49665_ (_07739_, \uc8051golden_1.IRAM[122] [7]);
  buf _49666_ (_07740_, \uc8051golden_1.IRAM[123] [0]);
  buf _49667_ (_07741_, \uc8051golden_1.IRAM[123] [1]);
  buf _49668_ (_07742_, \uc8051golden_1.IRAM[123] [2]);
  buf _49669_ (_07743_, \uc8051golden_1.IRAM[123] [3]);
  buf _49670_ (_07744_, \uc8051golden_1.IRAM[123] [4]);
  buf _49671_ (_07745_, \uc8051golden_1.IRAM[123] [5]);
  buf _49672_ (_07746_, \uc8051golden_1.IRAM[123] [6]);
  buf _49673_ (_07747_, \uc8051golden_1.IRAM[123] [7]);
  buf _49674_ (_07748_, \uc8051golden_1.IRAM[124] [0]);
  buf _49675_ (_07749_, \uc8051golden_1.IRAM[124] [1]);
  buf _49676_ (_07750_, \uc8051golden_1.IRAM[124] [2]);
  buf _49677_ (_07751_, \uc8051golden_1.IRAM[124] [3]);
  buf _49678_ (_07752_, \uc8051golden_1.IRAM[124] [4]);
  buf _49679_ (_07753_, \uc8051golden_1.IRAM[124] [5]);
  buf _49680_ (_07754_, \uc8051golden_1.IRAM[124] [6]);
  buf _49681_ (_07755_, \uc8051golden_1.IRAM[124] [7]);
  buf _49682_ (_07756_, \uc8051golden_1.IRAM[125] [0]);
  buf _49683_ (_07757_, \uc8051golden_1.IRAM[125] [1]);
  buf _49684_ (_07758_, \uc8051golden_1.IRAM[125] [2]);
  buf _49685_ (_07759_, \uc8051golden_1.IRAM[125] [3]);
  buf _49686_ (_07760_, \uc8051golden_1.IRAM[125] [4]);
  buf _49687_ (_07761_, \uc8051golden_1.IRAM[125] [5]);
  buf _49688_ (_07762_, \uc8051golden_1.IRAM[125] [6]);
  buf _49689_ (_07764_, \uc8051golden_1.IRAM[125] [7]);
  buf _49690_ (_07765_, \uc8051golden_1.IRAM[126] [0]);
  buf _49691_ (_07766_, \uc8051golden_1.IRAM[126] [1]);
  buf _49692_ (_07767_, \uc8051golden_1.IRAM[126] [2]);
  buf _49693_ (_07768_, \uc8051golden_1.IRAM[126] [3]);
  buf _49694_ (_07769_, \uc8051golden_1.IRAM[126] [4]);
  buf _49695_ (_07770_, \uc8051golden_1.IRAM[126] [5]);
  buf _49696_ (_07771_, \uc8051golden_1.IRAM[126] [6]);
  buf _49697_ (_07772_, \uc8051golden_1.IRAM[126] [7]);
  buf _49698_ (_07773_, \uc8051golden_1.IRAM[127] [0]);
  buf _49699_ (_07774_, \uc8051golden_1.IRAM[127] [1]);
  buf _49700_ (_07775_, \uc8051golden_1.IRAM[127] [2]);
  buf _49701_ (_07776_, \uc8051golden_1.IRAM[127] [3]);
  buf _49702_ (_07777_, \uc8051golden_1.IRAM[127] [4]);
  buf _49703_ (_07778_, \uc8051golden_1.IRAM[127] [5]);
  buf _49704_ (_07779_, \uc8051golden_1.IRAM[127] [6]);
  buf _49705_ (_07780_, \uc8051golden_1.IRAM[127] [7]);
  buf _49706_ (_07781_, \uc8051golden_1.IRAM[128] [0]);
  buf _49707_ (_07782_, \uc8051golden_1.IRAM[128] [1]);
  buf _49708_ (_07783_, \uc8051golden_1.IRAM[128] [2]);
  buf _49709_ (_07784_, \uc8051golden_1.IRAM[128] [3]);
  buf _49710_ (_07785_, \uc8051golden_1.IRAM[128] [4]);
  buf _49711_ (_07786_, \uc8051golden_1.IRAM[128] [5]);
  buf _49712_ (_07787_, \uc8051golden_1.IRAM[128] [6]);
  buf _49713_ (_07788_, \uc8051golden_1.IRAM[128] [7]);
  buf _49714_ (_07789_, \uc8051golden_1.IRAM[129] [0]);
  buf _49715_ (_07790_, \uc8051golden_1.IRAM[129] [1]);
  buf _49716_ (_07791_, \uc8051golden_1.IRAM[129] [2]);
  buf _49717_ (_07792_, \uc8051golden_1.IRAM[129] [3]);
  buf _49718_ (_07793_, \uc8051golden_1.IRAM[129] [4]);
  buf _49719_ (_07794_, \uc8051golden_1.IRAM[129] [5]);
  buf _49720_ (_07795_, \uc8051golden_1.IRAM[129] [6]);
  buf _49721_ (_07797_, \uc8051golden_1.IRAM[129] [7]);
  buf _49722_ (_07798_, \uc8051golden_1.IRAM[130] [0]);
  buf _49723_ (_07799_, \uc8051golden_1.IRAM[130] [1]);
  buf _49724_ (_07800_, \uc8051golden_1.IRAM[130] [2]);
  buf _49725_ (_07801_, \uc8051golden_1.IRAM[130] [3]);
  buf _49726_ (_07802_, \uc8051golden_1.IRAM[130] [4]);
  buf _49727_ (_07803_, \uc8051golden_1.IRAM[130] [5]);
  buf _49728_ (_07804_, \uc8051golden_1.IRAM[130] [6]);
  buf _49729_ (_07805_, \uc8051golden_1.IRAM[130] [7]);
  buf _49730_ (_07806_, \uc8051golden_1.IRAM[131] [0]);
  buf _49731_ (_07807_, \uc8051golden_1.IRAM[131] [1]);
  buf _49732_ (_07808_, \uc8051golden_1.IRAM[131] [2]);
  buf _49733_ (_07809_, \uc8051golden_1.IRAM[131] [3]);
  buf _49734_ (_07810_, \uc8051golden_1.IRAM[131] [4]);
  buf _49735_ (_07811_, \uc8051golden_1.IRAM[131] [5]);
  buf _49736_ (_07812_, \uc8051golden_1.IRAM[131] [6]);
  buf _49737_ (_07813_, \uc8051golden_1.IRAM[131] [7]);
  buf _49738_ (_07814_, \uc8051golden_1.IRAM[132] [0]);
  buf _49739_ (_07815_, \uc8051golden_1.IRAM[132] [1]);
  buf _49740_ (_07816_, \uc8051golden_1.IRAM[132] [2]);
  buf _49741_ (_07817_, \uc8051golden_1.IRAM[132] [3]);
  buf _49742_ (_07818_, \uc8051golden_1.IRAM[132] [4]);
  buf _49743_ (_07819_, \uc8051golden_1.IRAM[132] [5]);
  buf _49744_ (_07820_, \uc8051golden_1.IRAM[132] [6]);
  buf _49745_ (_07821_, \uc8051golden_1.IRAM[132] [7]);
  buf _49746_ (_07822_, \uc8051golden_1.IRAM[133] [0]);
  buf _49747_ (_07823_, \uc8051golden_1.IRAM[133] [1]);
  buf _49748_ (_07824_, \uc8051golden_1.IRAM[133] [2]);
  buf _49749_ (_07825_, \uc8051golden_1.IRAM[133] [3]);
  buf _49750_ (_07826_, \uc8051golden_1.IRAM[133] [4]);
  buf _49751_ (_07827_, \uc8051golden_1.IRAM[133] [5]);
  buf _49752_ (_07828_, \uc8051golden_1.IRAM[133] [6]);
  buf _49753_ (_07829_, \uc8051golden_1.IRAM[133] [7]);
  buf _49754_ (_07831_, \uc8051golden_1.IRAM[134] [0]);
  buf _49755_ (_07832_, \uc8051golden_1.IRAM[134] [1]);
  buf _49756_ (_07833_, \uc8051golden_1.IRAM[134] [2]);
  buf _49757_ (_07834_, \uc8051golden_1.IRAM[134] [3]);
  buf _49758_ (_07835_, \uc8051golden_1.IRAM[134] [4]);
  buf _49759_ (_07836_, \uc8051golden_1.IRAM[134] [5]);
  buf _49760_ (_07837_, \uc8051golden_1.IRAM[134] [6]);
  buf _49761_ (_07838_, \uc8051golden_1.IRAM[134] [7]);
  buf _49762_ (_07839_, \uc8051golden_1.IRAM[135] [0]);
  buf _49763_ (_07840_, \uc8051golden_1.IRAM[135] [1]);
  buf _49764_ (_07841_, \uc8051golden_1.IRAM[135] [2]);
  buf _49765_ (_07842_, \uc8051golden_1.IRAM[135] [3]);
  buf _49766_ (_07843_, \uc8051golden_1.IRAM[135] [4]);
  buf _49767_ (_07844_, \uc8051golden_1.IRAM[135] [5]);
  buf _49768_ (_07845_, \uc8051golden_1.IRAM[135] [6]);
  buf _49769_ (_07846_, \uc8051golden_1.IRAM[135] [7]);
  buf _49770_ (_07847_, \uc8051golden_1.IRAM[136] [0]);
  buf _49771_ (_07848_, \uc8051golden_1.IRAM[136] [1]);
  buf _49772_ (_07849_, \uc8051golden_1.IRAM[136] [2]);
  buf _49773_ (_07850_, \uc8051golden_1.IRAM[136] [3]);
  buf _49774_ (_07851_, \uc8051golden_1.IRAM[136] [4]);
  buf _49775_ (_07852_, \uc8051golden_1.IRAM[136] [5]);
  buf _49776_ (_07853_, \uc8051golden_1.IRAM[136] [6]);
  buf _49777_ (_07854_, \uc8051golden_1.IRAM[136] [7]);
  buf _49778_ (_07855_, \uc8051golden_1.IRAM[137] [0]);
  buf _49779_ (_07856_, \uc8051golden_1.IRAM[137] [1]);
  buf _49780_ (_07857_, \uc8051golden_1.IRAM[137] [2]);
  buf _49781_ (_07858_, \uc8051golden_1.IRAM[137] [3]);
  buf _49782_ (_07859_, \uc8051golden_1.IRAM[137] [4]);
  buf _49783_ (_07860_, \uc8051golden_1.IRAM[137] [5]);
  buf _49784_ (_07861_, \uc8051golden_1.IRAM[137] [6]);
  buf _49785_ (_07862_, \uc8051golden_1.IRAM[137] [7]);
  buf _49786_ (_07863_, \uc8051golden_1.IRAM[138] [0]);
  buf _49787_ (_07865_, \uc8051golden_1.IRAM[138] [1]);
  buf _49788_ (_07866_, \uc8051golden_1.IRAM[138] [2]);
  buf _49789_ (_07867_, \uc8051golden_1.IRAM[138] [3]);
  buf _49790_ (_07868_, \uc8051golden_1.IRAM[138] [4]);
  buf _49791_ (_07869_, \uc8051golden_1.IRAM[138] [5]);
  buf _49792_ (_07870_, \uc8051golden_1.IRAM[138] [6]);
  buf _49793_ (_07871_, \uc8051golden_1.IRAM[138] [7]);
  buf _49794_ (_07872_, \uc8051golden_1.IRAM[139] [0]);
  buf _49795_ (_07873_, \uc8051golden_1.IRAM[139] [1]);
  buf _49796_ (_07874_, \uc8051golden_1.IRAM[139] [2]);
  buf _49797_ (_07875_, \uc8051golden_1.IRAM[139] [3]);
  buf _49798_ (_07876_, \uc8051golden_1.IRAM[139] [4]);
  buf _49799_ (_07877_, \uc8051golden_1.IRAM[139] [5]);
  buf _49800_ (_07878_, \uc8051golden_1.IRAM[139] [6]);
  buf _49801_ (_07879_, \uc8051golden_1.IRAM[139] [7]);
  buf _49802_ (_07880_, \uc8051golden_1.IRAM[140] [0]);
  buf _49803_ (_07881_, \uc8051golden_1.IRAM[140] [1]);
  buf _49804_ (_07882_, \uc8051golden_1.IRAM[140] [2]);
  buf _49805_ (_07883_, \uc8051golden_1.IRAM[140] [3]);
  buf _49806_ (_07884_, \uc8051golden_1.IRAM[140] [4]);
  buf _49807_ (_07885_, \uc8051golden_1.IRAM[140] [5]);
  buf _49808_ (_07886_, \uc8051golden_1.IRAM[140] [6]);
  buf _49809_ (_07887_, \uc8051golden_1.IRAM[140] [7]);
  buf _49810_ (_07888_, \uc8051golden_1.IRAM[141] [0]);
  buf _49811_ (_07889_, \uc8051golden_1.IRAM[141] [1]);
  buf _49812_ (_07890_, \uc8051golden_1.IRAM[141] [2]);
  buf _49813_ (_07891_, \uc8051golden_1.IRAM[141] [3]);
  buf _49814_ (_07892_, \uc8051golden_1.IRAM[141] [4]);
  buf _49815_ (_07893_, \uc8051golden_1.IRAM[141] [5]);
  buf _49816_ (_07894_, \uc8051golden_1.IRAM[141] [6]);
  buf _49817_ (_07895_, \uc8051golden_1.IRAM[141] [7]);
  buf _49818_ (_07896_, \uc8051golden_1.IRAM[142] [0]);
  buf _49819_ (_07897_, \uc8051golden_1.IRAM[142] [1]);
  buf _49820_ (_07898_, \uc8051golden_1.IRAM[142] [2]);
  buf _49821_ (_07900_, \uc8051golden_1.IRAM[142] [3]);
  buf _49822_ (_07901_, \uc8051golden_1.IRAM[142] [4]);
  buf _49823_ (_07902_, \uc8051golden_1.IRAM[142] [5]);
  buf _49824_ (_07903_, \uc8051golden_1.IRAM[142] [6]);
  buf _49825_ (_07904_, \uc8051golden_1.IRAM[142] [7]);
  buf _49826_ (_07905_, \uc8051golden_1.IRAM[143] [0]);
  buf _49827_ (_07906_, \uc8051golden_1.IRAM[143] [1]);
  buf _49828_ (_07907_, \uc8051golden_1.IRAM[143] [2]);
  buf _49829_ (_07908_, \uc8051golden_1.IRAM[143] [3]);
  buf _49830_ (_07909_, \uc8051golden_1.IRAM[143] [4]);
  buf _49831_ (_07910_, \uc8051golden_1.IRAM[143] [5]);
  buf _49832_ (_07911_, \uc8051golden_1.IRAM[143] [6]);
  buf _49833_ (_07912_, \uc8051golden_1.IRAM[143] [7]);
  buf _49834_ (_07913_, \uc8051golden_1.IRAM[144] [0]);
  buf _49835_ (_07914_, \uc8051golden_1.IRAM[144] [1]);
  buf _49836_ (_07915_, \uc8051golden_1.IRAM[144] [2]);
  buf _49837_ (_07916_, \uc8051golden_1.IRAM[144] [3]);
  buf _49838_ (_07917_, \uc8051golden_1.IRAM[144] [4]);
  buf _49839_ (_07918_, \uc8051golden_1.IRAM[144] [5]);
  buf _49840_ (_07919_, \uc8051golden_1.IRAM[144] [6]);
  buf _49841_ (_07920_, \uc8051golden_1.IRAM[144] [7]);
  buf _49842_ (_07921_, \uc8051golden_1.IRAM[145] [0]);
  buf _49843_ (_07922_, \uc8051golden_1.IRAM[145] [1]);
  buf _49844_ (_07923_, \uc8051golden_1.IRAM[145] [2]);
  buf _49845_ (_07924_, \uc8051golden_1.IRAM[145] [3]);
  buf _49846_ (_07925_, \uc8051golden_1.IRAM[145] [4]);
  buf _49847_ (_07926_, \uc8051golden_1.IRAM[145] [5]);
  buf _49848_ (_07927_, \uc8051golden_1.IRAM[145] [6]);
  buf _49849_ (_07928_, \uc8051golden_1.IRAM[145] [7]);
  buf _49850_ (_07929_, \uc8051golden_1.IRAM[146] [0]);
  buf _49851_ (_07930_, \uc8051golden_1.IRAM[146] [1]);
  buf _49852_ (_07931_, \uc8051golden_1.IRAM[146] [2]);
  buf _49853_ (_07932_, \uc8051golden_1.IRAM[146] [3]);
  buf _49854_ (_07934_, \uc8051golden_1.IRAM[146] [4]);
  buf _49855_ (_07935_, \uc8051golden_1.IRAM[146] [5]);
  buf _49856_ (_07936_, \uc8051golden_1.IRAM[146] [6]);
  buf _49857_ (_07937_, \uc8051golden_1.IRAM[146] [7]);
  buf _49858_ (_07938_, \uc8051golden_1.IRAM[147] [0]);
  buf _49859_ (_07939_, \uc8051golden_1.IRAM[147] [1]);
  buf _49860_ (_07940_, \uc8051golden_1.IRAM[147] [2]);
  buf _49861_ (_07941_, \uc8051golden_1.IRAM[147] [3]);
  buf _49862_ (_07942_, \uc8051golden_1.IRAM[147] [4]);
  buf _49863_ (_07943_, \uc8051golden_1.IRAM[147] [5]);
  buf _49864_ (_07944_, \uc8051golden_1.IRAM[147] [6]);
  buf _49865_ (_07945_, \uc8051golden_1.IRAM[147] [7]);
  buf _49866_ (_07946_, \uc8051golden_1.IRAM[148] [0]);
  buf _49867_ (_07947_, \uc8051golden_1.IRAM[148] [1]);
  buf _49868_ (_07948_, \uc8051golden_1.IRAM[148] [2]);
  buf _49869_ (_07949_, \uc8051golden_1.IRAM[148] [3]);
  buf _49870_ (_07950_, \uc8051golden_1.IRAM[148] [4]);
  buf _49871_ (_07951_, \uc8051golden_1.IRAM[148] [5]);
  buf _49872_ (_07952_, \uc8051golden_1.IRAM[148] [6]);
  buf _49873_ (_07953_, \uc8051golden_1.IRAM[148] [7]);
  buf _49874_ (_07954_, \uc8051golden_1.IRAM[149] [0]);
  buf _49875_ (_07955_, \uc8051golden_1.IRAM[149] [1]);
  buf _49876_ (_07956_, \uc8051golden_1.IRAM[149] [2]);
  buf _49877_ (_07957_, \uc8051golden_1.IRAM[149] [3]);
  buf _49878_ (_07958_, \uc8051golden_1.IRAM[149] [4]);
  buf _49879_ (_07959_, \uc8051golden_1.IRAM[149] [5]);
  buf _49880_ (_07960_, \uc8051golden_1.IRAM[149] [6]);
  buf _49881_ (_07961_, \uc8051golden_1.IRAM[149] [7]);
  buf _49882_ (_07962_, \uc8051golden_1.IRAM[150] [0]);
  buf _49883_ (_07963_, \uc8051golden_1.IRAM[150] [1]);
  buf _49884_ (_07964_, \uc8051golden_1.IRAM[150] [2]);
  buf _49885_ (_07965_, \uc8051golden_1.IRAM[150] [3]);
  buf _49886_ (_07966_, \uc8051golden_1.IRAM[150] [4]);
  buf _49887_ (_07968_, \uc8051golden_1.IRAM[150] [5]);
  buf _49888_ (_07969_, \uc8051golden_1.IRAM[150] [6]);
  buf _49889_ (_07970_, \uc8051golden_1.IRAM[150] [7]);
  buf _49890_ (_07971_, \uc8051golden_1.IRAM[151] [0]);
  buf _49891_ (_07972_, \uc8051golden_1.IRAM[151] [1]);
  buf _49892_ (_07973_, \uc8051golden_1.IRAM[151] [2]);
  buf _49893_ (_07974_, \uc8051golden_1.IRAM[151] [3]);
  buf _49894_ (_07975_, \uc8051golden_1.IRAM[151] [4]);
  buf _49895_ (_07976_, \uc8051golden_1.IRAM[151] [5]);
  buf _49896_ (_07977_, \uc8051golden_1.IRAM[151] [6]);
  buf _49897_ (_07978_, \uc8051golden_1.IRAM[151] [7]);
  buf _49898_ (_07979_, \uc8051golden_1.IRAM[152] [0]);
  buf _49899_ (_07980_, \uc8051golden_1.IRAM[152] [1]);
  buf _49900_ (_07981_, \uc8051golden_1.IRAM[152] [2]);
  buf _49901_ (_07982_, \uc8051golden_1.IRAM[152] [3]);
  buf _49902_ (_07983_, \uc8051golden_1.IRAM[152] [4]);
  buf _49903_ (_07984_, \uc8051golden_1.IRAM[152] [5]);
  buf _49904_ (_07985_, \uc8051golden_1.IRAM[152] [6]);
  buf _49905_ (_07986_, \uc8051golden_1.IRAM[152] [7]);
  buf _49906_ (_07987_, \uc8051golden_1.IRAM[153] [0]);
  buf _49907_ (_07988_, \uc8051golden_1.IRAM[153] [1]);
  buf _49908_ (_07989_, \uc8051golden_1.IRAM[153] [2]);
  buf _49909_ (_07990_, \uc8051golden_1.IRAM[153] [3]);
  buf _49910_ (_07991_, \uc8051golden_1.IRAM[153] [4]);
  buf _49911_ (_07992_, \uc8051golden_1.IRAM[153] [5]);
  buf _49912_ (_07993_, \uc8051golden_1.IRAM[153] [6]);
  buf _49913_ (_07994_, \uc8051golden_1.IRAM[153] [7]);
  buf _49914_ (_07995_, \uc8051golden_1.IRAM[154] [0]);
  buf _49915_ (_07996_, \uc8051golden_1.IRAM[154] [1]);
  buf _49916_ (_07997_, \uc8051golden_1.IRAM[154] [2]);
  buf _49917_ (_07998_, \uc8051golden_1.IRAM[154] [3]);
  buf _49918_ (_07999_, \uc8051golden_1.IRAM[154] [4]);
  buf _49919_ (_08000_, \uc8051golden_1.IRAM[154] [5]);
  buf _49920_ (_08002_, \uc8051golden_1.IRAM[154] [6]);
  buf _49921_ (_08003_, \uc8051golden_1.IRAM[154] [7]);
  buf _49922_ (_08004_, \uc8051golden_1.IRAM[155] [0]);
  buf _49923_ (_08005_, \uc8051golden_1.IRAM[155] [1]);
  buf _49924_ (_08006_, \uc8051golden_1.IRAM[155] [2]);
  buf _49925_ (_08007_, \uc8051golden_1.IRAM[155] [3]);
  buf _49926_ (_08008_, \uc8051golden_1.IRAM[155] [4]);
  buf _49927_ (_08009_, \uc8051golden_1.IRAM[155] [5]);
  buf _49928_ (_08010_, \uc8051golden_1.IRAM[155] [6]);
  buf _49929_ (_08011_, \uc8051golden_1.IRAM[155] [7]);
  buf _49930_ (_08012_, \uc8051golden_1.IRAM[156] [0]);
  buf _49931_ (_08013_, \uc8051golden_1.IRAM[156] [1]);
  buf _49932_ (_08014_, \uc8051golden_1.IRAM[156] [2]);
  buf _49933_ (_08015_, \uc8051golden_1.IRAM[156] [3]);
  buf _49934_ (_08016_, \uc8051golden_1.IRAM[156] [4]);
  buf _49935_ (_08017_, \uc8051golden_1.IRAM[156] [5]);
  buf _49936_ (_08018_, \uc8051golden_1.IRAM[156] [6]);
  buf _49937_ (_08019_, \uc8051golden_1.IRAM[156] [7]);
  buf _49938_ (_08020_, \uc8051golden_1.IRAM[157] [0]);
  buf _49939_ (_08021_, \uc8051golden_1.IRAM[157] [1]);
  buf _49940_ (_08022_, \uc8051golden_1.IRAM[157] [2]);
  buf _49941_ (_08023_, \uc8051golden_1.IRAM[157] [3]);
  buf _49942_ (_08024_, \uc8051golden_1.IRAM[157] [4]);
  buf _49943_ (_08025_, \uc8051golden_1.IRAM[157] [5]);
  buf _49944_ (_08026_, \uc8051golden_1.IRAM[157] [6]);
  buf _49945_ (_08027_, \uc8051golden_1.IRAM[157] [7]);
  buf _49946_ (_08028_, \uc8051golden_1.IRAM[158] [0]);
  buf _49947_ (_08029_, \uc8051golden_1.IRAM[158] [1]);
  buf _49948_ (_08030_, \uc8051golden_1.IRAM[158] [2]);
  buf _49949_ (_08031_, \uc8051golden_1.IRAM[158] [3]);
  buf _49950_ (_08032_, \uc8051golden_1.IRAM[158] [4]);
  buf _49951_ (_08033_, \uc8051golden_1.IRAM[158] [5]);
  buf _49952_ (_08034_, \uc8051golden_1.IRAM[158] [6]);
  buf _49953_ (_08035_, \uc8051golden_1.IRAM[158] [7]);
  buf _49954_ (_08037_, \uc8051golden_1.IRAM[159] [0]);
  buf _49955_ (_08038_, \uc8051golden_1.IRAM[159] [1]);
  buf _49956_ (_08039_, \uc8051golden_1.IRAM[159] [2]);
  buf _49957_ (_08040_, \uc8051golden_1.IRAM[159] [3]);
  buf _49958_ (_08041_, \uc8051golden_1.IRAM[159] [4]);
  buf _49959_ (_08042_, \uc8051golden_1.IRAM[159] [5]);
  buf _49960_ (_08043_, \uc8051golden_1.IRAM[159] [6]);
  buf _49961_ (_08044_, \uc8051golden_1.IRAM[159] [7]);
  buf _49962_ (_08045_, \uc8051golden_1.IRAM[160] [0]);
  buf _49963_ (_08046_, \uc8051golden_1.IRAM[160] [1]);
  buf _49964_ (_08047_, \uc8051golden_1.IRAM[160] [2]);
  buf _49965_ (_08048_, \uc8051golden_1.IRAM[160] [3]);
  buf _49966_ (_08049_, \uc8051golden_1.IRAM[160] [4]);
  buf _49967_ (_08050_, \uc8051golden_1.IRAM[160] [5]);
  buf _49968_ (_08051_, \uc8051golden_1.IRAM[160] [6]);
  buf _49969_ (_08052_, \uc8051golden_1.IRAM[160] [7]);
  buf _49970_ (_08053_, \uc8051golden_1.IRAM[161] [0]);
  buf _49971_ (_08054_, \uc8051golden_1.IRAM[161] [1]);
  buf _49972_ (_08055_, \uc8051golden_1.IRAM[161] [2]);
  buf _49973_ (_08056_, \uc8051golden_1.IRAM[161] [3]);
  buf _49974_ (_08057_, \uc8051golden_1.IRAM[161] [4]);
  buf _49975_ (_08058_, \uc8051golden_1.IRAM[161] [5]);
  buf _49976_ (_08059_, \uc8051golden_1.IRAM[161] [6]);
  buf _49977_ (_08060_, \uc8051golden_1.IRAM[161] [7]);
  buf _49978_ (_08061_, \uc8051golden_1.IRAM[162] [0]);
  buf _49979_ (_08062_, \uc8051golden_1.IRAM[162] [1]);
  buf _49980_ (_08063_, \uc8051golden_1.IRAM[162] [2]);
  buf _49981_ (_08064_, \uc8051golden_1.IRAM[162] [3]);
  buf _49982_ (_08065_, \uc8051golden_1.IRAM[162] [4]);
  buf _49983_ (_08066_, \uc8051golden_1.IRAM[162] [5]);
  buf _49984_ (_08067_, \uc8051golden_1.IRAM[162] [6]);
  buf _49985_ (_08068_, \uc8051golden_1.IRAM[162] [7]);
  buf _49986_ (_08069_, \uc8051golden_1.IRAM[163] [0]);
  buf _49987_ (_08071_, \uc8051golden_1.IRAM[163] [1]);
  buf _49988_ (_08072_, \uc8051golden_1.IRAM[163] [2]);
  buf _49989_ (_08073_, \uc8051golden_1.IRAM[163] [3]);
  buf _49990_ (_08074_, \uc8051golden_1.IRAM[163] [4]);
  buf _49991_ (_08075_, \uc8051golden_1.IRAM[163] [5]);
  buf _49992_ (_08076_, \uc8051golden_1.IRAM[163] [6]);
  buf _49993_ (_08077_, \uc8051golden_1.IRAM[163] [7]);
  buf _49994_ (_08078_, \uc8051golden_1.IRAM[164] [0]);
  buf _49995_ (_08079_, \uc8051golden_1.IRAM[164] [1]);
  buf _49996_ (_08080_, \uc8051golden_1.IRAM[164] [2]);
  buf _49997_ (_08081_, \uc8051golden_1.IRAM[164] [3]);
  buf _49998_ (_08082_, \uc8051golden_1.IRAM[164] [4]);
  buf _49999_ (_08083_, \uc8051golden_1.IRAM[164] [5]);
  buf _50000_ (_08084_, \uc8051golden_1.IRAM[164] [6]);
  buf _50001_ (_08085_, \uc8051golden_1.IRAM[164] [7]);
  buf _50002_ (_08086_, \uc8051golden_1.IRAM[165] [0]);
  buf _50003_ (_08087_, \uc8051golden_1.IRAM[165] [1]);
  buf _50004_ (_08088_, \uc8051golden_1.IRAM[165] [2]);
  buf _50005_ (_08089_, \uc8051golden_1.IRAM[165] [3]);
  buf _50006_ (_08090_, \uc8051golden_1.IRAM[165] [4]);
  buf _50007_ (_08091_, \uc8051golden_1.IRAM[165] [5]);
  buf _50008_ (_08092_, \uc8051golden_1.IRAM[165] [6]);
  buf _50009_ (_08093_, \uc8051golden_1.IRAM[165] [7]);
  buf _50010_ (_08094_, \uc8051golden_1.IRAM[166] [0]);
  buf _50011_ (_08095_, \uc8051golden_1.IRAM[166] [1]);
  buf _50012_ (_08096_, \uc8051golden_1.IRAM[166] [2]);
  buf _50013_ (_08097_, \uc8051golden_1.IRAM[166] [3]);
  buf _50014_ (_08098_, \uc8051golden_1.IRAM[166] [4]);
  buf _50015_ (_08099_, \uc8051golden_1.IRAM[166] [5]);
  buf _50016_ (_08100_, \uc8051golden_1.IRAM[166] [6]);
  buf _50017_ (_08101_, \uc8051golden_1.IRAM[166] [7]);
  buf _50018_ (_08102_, \uc8051golden_1.IRAM[167] [0]);
  buf _50019_ (_08103_, \uc8051golden_1.IRAM[167] [1]);
  buf _50020_ (_08105_, \uc8051golden_1.IRAM[167] [2]);
  buf _50021_ (_08106_, \uc8051golden_1.IRAM[167] [3]);
  buf _50022_ (_08107_, \uc8051golden_1.IRAM[167] [4]);
  buf _50023_ (_08108_, \uc8051golden_1.IRAM[167] [5]);
  buf _50024_ (_08109_, \uc8051golden_1.IRAM[167] [6]);
  buf _50025_ (_08110_, \uc8051golden_1.IRAM[167] [7]);
  buf _50026_ (_08111_, \uc8051golden_1.IRAM[168] [0]);
  buf _50027_ (_08112_, \uc8051golden_1.IRAM[168] [1]);
  buf _50028_ (_08113_, \uc8051golden_1.IRAM[168] [2]);
  buf _50029_ (_08114_, \uc8051golden_1.IRAM[168] [3]);
  buf _50030_ (_08115_, \uc8051golden_1.IRAM[168] [4]);
  buf _50031_ (_08116_, \uc8051golden_1.IRAM[168] [5]);
  buf _50032_ (_08117_, \uc8051golden_1.IRAM[168] [6]);
  buf _50033_ (_08118_, \uc8051golden_1.IRAM[168] [7]);
  buf _50034_ (_08119_, \uc8051golden_1.IRAM[169] [0]);
  buf _50035_ (_08120_, \uc8051golden_1.IRAM[169] [1]);
  buf _50036_ (_08121_, \uc8051golden_1.IRAM[169] [2]);
  buf _50037_ (_08122_, \uc8051golden_1.IRAM[169] [3]);
  buf _50038_ (_08123_, \uc8051golden_1.IRAM[169] [4]);
  buf _50039_ (_08124_, \uc8051golden_1.IRAM[169] [5]);
  buf _50040_ (_08125_, \uc8051golden_1.IRAM[169] [6]);
  buf _50041_ (_08126_, \uc8051golden_1.IRAM[169] [7]);
  buf _50042_ (_08127_, \uc8051golden_1.IRAM[170] [0]);
  buf _50043_ (_08128_, \uc8051golden_1.IRAM[170] [1]);
  buf _50044_ (_08129_, \uc8051golden_1.IRAM[170] [2]);
  buf _50045_ (_08130_, \uc8051golden_1.IRAM[170] [3]);
  buf _50046_ (_08131_, \uc8051golden_1.IRAM[170] [4]);
  buf _50047_ (_08132_, \uc8051golden_1.IRAM[170] [5]);
  buf _50048_ (_08133_, \uc8051golden_1.IRAM[170] [6]);
  buf _50049_ (_08134_, \uc8051golden_1.IRAM[170] [7]);
  buf _50050_ (_08135_, \uc8051golden_1.IRAM[171] [0]);
  buf _50051_ (_08136_, \uc8051golden_1.IRAM[171] [1]);
  buf _50052_ (_08137_, \uc8051golden_1.IRAM[171] [2]);
  buf _50053_ (_08139_, \uc8051golden_1.IRAM[171] [3]);
  buf _50054_ (_08140_, \uc8051golden_1.IRAM[171] [4]);
  buf _50055_ (_08141_, \uc8051golden_1.IRAM[171] [5]);
  buf _50056_ (_08142_, \uc8051golden_1.IRAM[171] [6]);
  buf _50057_ (_08143_, \uc8051golden_1.IRAM[171] [7]);
  buf _50058_ (_08144_, \uc8051golden_1.IRAM[172] [0]);
  buf _50059_ (_08145_, \uc8051golden_1.IRAM[172] [1]);
  buf _50060_ (_08146_, \uc8051golden_1.IRAM[172] [2]);
  buf _50061_ (_08147_, \uc8051golden_1.IRAM[172] [3]);
  buf _50062_ (_08148_, \uc8051golden_1.IRAM[172] [4]);
  buf _50063_ (_08149_, \uc8051golden_1.IRAM[172] [5]);
  buf _50064_ (_08150_, \uc8051golden_1.IRAM[172] [6]);
  buf _50065_ (_08151_, \uc8051golden_1.IRAM[172] [7]);
  buf _50066_ (_08152_, \uc8051golden_1.IRAM[173] [0]);
  buf _50067_ (_08153_, \uc8051golden_1.IRAM[173] [1]);
  buf _50068_ (_08154_, \uc8051golden_1.IRAM[173] [2]);
  buf _50069_ (_08155_, \uc8051golden_1.IRAM[173] [3]);
  buf _50070_ (_08156_, \uc8051golden_1.IRAM[173] [4]);
  buf _50071_ (_08157_, \uc8051golden_1.IRAM[173] [5]);
  buf _50072_ (_08158_, \uc8051golden_1.IRAM[173] [6]);
  buf _50073_ (_08159_, \uc8051golden_1.IRAM[173] [7]);
  buf _50074_ (_08160_, \uc8051golden_1.IRAM[174] [0]);
  buf _50075_ (_08161_, \uc8051golden_1.IRAM[174] [1]);
  buf _50076_ (_08162_, \uc8051golden_1.IRAM[174] [2]);
  buf _50077_ (_08163_, \uc8051golden_1.IRAM[174] [3]);
  buf _50078_ (_08164_, \uc8051golden_1.IRAM[174] [4]);
  buf _50079_ (_08165_, \uc8051golden_1.IRAM[174] [5]);
  buf _50080_ (_08166_, \uc8051golden_1.IRAM[174] [6]);
  buf _50081_ (_08167_, \uc8051golden_1.IRAM[174] [7]);
  buf _50082_ (_08168_, \uc8051golden_1.IRAM[175] [0]);
  buf _50083_ (_08169_, \uc8051golden_1.IRAM[175] [1]);
  buf _50084_ (_08170_, \uc8051golden_1.IRAM[175] [2]);
  buf _50085_ (_08171_, \uc8051golden_1.IRAM[175] [3]);
  buf _50086_ (_08172_, \uc8051golden_1.IRAM[175] [4]);
  buf _50087_ (_08174_, \uc8051golden_1.IRAM[175] [5]);
  buf _50088_ (_08175_, \uc8051golden_1.IRAM[175] [6]);
  buf _50089_ (_08176_, \uc8051golden_1.IRAM[175] [7]);
  buf _50090_ (_08177_, \uc8051golden_1.IRAM[176] [0]);
  buf _50091_ (_08178_, \uc8051golden_1.IRAM[176] [1]);
  buf _50092_ (_08179_, \uc8051golden_1.IRAM[176] [2]);
  buf _50093_ (_08180_, \uc8051golden_1.IRAM[176] [3]);
  buf _50094_ (_08181_, \uc8051golden_1.IRAM[176] [4]);
  buf _50095_ (_08182_, \uc8051golden_1.IRAM[176] [5]);
  buf _50096_ (_08183_, \uc8051golden_1.IRAM[176] [6]);
  buf _50097_ (_08184_, \uc8051golden_1.IRAM[176] [7]);
  buf _50098_ (_08185_, \uc8051golden_1.IRAM[177] [0]);
  buf _50099_ (_08186_, \uc8051golden_1.IRAM[177] [1]);
  buf _50100_ (_08187_, \uc8051golden_1.IRAM[177] [2]);
  buf _50101_ (_08188_, \uc8051golden_1.IRAM[177] [3]);
  buf _50102_ (_08189_, \uc8051golden_1.IRAM[177] [4]);
  buf _50103_ (_08190_, \uc8051golden_1.IRAM[177] [5]);
  buf _50104_ (_08191_, \uc8051golden_1.IRAM[177] [6]);
  buf _50105_ (_08192_, \uc8051golden_1.IRAM[177] [7]);
  buf _50106_ (_08193_, \uc8051golden_1.IRAM[178] [0]);
  buf _50107_ (_08194_, \uc8051golden_1.IRAM[178] [1]);
  buf _50108_ (_08195_, \uc8051golden_1.IRAM[178] [2]);
  buf _50109_ (_08196_, \uc8051golden_1.IRAM[178] [3]);
  buf _50110_ (_08197_, \uc8051golden_1.IRAM[178] [4]);
  buf _50111_ (_08198_, \uc8051golden_1.IRAM[178] [5]);
  buf _50112_ (_08199_, \uc8051golden_1.IRAM[178] [6]);
  buf _50113_ (_08200_, \uc8051golden_1.IRAM[178] [7]);
  buf _50114_ (_08201_, \uc8051golden_1.IRAM[179] [0]);
  buf _50115_ (_08202_, \uc8051golden_1.IRAM[179] [1]);
  buf _50116_ (_08203_, \uc8051golden_1.IRAM[179] [2]);
  buf _50117_ (_08204_, \uc8051golden_1.IRAM[179] [3]);
  buf _50118_ (_08205_, \uc8051golden_1.IRAM[179] [4]);
  buf _50119_ (_08206_, \uc8051golden_1.IRAM[179] [5]);
  buf _50120_ (_08208_, \uc8051golden_1.IRAM[179] [6]);
  buf _50121_ (_08209_, \uc8051golden_1.IRAM[179] [7]);
  buf _50122_ (_08210_, \uc8051golden_1.IRAM[180] [0]);
  buf _50123_ (_08211_, \uc8051golden_1.IRAM[180] [1]);
  buf _50124_ (_08212_, \uc8051golden_1.IRAM[180] [2]);
  buf _50125_ (_08213_, \uc8051golden_1.IRAM[180] [3]);
  buf _50126_ (_08214_, \uc8051golden_1.IRAM[180] [4]);
  buf _50127_ (_08215_, \uc8051golden_1.IRAM[180] [5]);
  buf _50128_ (_08216_, \uc8051golden_1.IRAM[180] [6]);
  buf _50129_ (_08217_, \uc8051golden_1.IRAM[180] [7]);
  buf _50130_ (_08218_, \uc8051golden_1.IRAM[181] [0]);
  buf _50131_ (_08219_, \uc8051golden_1.IRAM[181] [1]);
  buf _50132_ (_08220_, \uc8051golden_1.IRAM[181] [2]);
  buf _50133_ (_08221_, \uc8051golden_1.IRAM[181] [3]);
  buf _50134_ (_08222_, \uc8051golden_1.IRAM[181] [4]);
  buf _50135_ (_08223_, \uc8051golden_1.IRAM[181] [5]);
  buf _50136_ (_08224_, \uc8051golden_1.IRAM[181] [6]);
  buf _50137_ (_08225_, \uc8051golden_1.IRAM[181] [7]);
  buf _50138_ (_08226_, \uc8051golden_1.IRAM[182] [0]);
  buf _50139_ (_08227_, \uc8051golden_1.IRAM[182] [1]);
  buf _50140_ (_08228_, \uc8051golden_1.IRAM[182] [2]);
  buf _50141_ (_08229_, \uc8051golden_1.IRAM[182] [3]);
  buf _50142_ (_08230_, \uc8051golden_1.IRAM[182] [4]);
  buf _50143_ (_08231_, \uc8051golden_1.IRAM[182] [5]);
  buf _50144_ (_08232_, \uc8051golden_1.IRAM[182] [6]);
  buf _50145_ (_08233_, \uc8051golden_1.IRAM[182] [7]);
  buf _50146_ (_08234_, \uc8051golden_1.IRAM[183] [0]);
  buf _50147_ (_08235_, \uc8051golden_1.IRAM[183] [1]);
  buf _50148_ (_08236_, \uc8051golden_1.IRAM[183] [2]);
  buf _50149_ (_08237_, \uc8051golden_1.IRAM[183] [3]);
  buf _50150_ (_08238_, \uc8051golden_1.IRAM[183] [4]);
  buf _50151_ (_08239_, \uc8051golden_1.IRAM[183] [5]);
  buf _50152_ (_08240_, \uc8051golden_1.IRAM[183] [6]);
  buf _50153_ (_08242_, \uc8051golden_1.IRAM[183] [7]);
  buf _50154_ (_08243_, \uc8051golden_1.IRAM[184] [0]);
  buf _50155_ (_08244_, \uc8051golden_1.IRAM[184] [1]);
  buf _50156_ (_08245_, \uc8051golden_1.IRAM[184] [2]);
  buf _50157_ (_08246_, \uc8051golden_1.IRAM[184] [3]);
  buf _50158_ (_08247_, \uc8051golden_1.IRAM[184] [4]);
  buf _50159_ (_08248_, \uc8051golden_1.IRAM[184] [5]);
  buf _50160_ (_08249_, \uc8051golden_1.IRAM[184] [6]);
  buf _50161_ (_08250_, \uc8051golden_1.IRAM[184] [7]);
  buf _50162_ (_08251_, \uc8051golden_1.IRAM[185] [0]);
  buf _50163_ (_08252_, \uc8051golden_1.IRAM[185] [1]);
  buf _50164_ (_08253_, \uc8051golden_1.IRAM[185] [2]);
  buf _50165_ (_08254_, \uc8051golden_1.IRAM[185] [3]);
  buf _50166_ (_08255_, \uc8051golden_1.IRAM[185] [4]);
  buf _50167_ (_08256_, \uc8051golden_1.IRAM[185] [5]);
  buf _50168_ (_08257_, \uc8051golden_1.IRAM[185] [6]);
  buf _50169_ (_08258_, \uc8051golden_1.IRAM[185] [7]);
  buf _50170_ (_08259_, \uc8051golden_1.IRAM[186] [0]);
  buf _50171_ (_08260_, \uc8051golden_1.IRAM[186] [1]);
  buf _50172_ (_08261_, \uc8051golden_1.IRAM[186] [2]);
  buf _50173_ (_08262_, \uc8051golden_1.IRAM[186] [3]);
  buf _50174_ (_08263_, \uc8051golden_1.IRAM[186] [4]);
  buf _50175_ (_08264_, \uc8051golden_1.IRAM[186] [5]);
  buf _50176_ (_08265_, \uc8051golden_1.IRAM[186] [6]);
  buf _50177_ (_08266_, \uc8051golden_1.IRAM[186] [7]);
  buf _50178_ (_08267_, \uc8051golden_1.IRAM[187] [0]);
  buf _50179_ (_08268_, \uc8051golden_1.IRAM[187] [1]);
  buf _50180_ (_08269_, \uc8051golden_1.IRAM[187] [2]);
  buf _50181_ (_08270_, \uc8051golden_1.IRAM[187] [3]);
  buf _50182_ (_08271_, \uc8051golden_1.IRAM[187] [4]);
  buf _50183_ (_08272_, \uc8051golden_1.IRAM[187] [5]);
  buf _50184_ (_08273_, \uc8051golden_1.IRAM[187] [6]);
  buf _50185_ (_08274_, \uc8051golden_1.IRAM[187] [7]);
  buf _50186_ (_08276_, \uc8051golden_1.IRAM[188] [0]);
  buf _50187_ (_08277_, \uc8051golden_1.IRAM[188] [1]);
  buf _50188_ (_08278_, \uc8051golden_1.IRAM[188] [2]);
  buf _50189_ (_08279_, \uc8051golden_1.IRAM[188] [3]);
  buf _50190_ (_08280_, \uc8051golden_1.IRAM[188] [4]);
  buf _50191_ (_08281_, \uc8051golden_1.IRAM[188] [5]);
  buf _50192_ (_08282_, \uc8051golden_1.IRAM[188] [6]);
  buf _50193_ (_08283_, \uc8051golden_1.IRAM[188] [7]);
  buf _50194_ (_08284_, \uc8051golden_1.IRAM[189] [0]);
  buf _50195_ (_08285_, \uc8051golden_1.IRAM[189] [1]);
  buf _50196_ (_08286_, \uc8051golden_1.IRAM[189] [2]);
  buf _50197_ (_08287_, \uc8051golden_1.IRAM[189] [3]);
  buf _50198_ (_08288_, \uc8051golden_1.IRAM[189] [4]);
  buf _50199_ (_08289_, \uc8051golden_1.IRAM[189] [5]);
  buf _50200_ (_08290_, \uc8051golden_1.IRAM[189] [6]);
  buf _50201_ (_08291_, \uc8051golden_1.IRAM[189] [7]);
  buf _50202_ (_08292_, \uc8051golden_1.IRAM[190] [0]);
  buf _50203_ (_08293_, \uc8051golden_1.IRAM[190] [1]);
  buf _50204_ (_08294_, \uc8051golden_1.IRAM[190] [2]);
  buf _50205_ (_08295_, \uc8051golden_1.IRAM[190] [3]);
  buf _50206_ (_08296_, \uc8051golden_1.IRAM[190] [4]);
  buf _50207_ (_08297_, \uc8051golden_1.IRAM[190] [5]);
  buf _50208_ (_08298_, \uc8051golden_1.IRAM[190] [6]);
  buf _50209_ (_08299_, \uc8051golden_1.IRAM[190] [7]);
  buf _50210_ (_08300_, \uc8051golden_1.IRAM[191] [0]);
  buf _50211_ (_08301_, \uc8051golden_1.IRAM[191] [1]);
  buf _50212_ (_08302_, \uc8051golden_1.IRAM[191] [2]);
  buf _50213_ (_08303_, \uc8051golden_1.IRAM[191] [3]);
  buf _50214_ (_08304_, \uc8051golden_1.IRAM[191] [4]);
  buf _50215_ (_08305_, \uc8051golden_1.IRAM[191] [5]);
  buf _50216_ (_08306_, \uc8051golden_1.IRAM[191] [6]);
  buf _50217_ (_08307_, \uc8051golden_1.IRAM[191] [7]);
  buf _50218_ (_08308_, \uc8051golden_1.IRAM[192] [0]);
  buf _50219_ (_08310_, \uc8051golden_1.IRAM[192] [1]);
  buf _50220_ (_08311_, \uc8051golden_1.IRAM[192] [2]);
  buf _50221_ (_08312_, \uc8051golden_1.IRAM[192] [3]);
  buf _50222_ (_08313_, \uc8051golden_1.IRAM[192] [4]);
  buf _50223_ (_08314_, \uc8051golden_1.IRAM[192] [5]);
  buf _50224_ (_08315_, \uc8051golden_1.IRAM[192] [6]);
  buf _50225_ (_08316_, \uc8051golden_1.IRAM[192] [7]);
  buf _50226_ (_08317_, \uc8051golden_1.IRAM[193] [0]);
  buf _50227_ (_08318_, \uc8051golden_1.IRAM[193] [1]);
  buf _50228_ (_08319_, \uc8051golden_1.IRAM[193] [2]);
  buf _50229_ (_08320_, \uc8051golden_1.IRAM[193] [3]);
  buf _50230_ (_08321_, \uc8051golden_1.IRAM[193] [4]);
  buf _50231_ (_08322_, \uc8051golden_1.IRAM[193] [5]);
  buf _50232_ (_08323_, \uc8051golden_1.IRAM[193] [6]);
  buf _50233_ (_08324_, \uc8051golden_1.IRAM[193] [7]);
  buf _50234_ (_08325_, \uc8051golden_1.IRAM[194] [0]);
  buf _50235_ (_08326_, \uc8051golden_1.IRAM[194] [1]);
  buf _50236_ (_08327_, \uc8051golden_1.IRAM[194] [2]);
  buf _50237_ (_08328_, \uc8051golden_1.IRAM[194] [3]);
  buf _50238_ (_08329_, \uc8051golden_1.IRAM[194] [4]);
  buf _50239_ (_08330_, \uc8051golden_1.IRAM[194] [5]);
  buf _50240_ (_08331_, \uc8051golden_1.IRAM[194] [6]);
  buf _50241_ (_08332_, \uc8051golden_1.IRAM[194] [7]);
  buf _50242_ (_08333_, \uc8051golden_1.IRAM[195] [0]);
  buf _50243_ (_08334_, \uc8051golden_1.IRAM[195] [1]);
  buf _50244_ (_08335_, \uc8051golden_1.IRAM[195] [2]);
  buf _50245_ (_08336_, \uc8051golden_1.IRAM[195] [3]);
  buf _50246_ (_08337_, \uc8051golden_1.IRAM[195] [4]);
  buf _50247_ (_08338_, \uc8051golden_1.IRAM[195] [5]);
  buf _50248_ (_08339_, \uc8051golden_1.IRAM[195] [6]);
  buf _50249_ (_08340_, \uc8051golden_1.IRAM[195] [7]);
  buf _50250_ (_08341_, \uc8051golden_1.IRAM[196] [0]);
  buf _50251_ (_08342_, \uc8051golden_1.IRAM[196] [1]);
  buf _50252_ (_08344_, \uc8051golden_1.IRAM[196] [2]);
  buf _50253_ (_08345_, \uc8051golden_1.IRAM[196] [3]);
  buf _50254_ (_08346_, \uc8051golden_1.IRAM[196] [4]);
  buf _50255_ (_08347_, \uc8051golden_1.IRAM[196] [5]);
  buf _50256_ (_08348_, \uc8051golden_1.IRAM[196] [6]);
  buf _50257_ (_08349_, \uc8051golden_1.IRAM[196] [7]);
  buf _50258_ (_08350_, \uc8051golden_1.IRAM[197] [0]);
  buf _50259_ (_08351_, \uc8051golden_1.IRAM[197] [1]);
  buf _50260_ (_08352_, \uc8051golden_1.IRAM[197] [2]);
  buf _50261_ (_08353_, \uc8051golden_1.IRAM[197] [3]);
  buf _50262_ (_08354_, \uc8051golden_1.IRAM[197] [4]);
  buf _50263_ (_08355_, \uc8051golden_1.IRAM[197] [5]);
  buf _50264_ (_08356_, \uc8051golden_1.IRAM[197] [6]);
  buf _50265_ (_08357_, \uc8051golden_1.IRAM[197] [7]);
  buf _50266_ (_08358_, \uc8051golden_1.IRAM[198] [0]);
  buf _50267_ (_08359_, \uc8051golden_1.IRAM[198] [1]);
  buf _50268_ (_08360_, \uc8051golden_1.IRAM[198] [2]);
  buf _50269_ (_08361_, \uc8051golden_1.IRAM[198] [3]);
  buf _50270_ (_08362_, \uc8051golden_1.IRAM[198] [4]);
  buf _50271_ (_08363_, \uc8051golden_1.IRAM[198] [5]);
  buf _50272_ (_08364_, \uc8051golden_1.IRAM[198] [6]);
  buf _50273_ (_08365_, \uc8051golden_1.IRAM[198] [7]);
  buf _50274_ (_08366_, \uc8051golden_1.IRAM[199] [0]);
  buf _50275_ (_08367_, \uc8051golden_1.IRAM[199] [1]);
  buf _50276_ (_08368_, \uc8051golden_1.IRAM[199] [2]);
  buf _50277_ (_08369_, \uc8051golden_1.IRAM[199] [3]);
  buf _50278_ (_08370_, \uc8051golden_1.IRAM[199] [4]);
  buf _50279_ (_08371_, \uc8051golden_1.IRAM[199] [5]);
  buf _50280_ (_08372_, \uc8051golden_1.IRAM[199] [6]);
  buf _50281_ (_08373_, \uc8051golden_1.IRAM[199] [7]);
  buf _50282_ (_08374_, \uc8051golden_1.IRAM[200] [0]);
  buf _50283_ (_08375_, \uc8051golden_1.IRAM[200] [1]);
  buf _50284_ (_08376_, \uc8051golden_1.IRAM[200] [2]);
  buf _50285_ (_08377_, \uc8051golden_1.IRAM[200] [3]);
  buf _50286_ (_08379_, \uc8051golden_1.IRAM[200] [4]);
  buf _50287_ (_08380_, \uc8051golden_1.IRAM[200] [5]);
  buf _50288_ (_08381_, \uc8051golden_1.IRAM[200] [6]);
  buf _50289_ (_08382_, \uc8051golden_1.IRAM[200] [7]);
  buf _50290_ (_08383_, \uc8051golden_1.IRAM[201] [0]);
  buf _50291_ (_08384_, \uc8051golden_1.IRAM[201] [1]);
  buf _50292_ (_08385_, \uc8051golden_1.IRAM[201] [2]);
  buf _50293_ (_08386_, \uc8051golden_1.IRAM[201] [3]);
  buf _50294_ (_08387_, \uc8051golden_1.IRAM[201] [4]);
  buf _50295_ (_08388_, \uc8051golden_1.IRAM[201] [5]);
  buf _50296_ (_08389_, \uc8051golden_1.IRAM[201] [6]);
  buf _50297_ (_08390_, \uc8051golden_1.IRAM[201] [7]);
  buf _50298_ (_08391_, \uc8051golden_1.IRAM[202] [0]);
  buf _50299_ (_08392_, \uc8051golden_1.IRAM[202] [1]);
  buf _50300_ (_08393_, \uc8051golden_1.IRAM[202] [2]);
  buf _50301_ (_08394_, \uc8051golden_1.IRAM[202] [3]);
  buf _50302_ (_08395_, \uc8051golden_1.IRAM[202] [4]);
  buf _50303_ (_08396_, \uc8051golden_1.IRAM[202] [5]);
  buf _50304_ (_08397_, \uc8051golden_1.IRAM[202] [6]);
  buf _50305_ (_08398_, \uc8051golden_1.IRAM[202] [7]);
  buf _50306_ (_08399_, \uc8051golden_1.IRAM[203] [0]);
  buf _50307_ (_08400_, \uc8051golden_1.IRAM[203] [1]);
  buf _50308_ (_08401_, \uc8051golden_1.IRAM[203] [2]);
  buf _50309_ (_08402_, \uc8051golden_1.IRAM[203] [3]);
  buf _50310_ (_08403_, \uc8051golden_1.IRAM[203] [4]);
  buf _50311_ (_08404_, \uc8051golden_1.IRAM[203] [5]);
  buf _50312_ (_08405_, \uc8051golden_1.IRAM[203] [6]);
  buf _50313_ (_08406_, \uc8051golden_1.IRAM[203] [7]);
  buf _50314_ (_08407_, \uc8051golden_1.IRAM[204] [0]);
  buf _50315_ (_08408_, \uc8051golden_1.IRAM[204] [1]);
  buf _50316_ (_08409_, \uc8051golden_1.IRAM[204] [2]);
  buf _50317_ (_08410_, \uc8051golden_1.IRAM[204] [3]);
  buf _50318_ (_08411_, \uc8051golden_1.IRAM[204] [4]);
  buf _50319_ (_08413_, \uc8051golden_1.IRAM[204] [5]);
  buf _50320_ (_08414_, \uc8051golden_1.IRAM[204] [6]);
  buf _50321_ (_08415_, \uc8051golden_1.IRAM[204] [7]);
  buf _50322_ (_08416_, \uc8051golden_1.IRAM[205] [0]);
  buf _50323_ (_08417_, \uc8051golden_1.IRAM[205] [1]);
  buf _50324_ (_08418_, \uc8051golden_1.IRAM[205] [2]);
  buf _50325_ (_08419_, \uc8051golden_1.IRAM[205] [3]);
  buf _50326_ (_08420_, \uc8051golden_1.IRAM[205] [4]);
  buf _50327_ (_08421_, \uc8051golden_1.IRAM[205] [5]);
  buf _50328_ (_08422_, \uc8051golden_1.IRAM[205] [6]);
  buf _50329_ (_08423_, \uc8051golden_1.IRAM[205] [7]);
  buf _50330_ (_08424_, \uc8051golden_1.IRAM[206] [0]);
  buf _50331_ (_08425_, \uc8051golden_1.IRAM[206] [1]);
  buf _50332_ (_08426_, \uc8051golden_1.IRAM[206] [2]);
  buf _50333_ (_08427_, \uc8051golden_1.IRAM[206] [3]);
  buf _50334_ (_08428_, \uc8051golden_1.IRAM[206] [4]);
  buf _50335_ (_08429_, \uc8051golden_1.IRAM[206] [5]);
  buf _50336_ (_08430_, \uc8051golden_1.IRAM[206] [6]);
  buf _50337_ (_08431_, \uc8051golden_1.IRAM[206] [7]);
  buf _50338_ (_08432_, \uc8051golden_1.IRAM[207] [0]);
  buf _50339_ (_08433_, \uc8051golden_1.IRAM[207] [1]);
  buf _50340_ (_08434_, \uc8051golden_1.IRAM[207] [2]);
  buf _50341_ (_08435_, \uc8051golden_1.IRAM[207] [3]);
  buf _50342_ (_08436_, \uc8051golden_1.IRAM[207] [4]);
  buf _50343_ (_08437_, \uc8051golden_1.IRAM[207] [5]);
  buf _50344_ (_08438_, \uc8051golden_1.IRAM[207] [6]);
  buf _50345_ (_08439_, \uc8051golden_1.IRAM[207] [7]);
  buf _50346_ (_08440_, \uc8051golden_1.IRAM[208] [0]);
  buf _50347_ (_08441_, \uc8051golden_1.IRAM[208] [1]);
  buf _50348_ (_08442_, \uc8051golden_1.IRAM[208] [2]);
  buf _50349_ (_08443_, \uc8051golden_1.IRAM[208] [3]);
  buf _50350_ (_08444_, \uc8051golden_1.IRAM[208] [4]);
  buf _50351_ (_08445_, \uc8051golden_1.IRAM[208] [5]);
  buf _50352_ (_08447_, \uc8051golden_1.IRAM[208] [6]);
  buf _50353_ (_08448_, \uc8051golden_1.IRAM[208] [7]);
  buf _50354_ (_08449_, \uc8051golden_1.IRAM[209] [0]);
  buf _50355_ (_08450_, \uc8051golden_1.IRAM[209] [1]);
  buf _50356_ (_08451_, \uc8051golden_1.IRAM[209] [2]);
  buf _50357_ (_08452_, \uc8051golden_1.IRAM[209] [3]);
  buf _50358_ (_08453_, \uc8051golden_1.IRAM[209] [4]);
  buf _50359_ (_08454_, \uc8051golden_1.IRAM[209] [5]);
  buf _50360_ (_08455_, \uc8051golden_1.IRAM[209] [6]);
  buf _50361_ (_08456_, \uc8051golden_1.IRAM[209] [7]);
  buf _50362_ (_08457_, \uc8051golden_1.IRAM[210] [0]);
  buf _50363_ (_08458_, \uc8051golden_1.IRAM[210] [1]);
  buf _50364_ (_08459_, \uc8051golden_1.IRAM[210] [2]);
  buf _50365_ (_08460_, \uc8051golden_1.IRAM[210] [3]);
  buf _50366_ (_08461_, \uc8051golden_1.IRAM[210] [4]);
  buf _50367_ (_08462_, \uc8051golden_1.IRAM[210] [5]);
  buf _50368_ (_08463_, \uc8051golden_1.IRAM[210] [6]);
  buf _50369_ (_08464_, \uc8051golden_1.IRAM[210] [7]);
  buf _50370_ (_08465_, \uc8051golden_1.IRAM[211] [0]);
  buf _50371_ (_08466_, \uc8051golden_1.IRAM[211] [1]);
  buf _50372_ (_08467_, \uc8051golden_1.IRAM[211] [2]);
  buf _50373_ (_08468_, \uc8051golden_1.IRAM[211] [3]);
  buf _50374_ (_08469_, \uc8051golden_1.IRAM[211] [4]);
  buf _50375_ (_08470_, \uc8051golden_1.IRAM[211] [5]);
  buf _50376_ (_08471_, \uc8051golden_1.IRAM[211] [6]);
  buf _50377_ (_08472_, \uc8051golden_1.IRAM[211] [7]);
  buf _50378_ (_08473_, \uc8051golden_1.IRAM[212] [0]);
  buf _50379_ (_08474_, \uc8051golden_1.IRAM[212] [1]);
  buf _50380_ (_08475_, \uc8051golden_1.IRAM[212] [2]);
  buf _50381_ (_08476_, \uc8051golden_1.IRAM[212] [3]);
  buf _50382_ (_08477_, \uc8051golden_1.IRAM[212] [4]);
  buf _50383_ (_08478_, \uc8051golden_1.IRAM[212] [5]);
  buf _50384_ (_08479_, \uc8051golden_1.IRAM[212] [6]);
  buf _50385_ (_08480_, \uc8051golden_1.IRAM[212] [7]);
  buf _50386_ (_08482_, \uc8051golden_1.IRAM[213] [0]);
  buf _50387_ (_08483_, \uc8051golden_1.IRAM[213] [1]);
  buf _50388_ (_08484_, \uc8051golden_1.IRAM[213] [2]);
  buf _50389_ (_08485_, \uc8051golden_1.IRAM[213] [3]);
  buf _50390_ (_08486_, \uc8051golden_1.IRAM[213] [4]);
  buf _50391_ (_08487_, \uc8051golden_1.IRAM[213] [5]);
  buf _50392_ (_08488_, \uc8051golden_1.IRAM[213] [6]);
  buf _50393_ (_08489_, \uc8051golden_1.IRAM[213] [7]);
  buf _50394_ (_08490_, \uc8051golden_1.IRAM[214] [0]);
  buf _50395_ (_08491_, \uc8051golden_1.IRAM[214] [1]);
  buf _50396_ (_08492_, \uc8051golden_1.IRAM[214] [2]);
  buf _50397_ (_08493_, \uc8051golden_1.IRAM[214] [3]);
  buf _50398_ (_08494_, \uc8051golden_1.IRAM[214] [4]);
  buf _50399_ (_08495_, \uc8051golden_1.IRAM[214] [5]);
  buf _50400_ (_08496_, \uc8051golden_1.IRAM[214] [6]);
  buf _50401_ (_08497_, \uc8051golden_1.IRAM[214] [7]);
  buf _50402_ (_08498_, \uc8051golden_1.IRAM[215] [0]);
  buf _50403_ (_08499_, \uc8051golden_1.IRAM[215] [1]);
  buf _50404_ (_08500_, \uc8051golden_1.IRAM[215] [2]);
  buf _50405_ (_08501_, \uc8051golden_1.IRAM[215] [3]);
  buf _50406_ (_08502_, \uc8051golden_1.IRAM[215] [4]);
  buf _50407_ (_08503_, \uc8051golden_1.IRAM[215] [5]);
  buf _50408_ (_08504_, \uc8051golden_1.IRAM[215] [6]);
  buf _50409_ (_08505_, \uc8051golden_1.IRAM[215] [7]);
  buf _50410_ (_08506_, \uc8051golden_1.IRAM[216] [0]);
  buf _50411_ (_08507_, \uc8051golden_1.IRAM[216] [1]);
  buf _50412_ (_08508_, \uc8051golden_1.IRAM[216] [2]);
  buf _50413_ (_08509_, \uc8051golden_1.IRAM[216] [3]);
  buf _50414_ (_08510_, \uc8051golden_1.IRAM[216] [4]);
  buf _50415_ (_08511_, \uc8051golden_1.IRAM[216] [5]);
  buf _50416_ (_08512_, \uc8051golden_1.IRAM[216] [6]);
  buf _50417_ (_08513_, \uc8051golden_1.IRAM[216] [7]);
  buf _50418_ (_08514_, \uc8051golden_1.IRAM[217] [0]);
  buf _50419_ (_08516_, \uc8051golden_1.IRAM[217] [1]);
  buf _50420_ (_08517_, \uc8051golden_1.IRAM[217] [2]);
  buf _50421_ (_08518_, \uc8051golden_1.IRAM[217] [3]);
  buf _50422_ (_08519_, \uc8051golden_1.IRAM[217] [4]);
  buf _50423_ (_08520_, \uc8051golden_1.IRAM[217] [5]);
  buf _50424_ (_08521_, \uc8051golden_1.IRAM[217] [6]);
  buf _50425_ (_08522_, \uc8051golden_1.IRAM[217] [7]);
  buf _50426_ (_08523_, \uc8051golden_1.IRAM[218] [0]);
  buf _50427_ (_08524_, \uc8051golden_1.IRAM[218] [1]);
  buf _50428_ (_08525_, \uc8051golden_1.IRAM[218] [2]);
  buf _50429_ (_08526_, \uc8051golden_1.IRAM[218] [3]);
  buf _50430_ (_08527_, \uc8051golden_1.IRAM[218] [4]);
  buf _50431_ (_08528_, \uc8051golden_1.IRAM[218] [5]);
  buf _50432_ (_08529_, \uc8051golden_1.IRAM[218] [6]);
  buf _50433_ (_08530_, \uc8051golden_1.IRAM[218] [7]);
  buf _50434_ (_08531_, \uc8051golden_1.IRAM[219] [0]);
  buf _50435_ (_08532_, \uc8051golden_1.IRAM[219] [1]);
  buf _50436_ (_08533_, \uc8051golden_1.IRAM[219] [2]);
  buf _50437_ (_08534_, \uc8051golden_1.IRAM[219] [3]);
  buf _50438_ (_08535_, \uc8051golden_1.IRAM[219] [4]);
  buf _50439_ (_08536_, \uc8051golden_1.IRAM[219] [5]);
  buf _50440_ (_08537_, \uc8051golden_1.IRAM[219] [6]);
  buf _50441_ (_08538_, \uc8051golden_1.IRAM[219] [7]);
  buf _50442_ (_08539_, \uc8051golden_1.IRAM[220] [0]);
  buf _50443_ (_08540_, \uc8051golden_1.IRAM[220] [1]);
  buf _50444_ (_08541_, \uc8051golden_1.IRAM[220] [2]);
  buf _50445_ (_08542_, \uc8051golden_1.IRAM[220] [3]);
  buf _50446_ (_08543_, \uc8051golden_1.IRAM[220] [4]);
  buf _50447_ (_08544_, \uc8051golden_1.IRAM[220] [5]);
  buf _50448_ (_08545_, \uc8051golden_1.IRAM[220] [6]);
  buf _50449_ (_08546_, \uc8051golden_1.IRAM[220] [7]);
  buf _50450_ (_08547_, \uc8051golden_1.IRAM[221] [0]);
  buf _50451_ (_08548_, \uc8051golden_1.IRAM[221] [1]);
  buf _50452_ (_08550_, \uc8051golden_1.IRAM[221] [2]);
  buf _50453_ (_08551_, \uc8051golden_1.IRAM[221] [3]);
  buf _50454_ (_08552_, \uc8051golden_1.IRAM[221] [4]);
  buf _50455_ (_08553_, \uc8051golden_1.IRAM[221] [5]);
  buf _50456_ (_08554_, \uc8051golden_1.IRAM[221] [6]);
  buf _50457_ (_08555_, \uc8051golden_1.IRAM[221] [7]);
  buf _50458_ (_08556_, \uc8051golden_1.IRAM[222] [0]);
  buf _50459_ (_08557_, \uc8051golden_1.IRAM[222] [1]);
  buf _50460_ (_08558_, \uc8051golden_1.IRAM[222] [2]);
  buf _50461_ (_08559_, \uc8051golden_1.IRAM[222] [3]);
  buf _50462_ (_08560_, \uc8051golden_1.IRAM[222] [4]);
  buf _50463_ (_08561_, \uc8051golden_1.IRAM[222] [5]);
  buf _50464_ (_08562_, \uc8051golden_1.IRAM[222] [6]);
  buf _50465_ (_08563_, \uc8051golden_1.IRAM[222] [7]);
  buf _50466_ (_08564_, \uc8051golden_1.IRAM[223] [0]);
  buf _50467_ (_08565_, \uc8051golden_1.IRAM[223] [1]);
  buf _50468_ (_08566_, \uc8051golden_1.IRAM[223] [2]);
  buf _50469_ (_08567_, \uc8051golden_1.IRAM[223] [3]);
  buf _50470_ (_08568_, \uc8051golden_1.IRAM[223] [4]);
  buf _50471_ (_08569_, \uc8051golden_1.IRAM[223] [5]);
  buf _50472_ (_08570_, \uc8051golden_1.IRAM[223] [6]);
  buf _50473_ (_08571_, \uc8051golden_1.IRAM[223] [7]);
  buf _50474_ (_08572_, \uc8051golden_1.IRAM[224] [0]);
  buf _50475_ (_08573_, \uc8051golden_1.IRAM[224] [1]);
  buf _50476_ (_08574_, \uc8051golden_1.IRAM[224] [2]);
  buf _50477_ (_08575_, \uc8051golden_1.IRAM[224] [3]);
  buf _50478_ (_08576_, \uc8051golden_1.IRAM[224] [4]);
  buf _50479_ (_08577_, \uc8051golden_1.IRAM[224] [5]);
  buf _50480_ (_08578_, \uc8051golden_1.IRAM[224] [6]);
  buf _50481_ (_08579_, \uc8051golden_1.IRAM[224] [7]);
  buf _50482_ (_08580_, \uc8051golden_1.IRAM[225] [0]);
  buf _50483_ (_08581_, \uc8051golden_1.IRAM[225] [1]);
  buf _50484_ (_08582_, \uc8051golden_1.IRAM[225] [2]);
  buf _50485_ (_08584_, \uc8051golden_1.IRAM[225] [3]);
  buf _50486_ (_08585_, \uc8051golden_1.IRAM[225] [4]);
  buf _50487_ (_08586_, \uc8051golden_1.IRAM[225] [5]);
  buf _50488_ (_08587_, \uc8051golden_1.IRAM[225] [6]);
  buf _50489_ (_08588_, \uc8051golden_1.IRAM[225] [7]);
  buf _50490_ (_08589_, \uc8051golden_1.IRAM[226] [0]);
  buf _50491_ (_08590_, \uc8051golden_1.IRAM[226] [1]);
  buf _50492_ (_08591_, \uc8051golden_1.IRAM[226] [2]);
  buf _50493_ (_08592_, \uc8051golden_1.IRAM[226] [3]);
  buf _50494_ (_08593_, \uc8051golden_1.IRAM[226] [4]);
  buf _50495_ (_08594_, \uc8051golden_1.IRAM[226] [5]);
  buf _50496_ (_08595_, \uc8051golden_1.IRAM[226] [6]);
  buf _50497_ (_08596_, \uc8051golden_1.IRAM[226] [7]);
  buf _50498_ (_08597_, \uc8051golden_1.IRAM[227] [0]);
  buf _50499_ (_08598_, \uc8051golden_1.IRAM[227] [1]);
  buf _50500_ (_08599_, \uc8051golden_1.IRAM[227] [2]);
  buf _50501_ (_08600_, \uc8051golden_1.IRAM[227] [3]);
  buf _50502_ (_08601_, \uc8051golden_1.IRAM[227] [4]);
  buf _50503_ (_08602_, \uc8051golden_1.IRAM[227] [5]);
  buf _50504_ (_08603_, \uc8051golden_1.IRAM[227] [6]);
  buf _50505_ (_08604_, \uc8051golden_1.IRAM[227] [7]);
  buf _50506_ (_08605_, \uc8051golden_1.IRAM[228] [0]);
  buf _50507_ (_08606_, \uc8051golden_1.IRAM[228] [1]);
  buf _50508_ (_08607_, \uc8051golden_1.IRAM[228] [2]);
  buf _50509_ (_08608_, \uc8051golden_1.IRAM[228] [3]);
  buf _50510_ (_08609_, \uc8051golden_1.IRAM[228] [4]);
  buf _50511_ (_08610_, \uc8051golden_1.IRAM[228] [5]);
  buf _50512_ (_08611_, \uc8051golden_1.IRAM[228] [6]);
  buf _50513_ (_08612_, \uc8051golden_1.IRAM[228] [7]);
  buf _50514_ (_08613_, \uc8051golden_1.IRAM[229] [0]);
  buf _50515_ (_08614_, \uc8051golden_1.IRAM[229] [1]);
  buf _50516_ (_08615_, \uc8051golden_1.IRAM[229] [2]);
  buf _50517_ (_08616_, \uc8051golden_1.IRAM[229] [3]);
  buf _50518_ (_08618_, \uc8051golden_1.IRAM[229] [4]);
  buf _50519_ (_08619_, \uc8051golden_1.IRAM[229] [5]);
  buf _50520_ (_08620_, \uc8051golden_1.IRAM[229] [6]);
  buf _50521_ (_08621_, \uc8051golden_1.IRAM[229] [7]);
  buf _50522_ (_08622_, \uc8051golden_1.IRAM[230] [0]);
  buf _50523_ (_08623_, \uc8051golden_1.IRAM[230] [1]);
  buf _50524_ (_08624_, \uc8051golden_1.IRAM[230] [2]);
  buf _50525_ (_08625_, \uc8051golden_1.IRAM[230] [3]);
  buf _50526_ (_08626_, \uc8051golden_1.IRAM[230] [4]);
  buf _50527_ (_08627_, \uc8051golden_1.IRAM[230] [5]);
  buf _50528_ (_08628_, \uc8051golden_1.IRAM[230] [6]);
  buf _50529_ (_08629_, \uc8051golden_1.IRAM[230] [7]);
  buf _50530_ (_08630_, \uc8051golden_1.IRAM[231] [0]);
  buf _50531_ (_08631_, \uc8051golden_1.IRAM[231] [1]);
  buf _50532_ (_08632_, \uc8051golden_1.IRAM[231] [2]);
  buf _50533_ (_08633_, \uc8051golden_1.IRAM[231] [3]);
  buf _50534_ (_08634_, \uc8051golden_1.IRAM[231] [4]);
  buf _50535_ (_08635_, \uc8051golden_1.IRAM[231] [5]);
  buf _50536_ (_08636_, \uc8051golden_1.IRAM[231] [6]);
  buf _50537_ (_08637_, \uc8051golden_1.IRAM[231] [7]);
  buf _50538_ (_08638_, \uc8051golden_1.IRAM[232] [0]);
  buf _50539_ (_08639_, \uc8051golden_1.IRAM[232] [1]);
  buf _50540_ (_08640_, \uc8051golden_1.IRAM[232] [2]);
  buf _50541_ (_08641_, \uc8051golden_1.IRAM[232] [3]);
  buf _50542_ (_08642_, \uc8051golden_1.IRAM[232] [4]);
  buf _50543_ (_08643_, \uc8051golden_1.IRAM[232] [5]);
  buf _50544_ (_08644_, \uc8051golden_1.IRAM[232] [6]);
  buf _50545_ (_08645_, \uc8051golden_1.IRAM[232] [7]);
  buf _50546_ (_08646_, \uc8051golden_1.IRAM[233] [0]);
  buf _50547_ (_08647_, \uc8051golden_1.IRAM[233] [1]);
  buf _50548_ (_08648_, \uc8051golden_1.IRAM[233] [2]);
  buf _50549_ (_08649_, \uc8051golden_1.IRAM[233] [3]);
  buf _50550_ (_08650_, \uc8051golden_1.IRAM[233] [4]);
  buf _50551_ (_08651_, \uc8051golden_1.IRAM[233] [5]);
  buf _50552_ (_08653_, \uc8051golden_1.IRAM[233] [6]);
  buf _50553_ (_08654_, \uc8051golden_1.IRAM[233] [7]);
  buf _50554_ (_08655_, \uc8051golden_1.IRAM[234] [0]);
  buf _50555_ (_08656_, \uc8051golden_1.IRAM[234] [1]);
  buf _50556_ (_08657_, \uc8051golden_1.IRAM[234] [2]);
  buf _50557_ (_08658_, \uc8051golden_1.IRAM[234] [3]);
  buf _50558_ (_08659_, \uc8051golden_1.IRAM[234] [4]);
  buf _50559_ (_08660_, \uc8051golden_1.IRAM[234] [5]);
  buf _50560_ (_08661_, \uc8051golden_1.IRAM[234] [6]);
  buf _50561_ (_08662_, \uc8051golden_1.IRAM[234] [7]);
  buf _50562_ (_08663_, \uc8051golden_1.IRAM[235] [0]);
  buf _50563_ (_08664_, \uc8051golden_1.IRAM[235] [1]);
  buf _50564_ (_08665_, \uc8051golden_1.IRAM[235] [2]);
  buf _50565_ (_08666_, \uc8051golden_1.IRAM[235] [3]);
  buf _50566_ (_08667_, \uc8051golden_1.IRAM[235] [4]);
  buf _50567_ (_08668_, \uc8051golden_1.IRAM[235] [5]);
  buf _50568_ (_08669_, \uc8051golden_1.IRAM[235] [6]);
  buf _50569_ (_08670_, \uc8051golden_1.IRAM[235] [7]);
  buf _50570_ (_08671_, \uc8051golden_1.IRAM[236] [0]);
  buf _50571_ (_08672_, \uc8051golden_1.IRAM[236] [1]);
  buf _50572_ (_08673_, \uc8051golden_1.IRAM[236] [2]);
  buf _50573_ (_08674_, \uc8051golden_1.IRAM[236] [3]);
  buf _50574_ (_08675_, \uc8051golden_1.IRAM[236] [4]);
  buf _50575_ (_08676_, \uc8051golden_1.IRAM[236] [5]);
  buf _50576_ (_08677_, \uc8051golden_1.IRAM[236] [6]);
  buf _50577_ (_08678_, \uc8051golden_1.IRAM[236] [7]);
  buf _50578_ (_08679_, \uc8051golden_1.IRAM[237] [0]);
  buf _50579_ (_08680_, \uc8051golden_1.IRAM[237] [1]);
  buf _50580_ (_08681_, \uc8051golden_1.IRAM[237] [2]);
  buf _50581_ (_08682_, \uc8051golden_1.IRAM[237] [3]);
  buf _50582_ (_08683_, \uc8051golden_1.IRAM[237] [4]);
  buf _50583_ (_08684_, \uc8051golden_1.IRAM[237] [5]);
  buf _50584_ (_08685_, \uc8051golden_1.IRAM[237] [6]);
  buf _50585_ (_08687_, \uc8051golden_1.IRAM[237] [7]);
  buf _50586_ (_08688_, \uc8051golden_1.IRAM[238] [0]);
  buf _50587_ (_08689_, \uc8051golden_1.IRAM[238] [1]);
  buf _50588_ (_08690_, \uc8051golden_1.IRAM[238] [2]);
  buf _50589_ (_08691_, \uc8051golden_1.IRAM[238] [3]);
  buf _50590_ (_08692_, \uc8051golden_1.IRAM[238] [4]);
  buf _50591_ (_08693_, \uc8051golden_1.IRAM[238] [5]);
  buf _50592_ (_08694_, \uc8051golden_1.IRAM[238] [6]);
  buf _50593_ (_08695_, \uc8051golden_1.IRAM[238] [7]);
  buf _50594_ (_08696_, \uc8051golden_1.IRAM[239] [0]);
  buf _50595_ (_08697_, \uc8051golden_1.IRAM[239] [1]);
  buf _50596_ (_08698_, \uc8051golden_1.IRAM[239] [2]);
  buf _50597_ (_08699_, \uc8051golden_1.IRAM[239] [3]);
  buf _50598_ (_08700_, \uc8051golden_1.IRAM[239] [4]);
  buf _50599_ (_08701_, \uc8051golden_1.IRAM[239] [5]);
  buf _50600_ (_08702_, \uc8051golden_1.IRAM[239] [6]);
  buf _50601_ (_08703_, \uc8051golden_1.IRAM[239] [7]);
  buf _50602_ (_08704_, \uc8051golden_1.IRAM[240] [0]);
  buf _50603_ (_08705_, \uc8051golden_1.IRAM[240] [1]);
  buf _50604_ (_08706_, \uc8051golden_1.IRAM[240] [2]);
  buf _50605_ (_08707_, \uc8051golden_1.IRAM[240] [3]);
  buf _50606_ (_08708_, \uc8051golden_1.IRAM[240] [4]);
  buf _50607_ (_08709_, \uc8051golden_1.IRAM[240] [5]);
  buf _50608_ (_08710_, \uc8051golden_1.IRAM[240] [6]);
  buf _50609_ (_08711_, \uc8051golden_1.IRAM[240] [7]);
  buf _50610_ (_08712_, \uc8051golden_1.IRAM[241] [0]);
  buf _50611_ (_08713_, \uc8051golden_1.IRAM[241] [1]);
  buf _50612_ (_08714_, \uc8051golden_1.IRAM[241] [2]);
  buf _50613_ (_08715_, \uc8051golden_1.IRAM[241] [3]);
  buf _50614_ (_08716_, \uc8051golden_1.IRAM[241] [4]);
  buf _50615_ (_08717_, \uc8051golden_1.IRAM[241] [5]);
  buf _50616_ (_08718_, \uc8051golden_1.IRAM[241] [6]);
  buf _50617_ (_08719_, \uc8051golden_1.IRAM[241] [7]);
  buf _50618_ (_08721_, \uc8051golden_1.IRAM[242] [0]);
  buf _50619_ (_08722_, \uc8051golden_1.IRAM[242] [1]);
  buf _50620_ (_08723_, \uc8051golden_1.IRAM[242] [2]);
  buf _50621_ (_08724_, \uc8051golden_1.IRAM[242] [3]);
  buf _50622_ (_08725_, \uc8051golden_1.IRAM[242] [4]);
  buf _50623_ (_08726_, \uc8051golden_1.IRAM[242] [5]);
  buf _50624_ (_08727_, \uc8051golden_1.IRAM[242] [6]);
  buf _50625_ (_08728_, \uc8051golden_1.IRAM[242] [7]);
  buf _50626_ (_08729_, \uc8051golden_1.IRAM[243] [0]);
  buf _50627_ (_08730_, \uc8051golden_1.IRAM[243] [1]);
  buf _50628_ (_08731_, \uc8051golden_1.IRAM[243] [2]);
  buf _50629_ (_08732_, \uc8051golden_1.IRAM[243] [3]);
  buf _50630_ (_08733_, \uc8051golden_1.IRAM[243] [4]);
  buf _50631_ (_08734_, \uc8051golden_1.IRAM[243] [5]);
  buf _50632_ (_08735_, \uc8051golden_1.IRAM[243] [6]);
  buf _50633_ (_08736_, \uc8051golden_1.IRAM[243] [7]);
  buf _50634_ (_08737_, \uc8051golden_1.IRAM[244] [0]);
  buf _50635_ (_08738_, \uc8051golden_1.IRAM[244] [1]);
  buf _50636_ (_08739_, \uc8051golden_1.IRAM[244] [2]);
  buf _50637_ (_08740_, \uc8051golden_1.IRAM[244] [3]);
  buf _50638_ (_08741_, \uc8051golden_1.IRAM[244] [4]);
  buf _50639_ (_08742_, \uc8051golden_1.IRAM[244] [5]);
  buf _50640_ (_08743_, \uc8051golden_1.IRAM[244] [6]);
  buf _50641_ (_08744_, \uc8051golden_1.IRAM[244] [7]);
  buf _50642_ (_08745_, \uc8051golden_1.IRAM[245] [0]);
  buf _50643_ (_08746_, \uc8051golden_1.IRAM[245] [1]);
  buf _50644_ (_08747_, \uc8051golden_1.IRAM[245] [2]);
  buf _50645_ (_08748_, \uc8051golden_1.IRAM[245] [3]);
  buf _50646_ (_08749_, \uc8051golden_1.IRAM[245] [4]);
  buf _50647_ (_08750_, \uc8051golden_1.IRAM[245] [5]);
  buf _50648_ (_08751_, \uc8051golden_1.IRAM[245] [6]);
  buf _50649_ (_08752_, \uc8051golden_1.IRAM[245] [7]);
  buf _50650_ (_08753_, \uc8051golden_1.IRAM[246] [0]);
  buf _50651_ (_08755_, \uc8051golden_1.IRAM[246] [1]);
  buf _50652_ (_08756_, \uc8051golden_1.IRAM[246] [2]);
  buf _50653_ (_08757_, \uc8051golden_1.IRAM[246] [3]);
  buf _50654_ (_08758_, \uc8051golden_1.IRAM[246] [4]);
  buf _50655_ (_08759_, \uc8051golden_1.IRAM[246] [5]);
  buf _50656_ (_08760_, \uc8051golden_1.IRAM[246] [6]);
  buf _50657_ (_08761_, \uc8051golden_1.IRAM[246] [7]);
  buf _50658_ (_08762_, \uc8051golden_1.IRAM[247] [0]);
  buf _50659_ (_08763_, \uc8051golden_1.IRAM[247] [1]);
  buf _50660_ (_08764_, \uc8051golden_1.IRAM[247] [2]);
  buf _50661_ (_08765_, \uc8051golden_1.IRAM[247] [3]);
  buf _50662_ (_08766_, \uc8051golden_1.IRAM[247] [4]);
  buf _50663_ (_08767_, \uc8051golden_1.IRAM[247] [5]);
  buf _50664_ (_08768_, \uc8051golden_1.IRAM[247] [6]);
  buf _50665_ (_08769_, \uc8051golden_1.IRAM[247] [7]);
  buf _50666_ (_08770_, \uc8051golden_1.IRAM[248] [0]);
  buf _50667_ (_08771_, \uc8051golden_1.IRAM[248] [1]);
  buf _50668_ (_08772_, \uc8051golden_1.IRAM[248] [2]);
  buf _50669_ (_08773_, \uc8051golden_1.IRAM[248] [3]);
  buf _50670_ (_08774_, \uc8051golden_1.IRAM[248] [4]);
  buf _50671_ (_08775_, \uc8051golden_1.IRAM[248] [5]);
  buf _50672_ (_08776_, \uc8051golden_1.IRAM[248] [6]);
  buf _50673_ (_08777_, \uc8051golden_1.IRAM[248] [7]);
  buf _50674_ (_08778_, \uc8051golden_1.IRAM[249] [0]);
  buf _50675_ (_08779_, \uc8051golden_1.IRAM[249] [1]);
  buf _50676_ (_08780_, \uc8051golden_1.IRAM[249] [2]);
  buf _50677_ (_08781_, \uc8051golden_1.IRAM[249] [3]);
  buf _50678_ (_08782_, \uc8051golden_1.IRAM[249] [4]);
  buf _50679_ (_08783_, \uc8051golden_1.IRAM[249] [5]);
  buf _50680_ (_08784_, \uc8051golden_1.IRAM[249] [6]);
  buf _50681_ (_08785_, \uc8051golden_1.IRAM[249] [7]);
  buf _50682_ (_08786_, \uc8051golden_1.IRAM[250] [0]);
  buf _50683_ (_08787_, \uc8051golden_1.IRAM[250] [1]);
  buf _50684_ (_08788_, \uc8051golden_1.IRAM[250] [2]);
  buf _50685_ (_08790_, \uc8051golden_1.IRAM[250] [3]);
  buf _50686_ (_08791_, \uc8051golden_1.IRAM[250] [4]);
  buf _50687_ (_08792_, \uc8051golden_1.IRAM[250] [5]);
  buf _50688_ (_08793_, \uc8051golden_1.IRAM[250] [6]);
  buf _50689_ (_08794_, \uc8051golden_1.IRAM[250] [7]);
  buf _50690_ (_08795_, \uc8051golden_1.IRAM[251] [0]);
  buf _50691_ (_08796_, \uc8051golden_1.IRAM[251] [1]);
  buf _50692_ (_08797_, \uc8051golden_1.IRAM[251] [2]);
  buf _50693_ (_08798_, \uc8051golden_1.IRAM[251] [3]);
  buf _50694_ (_08799_, \uc8051golden_1.IRAM[251] [4]);
  buf _50695_ (_08800_, \uc8051golden_1.IRAM[251] [5]);
  buf _50696_ (_08801_, \uc8051golden_1.IRAM[251] [6]);
  buf _50697_ (_08802_, \uc8051golden_1.IRAM[251] [7]);
  buf _50698_ (_08803_, \uc8051golden_1.IRAM[252] [0]);
  buf _50699_ (_08804_, \uc8051golden_1.IRAM[252] [1]);
  buf _50700_ (_08805_, \uc8051golden_1.IRAM[252] [2]);
  buf _50701_ (_08806_, \uc8051golden_1.IRAM[252] [3]);
  buf _50702_ (_08807_, \uc8051golden_1.IRAM[252] [4]);
  buf _50703_ (_08808_, \uc8051golden_1.IRAM[252] [5]);
  buf _50704_ (_08809_, \uc8051golden_1.IRAM[252] [6]);
  buf _50705_ (_08810_, \uc8051golden_1.IRAM[252] [7]);
  buf _50706_ (_08811_, \uc8051golden_1.IRAM[253] [0]);
  buf _50707_ (_08812_, \uc8051golden_1.IRAM[253] [1]);
  buf _50708_ (_08813_, \uc8051golden_1.IRAM[253] [2]);
  buf _50709_ (_08814_, \uc8051golden_1.IRAM[253] [3]);
  buf _50710_ (_08815_, \uc8051golden_1.IRAM[253] [4]);
  buf _50711_ (_08816_, \uc8051golden_1.IRAM[253] [5]);
  buf _50712_ (_08817_, \uc8051golden_1.IRAM[253] [6]);
  buf _50713_ (_08818_, \uc8051golden_1.IRAM[253] [7]);
  buf _50714_ (_08819_, \uc8051golden_1.IRAM[254] [0]);
  buf _50715_ (_08820_, \uc8051golden_1.IRAM[254] [1]);
  buf _50716_ (_08821_, \uc8051golden_1.IRAM[254] [2]);
  buf _50717_ (_08822_, \uc8051golden_1.IRAM[254] [3]);
  buf _50718_ (_08824_, \uc8051golden_1.IRAM[254] [4]);
  buf _50719_ (_08825_, \uc8051golden_1.IRAM[254] [5]);
  buf _50720_ (_08826_, \uc8051golden_1.IRAM[254] [6]);
  buf _50721_ (_08827_, \uc8051golden_1.IRAM[254] [7]);
  buf _50722_ (_08828_, \uc8051golden_1.IRAM[255] [0]);
  buf _50723_ (_08829_, \uc8051golden_1.IRAM[255] [1]);
  buf _50724_ (_08830_, \uc8051golden_1.IRAM[255] [2]);
  buf _50725_ (_08831_, \uc8051golden_1.IRAM[255] [3]);
  buf _50726_ (_08832_, \uc8051golden_1.IRAM[255] [4]);
  buf _50727_ (_08833_, \uc8051golden_1.IRAM[255] [5]);
  buf _50728_ (_08834_, \uc8051golden_1.IRAM[255] [6]);
  dff _50729_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02979_, clk);
  dff _50730_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02989_, clk);
  dff _50731_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03009_, clk);
  dff _50732_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03028_, clk);
  dff _50733_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03048_, clk);
  dff _50734_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00912_, clk);
  dff _50735_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03058_, clk);
  dff _50736_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00881_, clk);
  dff _50737_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03069_, clk);
  dff _50738_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03079_, clk);
  dff _50739_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03089_, clk);
  dff _50740_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03100_, clk);
  dff _50741_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03110_, clk);
  dff _50742_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03121_, clk);
  dff _50743_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03131_, clk);
  dff _50744_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00933_, clk);
  dff _50745_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02734_, clk);
  dff _50746_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _25272_, clk);
  dff _50747_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02921_, clk);
  dff _50748_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _03120_, clk);
  dff _50749_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03308_, clk);
  dff _50750_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03499_, clk);
  dff _50751_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03687_, clk);
  dff _50752_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03875_, clk);
  dff _50753_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _04060_, clk);
  dff _50754_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04243_, clk);
  dff _50755_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04339_, clk);
  dff _50756_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04433_, clk);
  dff _50757_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04522_, clk);
  dff _50758_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04613_, clk);
  dff _50759_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04706_, clk);
  dff _50760_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04792_, clk);
  dff _50761_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04876_, clk);
  dff _50762_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _25273_, clk);
  dff _50763_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _06083_, clk);
  dff _50764_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _06084_, clk);
  dff _50765_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _06085_, clk);
  dff _50766_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _06086_, clk);
  dff _50767_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _06087_, clk);
  dff _50768_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _06088_, clk);
  dff _50769_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _06089_, clk);
  dff _50770_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06079_, clk);
  dff _50771_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _06090_, clk);
  dff _50772_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _06091_, clk);
  dff _50773_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _06092_, clk);
  dff _50774_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _06093_, clk);
  dff _50775_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _06094_, clk);
  dff _50776_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _06096_, clk);
  dff _50777_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _06097_, clk);
  dff _50778_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _06080_, clk);
  dff _50779_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _06098_, clk);
  dff _50780_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _06099_, clk);
  dff _50781_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _06100_, clk);
  dff _50782_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _06101_, clk);
  dff _50783_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _06102_, clk);
  dff _50784_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _06103_, clk);
  dff _50785_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _06104_, clk);
  dff _50786_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _06081_, clk);
  dff _50787_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _05706_, clk);
  dff _50788_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _05707_, clk);
  dff _50789_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _05692_, clk);
  dff _50790_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _05708_, clk);
  dff _50791_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _05709_, clk);
  dff _50792_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05693_, clk);
  dff _50793_ (\oc8051_top_1.oc8051_decoder1.state [0], _05710_, clk);
  dff _50794_ (\oc8051_top_1.oc8051_decoder1.state [1], _05694_, clk);
  dff _50795_ (\oc8051_top_1.oc8051_decoder1.op [0], _05711_, clk);
  dff _50796_ (\oc8051_top_1.oc8051_decoder1.op [1], _05712_, clk);
  dff _50797_ (\oc8051_top_1.oc8051_decoder1.op [2], _05713_, clk);
  dff _50798_ (\oc8051_top_1.oc8051_decoder1.op [3], _05714_, clk);
  dff _50799_ (\oc8051_top_1.oc8051_decoder1.op [4], _05715_, clk);
  dff _50800_ (\oc8051_top_1.oc8051_decoder1.op [5], _05716_, clk);
  dff _50801_ (\oc8051_top_1.oc8051_decoder1.op [6], _05717_, clk);
  dff _50802_ (\oc8051_top_1.oc8051_decoder1.op [7], _05695_, clk);
  dff _50803_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _05696_, clk);
  dff _50804_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05951_, clk);
  dff _50805_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05697_, clk);
  dff _50806_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _05952_, clk);
  dff _50807_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05698_, clk);
  dff _50808_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05953_, clk);
  dff _50809_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05954_, clk);
  dff _50810_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05699_, clk);
  dff _50811_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _05955_, clk);
  dff _50812_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _05956_, clk);
  dff _50813_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05700_, clk);
  dff _50814_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _05957_, clk);
  dff _50815_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05701_, clk);
  dff _50816_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _05958_, clk);
  dff _50817_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _05959_, clk);
  dff _50818_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _05960_, clk);
  dff _50819_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _05702_, clk);
  dff _50820_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _05961_, clk);
  dff _50821_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05703_, clk);
  dff _50822_ (\oc8051_top_1.oc8051_decoder1.wr , _05705_, clk);
  dff _50823_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _06419_, clk);
  dff _50824_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _06438_, clk);
  dff _50825_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _06439_, clk);
  dff _50826_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _06440_, clk);
  dff _50827_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _06441_, clk);
  dff _50828_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _06442_, clk);
  dff _50829_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _06443_, clk);
  dff _50830_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _06444_, clk);
  dff _50831_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _06420_, clk);
  dff _50832_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _06445_, clk);
  dff _50833_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _06446_, clk);
  dff _50834_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _06447_, clk);
  dff _50835_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _06448_, clk);
  dff _50836_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _06449_, clk);
  dff _50837_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _06450_, clk);
  dff _50838_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _06451_, clk);
  dff _50839_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _06421_, clk);
  dff _50840_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _06452_, clk);
  dff _50841_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _06453_, clk);
  dff _50842_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _06454_, clk);
  dff _50843_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _06455_, clk);
  dff _50844_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _06456_, clk);
  dff _50845_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _06457_, clk);
  dff _50846_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _06458_, clk);
  dff _50847_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _06422_, clk);
  dff _50848_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _06459_, clk);
  dff _50849_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _06460_, clk);
  dff _50850_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _06461_, clk);
  dff _50851_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _06462_, clk);
  dff _50852_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _06463_, clk);
  dff _50853_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _06464_, clk);
  dff _50854_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _06465_, clk);
  dff _50855_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _06423_, clk);
  dff _50856_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _06466_, clk);
  dff _50857_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _06467_, clk);
  dff _50858_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _06468_, clk);
  dff _50859_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _06469_, clk);
  dff _50860_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _06470_, clk);
  dff _50861_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _06471_, clk);
  dff _50862_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _06472_, clk);
  dff _50863_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _06424_, clk);
  dff _50864_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _06473_, clk);
  dff _50865_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _06474_, clk);
  dff _50866_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _06475_, clk);
  dff _50867_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _06476_, clk);
  dff _50868_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _06477_, clk);
  dff _50869_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _06478_, clk);
  dff _50870_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _06479_, clk);
  dff _50871_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _06425_, clk);
  dff _50872_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _06480_, clk);
  dff _50873_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _06481_, clk);
  dff _50874_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _06482_, clk);
  dff _50875_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _06483_, clk);
  dff _50876_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _06484_, clk);
  dff _50877_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _06486_, clk);
  dff _50878_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _06487_, clk);
  dff _50879_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _06426_, clk);
  dff _50880_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _06488_, clk);
  dff _50881_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _06489_, clk);
  dff _50882_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _06490_, clk);
  dff _50883_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _06491_, clk);
  dff _50884_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _06492_, clk);
  dff _50885_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _06493_, clk);
  dff _50886_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _06494_, clk);
  dff _50887_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _06427_, clk);
  dff _50888_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _06200_, clk);
  dff _50889_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _06201_, clk);
  dff _50890_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _06202_, clk);
  dff _50891_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _06203_, clk);
  dff _50892_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _06114_, clk);
  dff _50893_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _06150_, clk);
  dff _50894_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _06151_, clk);
  dff _50895_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _06152_, clk);
  dff _50896_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06154_, clk);
  dff _50897_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _06155_, clk);
  dff _50898_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _06156_, clk);
  dff _50899_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _06157_, clk);
  dff _50900_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _06158_, clk);
  dff _50901_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _06159_, clk);
  dff _50902_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _06160_, clk);
  dff _50903_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _06161_, clk);
  dff _50904_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _06162_, clk);
  dff _50905_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _06163_, clk);
  dff _50906_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _06164_, clk);
  dff _50907_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _06165_, clk);
  dff _50908_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _06107_, clk);
  dff _50909_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _06166_, clk);
  dff _50910_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _06167_, clk);
  dff _50911_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _06168_, clk);
  dff _50912_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _06169_, clk);
  dff _50913_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _06170_, clk);
  dff _50914_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _06171_, clk);
  dff _50915_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _06172_, clk);
  dff _50916_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _06173_, clk);
  dff _50917_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _06174_, clk);
  dff _50918_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _06175_, clk);
  dff _50919_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _06176_, clk);
  dff _50920_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _06177_, clk);
  dff _50921_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _06178_, clk);
  dff _50922_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _06179_, clk);
  dff _50923_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _06180_, clk);
  dff _50924_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _06108_, clk);
  dff _50925_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _06204_, clk);
  dff _50926_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _06205_, clk);
  dff _50927_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _06206_, clk);
  dff _50928_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _06207_, clk);
  dff _50929_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _06208_, clk);
  dff _50930_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _06209_, clk);
  dff _50931_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _06210_, clk);
  dff _50932_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _06211_, clk);
  dff _50933_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _06212_, clk);
  dff _50934_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _06213_, clk);
  dff _50935_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _06214_, clk);
  dff _50936_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _06215_, clk);
  dff _50937_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _06216_, clk);
  dff _50938_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _06217_, clk);
  dff _50939_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _06218_, clk);
  dff _50940_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _06219_, clk);
  dff _50941_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _06220_, clk);
  dff _50942_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _06221_, clk);
  dff _50943_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _06222_, clk);
  dff _50944_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _06223_, clk);
  dff _50945_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _06224_, clk);
  dff _50946_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _06225_, clk);
  dff _50947_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _06226_, clk);
  dff _50948_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _06227_, clk);
  dff _50949_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _06228_, clk);
  dff _50950_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _06229_, clk);
  dff _50951_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _06230_, clk);
  dff _50952_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _06231_, clk);
  dff _50953_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _06232_, clk);
  dff _50954_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _06233_, clk);
  dff _50955_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _06234_, clk);
  dff _50956_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _06136_, clk);
  dff _50957_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _06113_, clk);
  dff _50958_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _50959_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _06235_, clk);
  dff _50960_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _06236_, clk);
  dff _50961_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _06237_, clk);
  dff _50962_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _06238_, clk);
  dff _50963_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _06239_, clk);
  dff _50964_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _06240_, clk);
  dff _50965_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _06241_, clk);
  dff _50966_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _06115_, clk);
  dff _50967_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _06242_, clk);
  dff _50968_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _06243_, clk);
  dff _50969_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _06244_, clk);
  dff _50970_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _06245_, clk);
  dff _50971_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _06246_, clk);
  dff _50972_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _06247_, clk);
  dff _50973_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _06248_, clk);
  dff _50974_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _06116_, clk);
  dff _50975_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _06249_, clk);
  dff _50976_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _06250_, clk);
  dff _50977_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _06251_, clk);
  dff _50978_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _06252_, clk);
  dff _50979_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _06253_, clk);
  dff _50980_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _06254_, clk);
  dff _50981_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _06255_, clk);
  dff _50982_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _06117_, clk);
  dff _50983_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _06118_, clk);
  dff _50984_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _06119_, clk);
  dff _50985_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _06256_, clk);
  dff _50986_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _06258_, clk);
  dff _50987_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _06259_, clk);
  dff _50988_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _06260_, clk);
  dff _50989_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _06261_, clk);
  dff _50990_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _06262_, clk);
  dff _50991_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _06263_, clk);
  dff _50992_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _06120_, clk);
  dff _50993_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _06264_, clk);
  dff _50994_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _06265_, clk);
  dff _50995_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _06266_, clk);
  dff _50996_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _06267_, clk);
  dff _50997_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _06268_, clk);
  dff _50998_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _06269_, clk);
  dff _50999_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _06270_, clk);
  dff _51000_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _06271_, clk);
  dff _51001_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _06272_, clk);
  dff _51002_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _06273_, clk);
  dff _51003_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _06274_, clk);
  dff _51004_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _06275_, clk);
  dff _51005_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _06276_, clk);
  dff _51006_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _06277_, clk);
  dff _51007_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _06278_, clk);
  dff _51008_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _06121_, clk);
  dff _51009_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _06279_, clk);
  dff _51010_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _06280_, clk);
  dff _51011_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _06281_, clk);
  dff _51012_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _06282_, clk);
  dff _51013_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _06283_, clk);
  dff _51014_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _06284_, clk);
  dff _51015_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _06285_, clk);
  dff _51016_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _06286_, clk);
  dff _51017_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _06287_, clk);
  dff _51018_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _06288_, clk);
  dff _51019_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _06289_, clk);
  dff _51020_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _06290_, clk);
  dff _51021_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _06291_, clk);
  dff _51022_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _06292_, clk);
  dff _51023_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _06293_, clk);
  dff _51024_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _06122_, clk);
  dff _51025_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _06123_, clk);
  dff _51026_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _06125_, clk);
  dff _51027_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _06124_, clk);
  dff _51028_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _06294_, clk);
  dff _51029_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _06295_, clk);
  dff _51030_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06296_, clk);
  dff _51031_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _06297_, clk);
  dff _51032_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _06298_, clk);
  dff _51033_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _06299_, clk);
  dff _51034_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _06300_, clk);
  dff _51035_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _06126_, clk);
  dff _51036_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _06301_, clk);
  dff _51037_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _06302_, clk);
  dff _51038_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _06127_, clk);
  dff _51039_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _06303_, clk);
  dff _51040_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _06304_, clk);
  dff _51041_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _06305_, clk);
  dff _51042_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _06306_, clk);
  dff _51043_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _06307_, clk);
  dff _51044_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _06308_, clk);
  dff _51045_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _06309_, clk);
  dff _51046_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _06128_, clk);
  dff _51047_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _06310_, clk);
  dff _51048_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _06311_, clk);
  dff _51049_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _06312_, clk);
  dff _51050_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _06313_, clk);
  dff _51051_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _06314_, clk);
  dff _51052_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _06315_, clk);
  dff _51053_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _06316_, clk);
  dff _51054_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _06129_, clk);
  dff _51055_ (\oc8051_top_1.oc8051_memory_interface1.reti , _06130_, clk);
  dff _51056_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _06317_, clk);
  dff _51057_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _06318_, clk);
  dff _51058_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _06319_, clk);
  dff _51059_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _06320_, clk);
  dff _51060_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _06321_, clk);
  dff _51061_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _06322_, clk);
  dff _51062_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _06323_, clk);
  dff _51063_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _06131_, clk);
  dff _51064_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _06132_, clk);
  dff _51065_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _06134_, clk);
  dff _51066_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _06324_, clk);
  dff _51067_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _06325_, clk);
  dff _51068_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _06326_, clk);
  dff _51069_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _06135_, clk);
  dff _51070_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _06327_, clk);
  dff _51071_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _06328_, clk);
  dff _51072_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _06329_, clk);
  dff _51073_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _06330_, clk);
  dff _51074_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _06331_, clk);
  dff _51075_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _06332_, clk);
  dff _51076_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _06333_, clk);
  dff _51077_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _06334_, clk);
  dff _51078_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _06335_, clk);
  dff _51079_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _06336_, clk);
  dff _51080_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _06337_, clk);
  dff _51081_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _06338_, clk);
  dff _51082_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _06339_, clk);
  dff _51083_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _06340_, clk);
  dff _51084_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _06341_, clk);
  dff _51085_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _06342_, clk);
  dff _51086_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _06343_, clk);
  dff _51087_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _06344_, clk);
  dff _51088_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _06345_, clk);
  dff _51089_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _06346_, clk);
  dff _51090_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _06347_, clk);
  dff _51091_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _06348_, clk);
  dff _51092_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _06349_, clk);
  dff _51093_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _06350_, clk);
  dff _51094_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _06351_, clk);
  dff _51095_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _06352_, clk);
  dff _51096_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _06353_, clk);
  dff _51097_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _06354_, clk);
  dff _51098_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _06355_, clk);
  dff _51099_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _06356_, clk);
  dff _51100_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _06357_, clk);
  dff _51101_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _06137_, clk);
  dff _51102_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _06359_, clk);
  dff _51103_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _06360_, clk);
  dff _51104_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _06361_, clk);
  dff _51105_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _06362_, clk);
  dff _51106_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _06363_, clk);
  dff _51107_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _06364_, clk);
  dff _51108_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _06365_, clk);
  dff _51109_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _06138_, clk);
  dff _51110_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _06139_, clk);
  dff _51111_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _06140_, clk);
  dff _51112_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _06366_, clk);
  dff _51113_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _06367_, clk);
  dff _51114_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _06368_, clk);
  dff _51115_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _06369_, clk);
  dff _51116_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _06370_, clk);
  dff _51117_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _06371_, clk);
  dff _51118_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _06372_, clk);
  dff _51119_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _06373_, clk);
  dff _51120_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _06374_, clk);
  dff _51121_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _06375_, clk);
  dff _51122_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _06376_, clk);
  dff _51123_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _06377_, clk);
  dff _51124_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _06378_, clk);
  dff _51125_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _06379_, clk);
  dff _51126_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _06380_, clk);
  dff _51127_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _06141_, clk);
  dff _51128_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _06142_, clk);
  dff _51129_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _06143_, clk);
  dff _51130_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _06144_, clk);
  dff _51131_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _06381_, clk);
  dff _51132_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _06382_, clk);
  dff _51133_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _06383_, clk);
  dff _51134_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _06384_, clk);
  dff _51135_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _06385_, clk);
  dff _51136_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _06386_, clk);
  dff _51137_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _06387_, clk);
  dff _51138_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _06388_, clk);
  dff _51139_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _06389_, clk);
  dff _51140_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _06390_, clk);
  dff _51141_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _06391_, clk);
  dff _51142_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _06392_, clk);
  dff _51143_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _06393_, clk);
  dff _51144_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _06394_, clk);
  dff _51145_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _06395_, clk);
  dff _51146_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _06145_, clk);
  dff _51147_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _06146_, clk);
  dff _51148_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _06533_, clk);
  dff _51149_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _06538_, clk);
  dff _51150_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _06539_, clk);
  dff _51151_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _06540_, clk);
  dff _51152_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _06541_, clk);
  dff _51153_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _06542_, clk);
  dff _51154_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _06543_, clk);
  dff _51155_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _06544_, clk);
  dff _51156_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _06534_, clk);
  dff _51157_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _06535_, clk);
  dff _51158_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _06545_, clk);
  dff _51159_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _06546_, clk);
  dff _51160_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _06536_, clk);
  dff _51161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _12202_, clk);
  dff _51162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _12204_, clk);
  dff _51163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _12205_, clk);
  dff _51164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _12207_, clk);
  dff _51165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _12208_, clk);
  dff _51166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _12210_, clk);
  dff _51167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _12211_, clk);
  dff _51168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _12213_, clk);
  dff _51169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _12214_, clk);
  dff _51170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _12215_, clk);
  dff _51171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _12216_, clk);
  dff _51172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _12217_, clk);
  dff _51173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _12219_, clk);
  dff _51174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _12220_, clk);
  dff _51175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _12221_, clk);
  dff _51176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _12222_, clk);
  dff _51177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _12282_, clk);
  dff _51178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _12283_, clk);
  dff _51179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _12284_, clk);
  dff _51180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _12286_, clk);
  dff _51181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _12287_, clk);
  dff _51182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _12288_, clk);
  dff _51183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _12290_, clk);
  dff _51184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _12291_, clk);
  dff _51185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _12272_, clk);
  dff _51186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _12273_, clk);
  dff _51187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _12275_, clk);
  dff _51188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _12276_, clk);
  dff _51189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _12277_, clk);
  dff _51190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _12279_, clk);
  dff _51191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _12280_, clk);
  dff _51192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _12281_, clk);
  dff _51193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _12263_, clk);
  dff _51194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _12264_, clk);
  dff _51195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _12265_, clk);
  dff _51196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _12266_, clk);
  dff _51197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _12268_, clk);
  dff _51198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _12269_, clk);
  dff _51199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _12270_, clk);
  dff _51200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _12271_, clk);
  dff _51201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _12253_, clk);
  dff _51202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _12254_, clk);
  dff _51203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _12256_, clk);
  dff _51204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _12257_, clk);
  dff _51205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _12258_, clk);
  dff _51206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _12259_, clk);
  dff _51207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _12260_, clk);
  dff _51208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _12261_, clk);
  dff _51209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _12244_, clk);
  dff _51210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _12245_, clk);
  dff _51211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _12246_, clk);
  dff _51212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _12247_, clk);
  dff _51213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _12248_, clk);
  dff _51214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _12249_, clk);
  dff _51215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _12250_, clk);
  dff _51216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _12252_, clk);
  dff _51217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _12234_, clk);
  dff _51218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _12235_, clk);
  dff _51219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _12236_, clk);
  dff _51220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _12237_, clk);
  dff _51221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _12238_, clk);
  dff _51222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _12239_, clk);
  dff _51223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _12241_, clk);
  dff _51224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _12242_, clk);
  dff _51225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _12224_, clk);
  dff _51226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _12225_, clk);
  dff _51227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _12226_, clk);
  dff _51228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _12227_, clk);
  dff _51229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _12228_, clk);
  dff _51230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _12230_, clk);
  dff _51231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _12231_, clk);
  dff _51232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _12232_, clk);
  dff _51233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _13995_, clk);
  dff _51234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _13996_, clk);
  dff _51235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _13998_, clk);
  dff _51236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _13999_, clk);
  dff _51237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _14000_, clk);
  dff _51238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _14001_, clk);
  dff _51239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _14003_, clk);
  dff _51240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _14004_, clk);
  dff _51241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _13986_, clk);
  dff _51242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _13987_, clk);
  dff _51243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _13988_, clk);
  dff _51244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _13989_, clk);
  dff _51245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _13991_, clk);
  dff _51246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _13992_, clk);
  dff _51247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _13993_, clk);
  dff _51248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _13994_, clk);
  dff _51249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _13976_, clk);
  dff _51250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _13977_, clk);
  dff _51251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _13979_, clk);
  dff _51252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _13980_, clk);
  dff _51253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _13981_, clk);
  dff _51254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _13982_, clk);
  dff _51255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _13983_, clk);
  dff _51256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _13984_, clk);
  dff _51257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _13966_, clk);
  dff _51258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _13967_, clk);
  dff _51259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _13968_, clk);
  dff _51260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _13970_, clk);
  dff _51261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _13971_, clk);
  dff _51262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _13972_, clk);
  dff _51263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _13974_, clk);
  dff _51264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _13975_, clk);
  dff _51265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _13956_, clk);
  dff _51266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _13958_, clk);
  dff _51267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _13959_, clk);
  dff _51268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _13960_, clk);
  dff _51269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _13961_, clk);
  dff _51270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _13962_, clk);
  dff _51271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _13963_, clk);
  dff _51272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _13964_, clk);
  dff _51273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _13947_, clk);
  dff _51274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _13948_, clk);
  dff _51275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _13949_, clk);
  dff _51276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _13950_, clk);
  dff _51277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _13951_, clk);
  dff _51278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _13952_, clk);
  dff _51279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _13954_, clk);
  dff _51280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _13955_, clk);
  dff _51281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _13927_, clk);
  dff _51282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _13928_, clk);
  dff _51283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _13930_, clk);
  dff _51284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _13931_, clk);
  dff _51285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _13932_, clk);
  dff _51286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _13934_, clk);
  dff _51287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _13935_, clk);
  dff _51288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _13936_, clk);
  dff _51289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _13899_, clk);
  dff _51290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _13900_, clk);
  dff _51291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _13901_, clk);
  dff _51292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _13902_, clk);
  dff _51293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _13903_, clk);
  dff _51294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _13904_, clk);
  dff _51295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _13906_, clk);
  dff _51296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _13907_, clk);
  dff _51297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _13879_, clk);
  dff _51298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _13880_, clk);
  dff _51299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _13882_, clk);
  dff _51300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _13883_, clk);
  dff _51301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _13884_, clk);
  dff _51302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _13886_, clk);
  dff _51303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _13887_, clk);
  dff _51304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _13888_, clk);
  dff _51305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _13859_, clk);
  dff _51306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _13861_, clk);
  dff _51307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _13862_, clk);
  dff _51308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _13863_, clk);
  dff _51309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _13864_, clk);
  dff _51310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _13866_, clk);
  dff _51311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _13867_, clk);
  dff _51312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _13868_, clk);
  dff _51313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _13840_, clk);
  dff _51314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _13842_, clk);
  dff _51315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _13843_, clk);
  dff _51316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _13844_, clk);
  dff _51317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _13845_, clk);
  dff _51318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _13846_, clk);
  dff _51319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _13847_, clk);
  dff _51320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _13848_, clk);
  dff _51321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _13821_, clk);
  dff _51322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _13822_, clk);
  dff _51323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _13823_, clk);
  dff _51324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _13825_, clk);
  dff _51325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _13826_, clk);
  dff _51326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _13827_, clk);
  dff _51327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _13828_, clk);
  dff _51328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _13830_, clk);
  dff _51329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _13802_, clk);
  dff _51330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _13803_, clk);
  dff _51331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _13804_, clk);
  dff _51332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _13806_, clk);
  dff _51333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _13807_, clk);
  dff _51334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _13808_, clk);
  dff _51335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _13809_, clk);
  dff _51336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _13810_, clk);
  dff _51337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _13783_, clk);
  dff _51338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _13784_, clk);
  dff _51339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _13785_, clk);
  dff _51340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _13786_, clk);
  dff _51341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _13787_, clk);
  dff _51342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _13789_, clk);
  dff _51343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _13790_, clk);
  dff _51344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _13791_, clk);
  dff _51345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _13763_, clk);
  dff _51346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _13765_, clk);
  dff _51347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _13766_, clk);
  dff _51348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _13767_, clk);
  dff _51349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _13768_, clk);
  dff _51350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _13770_, clk);
  dff _51351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _13771_, clk);
  dff _51352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _13772_, clk);
  dff _51353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _13743_, clk);
  dff _51354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _13745_, clk);
  dff _51355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _13746_, clk);
  dff _51356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _13747_, clk);
  dff _51357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _13749_, clk);
  dff _51358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _13750_, clk);
  dff _51359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _13751_, clk);
  dff _51360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _13752_, clk);
  dff _51361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _13725_, clk);
  dff _51362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _13726_, clk);
  dff _51363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _13727_, clk);
  dff _51364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _13728_, clk);
  dff _51365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _13729_, clk);
  dff _51366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _13730_, clk);
  dff _51367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _13731_, clk);
  dff _51368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _13733_, clk);
  dff _51369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _13705_, clk);
  dff _51370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _13706_, clk);
  dff _51371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _13707_, clk);
  dff _51372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _13709_, clk);
  dff _51373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _13710_, clk);
  dff _51374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _13711_, clk);
  dff _51375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _13713_, clk);
  dff _51376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _13714_, clk);
  dff _51377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _13695_, clk);
  dff _51378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _13697_, clk);
  dff _51379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _13698_, clk);
  dff _51380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _13699_, clk);
  dff _51381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _13701_, clk);
  dff _51382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _13702_, clk);
  dff _51383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _13703_, clk);
  dff _51384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _13704_, clk);
  dff _51385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _13686_, clk);
  dff _51386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _13687_, clk);
  dff _51387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _13689_, clk);
  dff _51388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _13690_, clk);
  dff _51389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _13691_, clk);
  dff _51390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _13692_, clk);
  dff _51391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _13693_, clk);
  dff _51392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _13694_, clk);
  dff _51393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _13677_, clk);
  dff _51394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _13678_, clk);
  dff _51395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _13679_, clk);
  dff _51396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _13680_, clk);
  dff _51397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _13681_, clk);
  dff _51398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _13682_, clk);
  dff _51399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _13683_, clk);
  dff _51400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _13685_, clk);
  dff _51401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _13657_, clk);
  dff _51402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _13658_, clk);
  dff _51403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _13659_, clk);
  dff _51404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _13661_, clk);
  dff _51405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _13662_, clk);
  dff _51406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _13663_, clk);
  dff _51407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _13665_, clk);
  dff _51408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _13666_, clk);
  dff _51409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _13637_, clk);
  dff _51410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _13638_, clk);
  dff _51411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _13640_, clk);
  dff _51412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _13641_, clk);
  dff _51413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _13642_, clk);
  dff _51414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _13643_, clk);
  dff _51415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _13644_, clk);
  dff _51416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _13645_, clk);
  dff _51417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _13608_, clk);
  dff _51418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _13609_, clk);
  dff _51419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _13610_, clk);
  dff _51420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _13612_, clk);
  dff _51421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _13613_, clk);
  dff _51422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _13614_, clk);
  dff _51423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _13616_, clk);
  dff _51424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _13617_, clk);
  dff _51425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _13598_, clk);
  dff _51426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _13600_, clk);
  dff _51427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _13601_, clk);
  dff _51428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _13602_, clk);
  dff _51429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _13604_, clk);
  dff _51430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _13605_, clk);
  dff _51431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _13606_, clk);
  dff _51432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _13607_, clk);
  dff _51433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _13589_, clk);
  dff _51434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _13590_, clk);
  dff _51435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _13591_, clk);
  dff _51436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _13593_, clk);
  dff _51437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _13594_, clk);
  dff _51438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _13595_, clk);
  dff _51439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _13596_, clk);
  dff _51440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _13597_, clk);
  dff _51441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _13579_, clk);
  dff _51442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _13581_, clk);
  dff _51443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _13582_, clk);
  dff _51444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _13583_, clk);
  dff _51445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _13584_, clk);
  dff _51446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _13585_, clk);
  dff _51447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _13586_, clk);
  dff _51448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _13587_, clk);
  dff _51449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _13570_, clk);
  dff _51450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _13571_, clk);
  dff _51451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _13572_, clk);
  dff _51452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _13573_, clk);
  dff _51453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _13574_, clk);
  dff _51454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _13576_, clk);
  dff _51455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _13577_, clk);
  dff _51456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _13578_, clk);
  dff _51457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _13560_, clk);
  dff _51458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _13561_, clk);
  dff _51459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _13562_, clk);
  dff _51460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _13564_, clk);
  dff _51461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _13565_, clk);
  dff _51462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _13566_, clk);
  dff _51463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _13567_, clk);
  dff _51464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _13569_, clk);
  dff _51465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _13550_, clk);
  dff _51466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _13552_, clk);
  dff _51467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _13553_, clk);
  dff _51468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _13554_, clk);
  dff _51469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _13555_, clk);
  dff _51470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _13557_, clk);
  dff _51471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _13558_, clk);
  dff _51472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _13559_, clk);
  dff _51473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _13540_, clk);
  dff _51474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _13541_, clk);
  dff _51475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _13542_, clk);
  dff _51476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _13544_, clk);
  dff _51477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _13545_, clk);
  dff _51478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _13546_, clk);
  dff _51479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _13548_, clk);
  dff _51480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _13549_, clk);
  dff _51481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _13530_, clk);
  dff _51482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _13532_, clk);
  dff _51483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _13533_, clk);
  dff _51484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _13534_, clk);
  dff _51485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _13536_, clk);
  dff _51486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _13537_, clk);
  dff _51487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _13538_, clk);
  dff _51488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _13539_, clk);
  dff _51489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _13521_, clk);
  dff _51490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _13522_, clk);
  dff _51491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _13524_, clk);
  dff _51492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _13525_, clk);
  dff _51493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _13526_, clk);
  dff _51494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _13527_, clk);
  dff _51495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _13528_, clk);
  dff _51496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _13529_, clk);
  dff _51497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _13512_, clk);
  dff _51498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _13513_, clk);
  dff _51499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _13514_, clk);
  dff _51500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _13515_, clk);
  dff _51501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _13516_, clk);
  dff _51502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _13517_, clk);
  dff _51503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _13518_, clk);
  dff _51504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _13520_, clk);
  dff _51505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _13502_, clk);
  dff _51506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _13503_, clk);
  dff _51507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _13504_, clk);
  dff _51508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _13505_, clk);
  dff _51509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _13506_, clk);
  dff _51510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _13508_, clk);
  dff _51511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _13509_, clk);
  dff _51512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _13510_, clk);
  dff _51513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _13492_, clk);
  dff _51514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _13493_, clk);
  dff _51515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _13494_, clk);
  dff _51516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _13496_, clk);
  dff _51517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _13497_, clk);
  dff _51518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _13498_, clk);
  dff _51519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _13500_, clk);
  dff _51520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _13501_, clk);
  dff _51521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _13482_, clk);
  dff _51522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _13484_, clk);
  dff _51523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _13485_, clk);
  dff _51524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _13486_, clk);
  dff _51525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _13488_, clk);
  dff _51526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _13489_, clk);
  dff _51527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _13490_, clk);
  dff _51528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _13491_, clk);
  dff _51529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _12292_, clk);
  dff _51530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _12293_, clk);
  dff _51531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _12294_, clk);
  dff _51532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _12295_, clk);
  dff _51533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _12297_, clk);
  dff _51534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _12298_, clk);
  dff _51535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _12299_, clk);
  dff _51536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _12300_, clk);
  dff _51537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _13473_, clk);
  dff _51538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _13474_, clk);
  dff _51539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _13476_, clk);
  dff _51540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _13477_, clk);
  dff _51541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _13478_, clk);
  dff _51542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _13479_, clk);
  dff _51543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _13480_, clk);
  dff _51544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _13481_, clk);
  dff _51545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _13464_, clk);
  dff _51546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _13465_, clk);
  dff _51547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _13466_, clk);
  dff _51548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _13467_, clk);
  dff _51549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _13468_, clk);
  dff _51550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _13469_, clk);
  dff _51551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _13470_, clk);
  dff _51552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _13472_, clk);
  dff _51553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _13454_, clk);
  dff _51554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _13455_, clk);
  dff _51555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _13456_, clk);
  dff _51556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _13457_, clk);
  dff _51557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _13458_, clk);
  dff _51558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _13460_, clk);
  dff _51559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _13461_, clk);
  dff _51560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _13462_, clk);
  dff _51561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _13444_, clk);
  dff _51562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _13445_, clk);
  dff _51563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _13446_, clk);
  dff _51564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _13448_, clk);
  dff _51565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _13449_, clk);
  dff _51566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _13450_, clk);
  dff _51567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _13452_, clk);
  dff _51568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _13453_, clk);
  dff _51569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _13434_, clk);
  dff _51570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _13435_, clk);
  dff _51571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _13436_, clk);
  dff _51572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _13437_, clk);
  dff _51573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _13438_, clk);
  dff _51574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _13439_, clk);
  dff _51575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _13441_, clk);
  dff _51576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _13442_, clk);
  dff _51577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _13424_, clk);
  dff _51578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _13425_, clk);
  dff _51579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _13426_, clk);
  dff _51580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _13427_, clk);
  dff _51581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _13429_, clk);
  dff _51582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _13430_, clk);
  dff _51583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _13431_, clk);
  dff _51584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _13433_, clk);
  dff _51585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _13414_, clk);
  dff _51586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _13415_, clk);
  dff _51587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _13417_, clk);
  dff _51588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _13418_, clk);
  dff _51589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _13419_, clk);
  dff _51590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _13421_, clk);
  dff _51591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _13422_, clk);
  dff _51592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _13423_, clk);
  dff _51593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _13405_, clk);
  dff _51594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _13406_, clk);
  dff _51595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _13407_, clk);
  dff _51596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _13409_, clk);
  dff _51597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _13410_, clk);
  dff _51598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _13411_, clk);
  dff _51599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _13412_, clk);
  dff _51600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _13413_, clk);
  dff _51601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _13395_, clk);
  dff _51602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _13397_, clk);
  dff _51603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _13398_, clk);
  dff _51604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _13399_, clk);
  dff _51605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _13400_, clk);
  dff _51606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _13401_, clk);
  dff _51607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _13402_, clk);
  dff _51608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _13403_, clk);
  dff _51609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _13386_, clk);
  dff _51610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _13387_, clk);
  dff _51611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _13388_, clk);
  dff _51612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _13389_, clk);
  dff _51613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _13390_, clk);
  dff _51614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _13391_, clk);
  dff _51615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _13393_, clk);
  dff _51616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _13394_, clk);
  dff _51617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _13376_, clk);
  dff _51618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _13377_, clk);
  dff _51619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _13378_, clk);
  dff _51620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _13379_, clk);
  dff _51621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _13381_, clk);
  dff _51622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _13382_, clk);
  dff _51623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _13383_, clk);
  dff _51624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _13385_, clk);
  dff _51625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _13366_, clk);
  dff _51626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _13367_, clk);
  dff _51627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _13369_, clk);
  dff _51628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _13370_, clk);
  dff _51629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _13371_, clk);
  dff _51630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _13373_, clk);
  dff _51631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _13374_, clk);
  dff _51632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _13375_, clk);
  dff _51633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _13357_, clk);
  dff _51634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _13358_, clk);
  dff _51635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _13359_, clk);
  dff _51636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _13361_, clk);
  dff _51637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _13362_, clk);
  dff _51638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _13363_, clk);
  dff _51639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _13364_, clk);
  dff _51640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _13365_, clk);
  dff _51641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _13347_, clk);
  dff _51642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _13349_, clk);
  dff _51643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _13350_, clk);
  dff _51644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _13351_, clk);
  dff _51645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _13352_, clk);
  dff _51646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _13353_, clk);
  dff _51647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _13354_, clk);
  dff _51648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _13355_, clk);
  dff _51649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _13337_, clk);
  dff _51650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _13338_, clk);
  dff _51651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _13340_, clk);
  dff _51652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _13341_, clk);
  dff _51653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _13342_, clk);
  dff _51654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _13343_, clk);
  dff _51655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _13345_, clk);
  dff _51656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _13346_, clk);
  dff _51657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _13328_, clk);
  dff _51658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _13329_, clk);
  dff _51659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _13330_, clk);
  dff _51660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _13331_, clk);
  dff _51661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _13332_, clk);
  dff _51662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _13333_, clk);
  dff _51663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _13334_, clk);
  dff _51664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _13336_, clk);
  dff _51665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _13318_, clk);
  dff _51666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _13319_, clk);
  dff _51667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _13320_, clk);
  dff _51668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _13321_, clk);
  dff _51669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _13322_, clk);
  dff _51670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _13324_, clk);
  dff _51671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _13325_, clk);
  dff _51672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _13326_, clk);
  dff _51673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _13308_, clk);
  dff _51674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _13309_, clk);
  dff _51675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _13310_, clk);
  dff _51676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _13312_, clk);
  dff _51677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _13313_, clk);
  dff _51678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _13314_, clk);
  dff _51679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _13316_, clk);
  dff _51680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _13317_, clk);
  dff _51681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _13298_, clk);
  dff _51682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _13300_, clk);
  dff _51683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _13301_, clk);
  dff _51684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _13302_, clk);
  dff _51685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _13304_, clk);
  dff _51686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _13305_, clk);
  dff _51687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _13306_, clk);
  dff _51688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _13307_, clk);
  dff _51689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _13289_, clk);
  dff _51690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _13290_, clk);
  dff _51691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _13292_, clk);
  dff _51692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _13293_, clk);
  dff _51693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _13294_, clk);
  dff _51694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _13295_, clk);
  dff _51695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _13296_, clk);
  dff _51696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _13297_, clk);
  dff _51697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _13279_, clk);
  dff _51698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _13281_, clk);
  dff _51699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _13282_, clk);
  dff _51700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _13283_, clk);
  dff _51701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _13284_, clk);
  dff _51702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _13285_, clk);
  dff _51703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _13286_, clk);
  dff _51704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _13287_, clk);
  dff _51705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _13270_, clk);
  dff _51706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _13271_, clk);
  dff _51707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _13272_, clk);
  dff _51708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _13273_, clk);
  dff _51709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _13274_, clk);
  dff _51710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _13276_, clk);
  dff _51711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _13277_, clk);
  dff _51712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _13278_, clk);
  dff _51713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _13260_, clk);
  dff _51714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _13261_, clk);
  dff _51715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _13262_, clk);
  dff _51716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _13264_, clk);
  dff _51717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _13265_, clk);
  dff _51718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _13266_, clk);
  dff _51719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _13267_, clk);
  dff _51720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _13269_, clk);
  dff _51721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _13250_, clk);
  dff _51722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _13252_, clk);
  dff _51723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _13253_, clk);
  dff _51724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _13254_, clk);
  dff _51725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _13255_, clk);
  dff _51726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _13257_, clk);
  dff _51727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _13258_, clk);
  dff _51728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _13259_, clk);
  dff _51729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _13241_, clk);
  dff _51730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _13242_, clk);
  dff _51731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _13243_, clk);
  dff _51732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _13245_, clk);
  dff _51733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _13246_, clk);
  dff _51734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _13247_, clk);
  dff _51735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _13248_, clk);
  dff _51736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _13249_, clk);
  dff _51737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _13230_, clk);
  dff _51738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _13232_, clk);
  dff _51739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _13233_, clk);
  dff _51740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _13234_, clk);
  dff _51741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _13236_, clk);
  dff _51742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _13237_, clk);
  dff _51743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _13238_, clk);
  dff _51744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _13239_, clk);
  dff _51745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _13221_, clk);
  dff _51746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _13222_, clk);
  dff _51747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _13224_, clk);
  dff _51748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _13225_, clk);
  dff _51749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _13226_, clk);
  dff _51750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _13227_, clk);
  dff _51751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _13228_, clk);
  dff _51752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _13229_, clk);
  dff _51753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _13212_, clk);
  dff _51754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _13213_, clk);
  dff _51755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _13214_, clk);
  dff _51756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _13215_, clk);
  dff _51757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _13216_, clk);
  dff _51758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _13217_, clk);
  dff _51759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _13218_, clk);
  dff _51760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _13220_, clk);
  dff _51761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _13202_, clk);
  dff _51762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _13203_, clk);
  dff _51763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _13204_, clk);
  dff _51764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _13205_, clk);
  dff _51765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _13206_, clk);
  dff _51766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _13208_, clk);
  dff _51767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _13209_, clk);
  dff _51768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _13210_, clk);
  dff _51769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _13192_, clk);
  dff _51770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _13193_, clk);
  dff _51771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _13194_, clk);
  dff _51772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _13196_, clk);
  dff _51773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _13197_, clk);
  dff _51774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _13198_, clk);
  dff _51775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _13200_, clk);
  dff _51776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _13201_, clk);
  dff _51777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _13182_, clk);
  dff _51778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _13184_, clk);
  dff _51779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _13185_, clk);
  dff _51780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _13186_, clk);
  dff _51781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _13188_, clk);
  dff _51782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _13189_, clk);
  dff _51783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _13190_, clk);
  dff _51784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _13191_, clk);
  dff _51785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _13173_, clk);
  dff _51786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _13174_, clk);
  dff _51787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _13176_, clk);
  dff _51788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _13177_, clk);
  dff _51789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _13178_, clk);
  dff _51790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _13179_, clk);
  dff _51791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _13180_, clk);
  dff _51792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _13181_, clk);
  dff _51793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _13164_, clk);
  dff _51794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _13165_, clk);
  dff _51795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _13166_, clk);
  dff _51796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _13167_, clk);
  dff _51797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _13168_, clk);
  dff _51798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _13169_, clk);
  dff _51799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _13170_, clk);
  dff _51800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _13172_, clk);
  dff _51801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _13154_, clk);
  dff _51802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _13155_, clk);
  dff _51803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _13156_, clk);
  dff _51804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _13157_, clk);
  dff _51805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _13158_, clk);
  dff _51806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _13160_, clk);
  dff _51807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _13161_, clk);
  dff _51808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _13162_, clk);
  dff _51809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _13144_, clk);
  dff _51810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _13145_, clk);
  dff _51811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _13146_, clk);
  dff _51812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _13148_, clk);
  dff _51813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _13149_, clk);
  dff _51814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _13150_, clk);
  dff _51815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _13152_, clk);
  dff _51816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _13153_, clk);
  dff _51817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _13134_, clk);
  dff _51818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _13136_, clk);
  dff _51819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _13137_, clk);
  dff _51820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _13138_, clk);
  dff _51821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _13140_, clk);
  dff _51822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _13141_, clk);
  dff _51823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _13142_, clk);
  dff _51824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _13143_, clk);
  dff _51825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _13115_, clk);
  dff _51826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _13116_, clk);
  dff _51827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _13117_, clk);
  dff _51828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _13118_, clk);
  dff _51829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _13120_, clk);
  dff _51830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _13121_, clk);
  dff _51831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _13122_, clk);
  dff _51832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _13123_, clk);
  dff _51833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _13105_, clk);
  dff _51834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _13106_, clk);
  dff _51835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _13108_, clk);
  dff _51836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _13109_, clk);
  dff _51837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _13110_, clk);
  dff _51838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _13111_, clk);
  dff _51839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _13112_, clk);
  dff _51840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _13113_, clk);
  dff _51841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _13096_, clk);
  dff _51842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _13097_, clk);
  dff _51843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _13098_, clk);
  dff _51844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _13099_, clk);
  dff _51845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _13100_, clk);
  dff _51846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _13101_, clk);
  dff _51847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _13103_, clk);
  dff _51848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _13104_, clk);
  dff _51849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _13086_, clk);
  dff _51850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _13087_, clk);
  dff _51851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _13088_, clk);
  dff _51852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _13089_, clk);
  dff _51853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _13091_, clk);
  dff _51854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _13092_, clk);
  dff _51855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _13093_, clk);
  dff _51856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _13094_, clk);
  dff _51857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _13076_, clk);
  dff _51858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _13077_, clk);
  dff _51859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _13079_, clk);
  dff _51860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _13080_, clk);
  dff _51861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _13081_, clk);
  dff _51862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _13082_, clk);
  dff _51863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _13084_, clk);
  dff _51864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _13085_, clk);
  dff _51865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _13067_, clk);
  dff _51866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _13068_, clk);
  dff _51867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _13069_, clk);
  dff _51868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _13070_, clk);
  dff _51869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _13072_, clk);
  dff _51870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _13073_, clk);
  dff _51871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _13074_, clk);
  dff _51872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _13075_, clk);
  dff _51873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _13057_, clk);
  dff _51874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _13058_, clk);
  dff _51875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _13060_, clk);
  dff _51876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _13061_, clk);
  dff _51877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _13062_, clk);
  dff _51878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _13063_, clk);
  dff _51879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _13064_, clk);
  dff _51880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _13065_, clk);
  dff _51881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _13048_, clk);
  dff _51882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _13049_, clk);
  dff _51883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _13050_, clk);
  dff _51884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _13051_, clk);
  dff _51885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _13052_, clk);
  dff _51886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _13053_, clk);
  dff _51887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _13055_, clk);
  dff _51888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _13056_, clk);
  dff _51889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _13038_, clk);
  dff _51890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _13039_, clk);
  dff _51891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _13040_, clk);
  dff _51892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _13041_, clk);
  dff _51893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _13043_, clk);
  dff _51894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _13044_, clk);
  dff _51895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _13045_, clk);
  dff _51896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _13046_, clk);
  dff _51897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _13028_, clk);
  dff _51898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _13029_, clk);
  dff _51899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _13031_, clk);
  dff _51900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _13032_, clk);
  dff _51901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _13033_, clk);
  dff _51902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _13034_, clk);
  dff _51903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _13036_, clk);
  dff _51904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _13037_, clk);
  dff _51905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _13018_, clk);
  dff _51906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _13019_, clk);
  dff _51907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _13020_, clk);
  dff _51908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _13021_, clk);
  dff _51909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _13023_, clk);
  dff _51910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _13024_, clk);
  dff _51911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _13025_, clk);
  dff _51912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _13027_, clk);
  dff _51913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _13008_, clk);
  dff _51914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _13009_, clk);
  dff _51915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _13011_, clk);
  dff _51916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _13012_, clk);
  dff _51917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _13013_, clk);
  dff _51918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _13015_, clk);
  dff _51919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _13016_, clk);
  dff _51920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _13017_, clk);
  dff _51921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _12999_, clk);
  dff _51922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _13000_, clk);
  dff _51923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _13001_, clk);
  dff _51924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _13003_, clk);
  dff _51925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _13004_, clk);
  dff _51926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _13005_, clk);
  dff _51927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _13006_, clk);
  dff _51928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _13007_, clk);
  dff _51929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _12989_, clk);
  dff _51930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _12991_, clk);
  dff _51931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _12992_, clk);
  dff _51932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _12993_, clk);
  dff _51933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _12994_, clk);
  dff _51934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _12995_, clk);
  dff _51935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _12996_, clk);
  dff _51936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _12997_, clk);
  dff _51937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _12980_, clk);
  dff _51938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _12981_, clk);
  dff _51939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _12982_, clk);
  dff _51940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _12983_, clk);
  dff _51941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _12984_, clk);
  dff _51942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _12985_, clk);
  dff _51943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _12987_, clk);
  dff _51944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _12988_, clk);
  dff _51945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _12970_, clk);
  dff _51946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _12971_, clk);
  dff _51947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _12972_, clk);
  dff _51948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _12973_, clk);
  dff _51949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _12975_, clk);
  dff _51950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _12976_, clk);
  dff _51951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _12977_, clk);
  dff _51952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _12978_, clk);
  dff _51953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _12960_, clk);
  dff _51954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _12961_, clk);
  dff _51955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _12963_, clk);
  dff _51956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _12964_, clk);
  dff _51957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _12965_, clk);
  dff _51958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _12967_, clk);
  dff _51959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _12968_, clk);
  dff _51960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _12969_, clk);
  dff _51961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _12951_, clk);
  dff _51962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _12952_, clk);
  dff _51963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _12953_, clk);
  dff _51964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _12955_, clk);
  dff _51965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _12956_, clk);
  dff _51966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _12957_, clk);
  dff _51967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _12958_, clk);
  dff _51968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _12959_, clk);
  dff _51969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _12941_, clk);
  dff _51970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _12943_, clk);
  dff _51971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _12944_, clk);
  dff _51972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _12945_, clk);
  dff _51973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _12946_, clk);
  dff _51974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _12947_, clk);
  dff _51975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _12948_, clk);
  dff _51976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _12949_, clk);
  dff _51977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _12932_, clk);
  dff _51978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _12933_, clk);
  dff _51979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _12934_, clk);
  dff _51980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _12935_, clk);
  dff _51981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _12936_, clk);
  dff _51982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _12937_, clk);
  dff _51983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _12939_, clk);
  dff _51984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _12940_, clk);
  dff _51985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _12921_, clk);
  dff _51986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _12923_, clk);
  dff _51987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _12924_, clk);
  dff _51988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _12925_, clk);
  dff _51989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _12927_, clk);
  dff _51990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _12928_, clk);
  dff _51991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _12929_, clk);
  dff _51992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _12930_, clk);
  dff _51993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _12912_, clk);
  dff _51994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _12913_, clk);
  dff _51995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _12914_, clk);
  dff _51996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _12915_, clk);
  dff _51997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _12916_, clk);
  dff _51998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _12918_, clk);
  dff _51999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _12919_, clk);
  dff _52000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _12920_, clk);
  dff _52001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _12902_, clk);
  dff _52002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _12903_, clk);
  dff _52003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _12904_, clk);
  dff _52004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _12906_, clk);
  dff _52005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _12907_, clk);
  dff _52006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _12908_, clk);
  dff _52007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _12909_, clk);
  dff _52008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _12911_, clk);
  dff _52009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _12892_, clk);
  dff _52010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _12894_, clk);
  dff _52011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _12895_, clk);
  dff _52012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _12896_, clk);
  dff _52013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _12897_, clk);
  dff _52014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _12899_, clk);
  dff _52015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _12900_, clk);
  dff _52016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _12901_, clk);
  dff _52017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _12883_, clk);
  dff _52018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _12884_, clk);
  dff _52019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _12885_, clk);
  dff _52020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _12887_, clk);
  dff _52021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _12888_, clk);
  dff _52022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _12889_, clk);
  dff _52023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _12890_, clk);
  dff _52024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _12891_, clk);
  dff _52025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _12873_, clk);
  dff _52026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _12875_, clk);
  dff _52027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _12876_, clk);
  dff _52028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _12877_, clk);
  dff _52029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _12878_, clk);
  dff _52030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _12879_, clk);
  dff _52031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _12880_, clk);
  dff _52032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _12881_, clk);
  dff _52033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _12864_, clk);
  dff _52034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _12865_, clk);
  dff _52035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _12866_, clk);
  dff _52036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _12867_, clk);
  dff _52037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _12868_, clk);
  dff _52038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _12870_, clk);
  dff _52039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _12871_, clk);
  dff _52040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _12872_, clk);
  dff _52041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _12854_, clk);
  dff _52042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _12855_, clk);
  dff _52043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _12856_, clk);
  dff _52044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _12858_, clk);
  dff _52045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _12859_, clk);
  dff _52046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _12860_, clk);
  dff _52047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _12861_, clk);
  dff _52048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _12863_, clk);
  dff _52049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _12844_, clk);
  dff _52050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _12846_, clk);
  dff _52051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _12847_, clk);
  dff _52052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _12848_, clk);
  dff _52053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _12849_, clk);
  dff _52054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _12851_, clk);
  dff _52055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _12852_, clk);
  dff _52056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _12853_, clk);
  dff _52057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _12835_, clk);
  dff _52058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _12836_, clk);
  dff _52059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _12837_, clk);
  dff _52060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _12839_, clk);
  dff _52061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _12840_, clk);
  dff _52062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _12841_, clk);
  dff _52063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _12842_, clk);
  dff _52064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _12843_, clk);
  dff _52065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _12825_, clk);
  dff _52066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _12827_, clk);
  dff _52067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _12828_, clk);
  dff _52068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _12829_, clk);
  dff _52069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _12830_, clk);
  dff _52070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _12831_, clk);
  dff _52071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _12832_, clk);
  dff _52072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _12833_, clk);
  dff _52073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _12815_, clk);
  dff _52074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _12816_, clk);
  dff _52075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _12817_, clk);
  dff _52076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _12819_, clk);
  dff _52077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _12820_, clk);
  dff _52078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _12821_, clk);
  dff _52079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _12822_, clk);
  dff _52080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _12824_, clk);
  dff _52081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _12805_, clk);
  dff _52082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _12807_, clk);
  dff _52083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _12808_, clk);
  dff _52084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _12809_, clk);
  dff _52085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _12810_, clk);
  dff _52086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _12811_, clk);
  dff _52087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _12812_, clk);
  dff _52088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _12813_, clk);
  dff _52089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _12796_, clk);
  dff _52090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _12797_, clk);
  dff _52091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _12798_, clk);
  dff _52092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _12799_, clk);
  dff _52093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _12800_, clk);
  dff _52094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _12801_, clk);
  dff _52095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _12803_, clk);
  dff _52096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _12804_, clk);
  dff _52097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _12786_, clk);
  dff _52098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _12787_, clk);
  dff _52099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _12788_, clk);
  dff _52100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _12789_, clk);
  dff _52101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _12791_, clk);
  dff _52102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _12792_, clk);
  dff _52103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _12793_, clk);
  dff _52104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _12794_, clk);
  dff _52105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _12776_, clk);
  dff _52106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _12777_, clk);
  dff _52107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _12779_, clk);
  dff _52108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _12780_, clk);
  dff _52109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _12781_, clk);
  dff _52110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _12783_, clk);
  dff _52111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _12784_, clk);
  dff _52112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _12785_, clk);
  dff _52113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _12767_, clk);
  dff _52114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _12768_, clk);
  dff _52115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _12769_, clk);
  dff _52116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _12771_, clk);
  dff _52117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _12772_, clk);
  dff _52118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _12773_, clk);
  dff _52119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _12774_, clk);
  dff _52120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _12775_, clk);
  dff _52121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _12757_, clk);
  dff _52122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _12759_, clk);
  dff _52123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _12760_, clk);
  dff _52124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _12761_, clk);
  dff _52125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _12762_, clk);
  dff _52126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _12763_, clk);
  dff _52127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _12764_, clk);
  dff _52128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _12765_, clk);
  dff _52129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _12748_, clk);
  dff _52130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _12749_, clk);
  dff _52131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _12750_, clk);
  dff _52132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _12751_, clk);
  dff _52133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _12752_, clk);
  dff _52134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _12753_, clk);
  dff _52135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _12755_, clk);
  dff _52136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _12756_, clk);
  dff _52137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _12738_, clk);
  dff _52138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _12739_, clk);
  dff _52139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _12740_, clk);
  dff _52140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _12741_, clk);
  dff _52141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _12743_, clk);
  dff _52142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _12744_, clk);
  dff _52143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _12745_, clk);
  dff _52144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _12746_, clk);
  dff _52145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _12728_, clk);
  dff _52146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _12729_, clk);
  dff _52147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _12731_, clk);
  dff _52148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _12732_, clk);
  dff _52149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _12733_, clk);
  dff _52150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _12735_, clk);
  dff _52151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _12736_, clk);
  dff _52152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _12737_, clk);
  dff _52153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _12719_, clk);
  dff _52154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _12720_, clk);
  dff _52155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _12721_, clk);
  dff _52156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _12723_, clk);
  dff _52157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _12724_, clk);
  dff _52158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _12725_, clk);
  dff _52159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _12726_, clk);
  dff _52160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _12727_, clk);
  dff _52161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _12708_, clk);
  dff _52162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _12710_, clk);
  dff _52163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _12711_, clk);
  dff _52164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _12712_, clk);
  dff _52165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _12713_, clk);
  dff _52166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _12715_, clk);
  dff _52167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _12716_, clk);
  dff _52168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _12717_, clk);
  dff _52169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _12699_, clk);
  dff _52170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _12700_, clk);
  dff _52171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _12701_, clk);
  dff _52172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _12703_, clk);
  dff _52173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _12704_, clk);
  dff _52174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _12705_, clk);
  dff _52175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _12706_, clk);
  dff _52176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _12707_, clk);
  dff _52177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _12689_, clk);
  dff _52178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _12691_, clk);
  dff _52179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _12692_, clk);
  dff _52180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _12693_, clk);
  dff _52181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _12694_, clk);
  dff _52182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _12695_, clk);
  dff _52183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _12696_, clk);
  dff _52184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _12697_, clk);
  dff _52185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _12680_, clk);
  dff _52186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _12681_, clk);
  dff _52187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _12682_, clk);
  dff _52188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _12683_, clk);
  dff _52189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _12684_, clk);
  dff _52190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _12686_, clk);
  dff _52191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _12687_, clk);
  dff _52192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _12688_, clk);
  dff _52193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _12670_, clk);
  dff _52194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _12671_, clk);
  dff _52195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _12672_, clk);
  dff _52196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _12674_, clk);
  dff _52197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _12675_, clk);
  dff _52198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _12676_, clk);
  dff _52199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _12677_, clk);
  dff _52200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _12679_, clk);
  dff _52201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _12660_, clk);
  dff _52202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _12661_, clk);
  dff _52203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _12663_, clk);
  dff _52204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _12664_, clk);
  dff _52205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _12665_, clk);
  dff _52206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _12667_, clk);
  dff _52207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _12668_, clk);
  dff _52208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _12669_, clk);
  dff _52209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _12651_, clk);
  dff _52210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _12652_, clk);
  dff _52211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _12653_, clk);
  dff _52212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _12655_, clk);
  dff _52213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _12656_, clk);
  dff _52214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _12657_, clk);
  dff _52215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _12658_, clk);
  dff _52216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _12659_, clk);
  dff _52217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _12641_, clk);
  dff _52218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _12643_, clk);
  dff _52219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _12644_, clk);
  dff _52220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _12645_, clk);
  dff _52221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _12646_, clk);
  dff _52222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _12647_, clk);
  dff _52223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _12648_, clk);
  dff _52224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _12649_, clk);
  dff _52225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _12632_, clk);
  dff _52226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _12633_, clk);
  dff _52227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _12634_, clk);
  dff _52228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _12635_, clk);
  dff _52229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _12636_, clk);
  dff _52230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _12637_, clk);
  dff _52231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _12639_, clk);
  dff _52232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _12640_, clk);
  dff _52233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _12622_, clk);
  dff _52234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _12623_, clk);
  dff _52235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _12624_, clk);
  dff _52236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _12625_, clk);
  dff _52237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _12627_, clk);
  dff _52238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _12628_, clk);
  dff _52239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _12629_, clk);
  dff _52240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _12630_, clk);
  dff _52241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _12612_, clk);
  dff _52242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _12613_, clk);
  dff _52243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _12615_, clk);
  dff _52244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _12616_, clk);
  dff _52245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _12617_, clk);
  dff _52246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _12619_, clk);
  dff _52247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _12620_, clk);
  dff _52248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _12621_, clk);
  dff _52249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _12602_, clk);
  dff _52250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _12603_, clk);
  dff _52251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _12604_, clk);
  dff _52252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _12606_, clk);
  dff _52253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _12607_, clk);
  dff _52254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _12608_, clk);
  dff _52255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _12609_, clk);
  dff _52256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _12611_, clk);
  dff _52257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _12592_, clk);
  dff _52258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _12594_, clk);
  dff _52259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _12595_, clk);
  dff _52260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _12596_, clk);
  dff _52261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _12597_, clk);
  dff _52262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _12599_, clk);
  dff _52263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _12600_, clk);
  dff _52264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _12601_, clk);
  dff _52265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _12583_, clk);
  dff _52266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _12584_, clk);
  dff _52267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _12585_, clk);
  dff _52268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _12587_, clk);
  dff _52269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _12588_, clk);
  dff _52270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _12589_, clk);
  dff _52271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _12590_, clk);
  dff _52272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _12591_, clk);
  dff _52273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _12573_, clk);
  dff _52274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _12575_, clk);
  dff _52275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _12576_, clk);
  dff _52276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _12577_, clk);
  dff _52277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _12578_, clk);
  dff _52278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _12579_, clk);
  dff _52279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _12580_, clk);
  dff _52280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _12581_, clk);
  dff _52281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _12564_, clk);
  dff _52282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _12565_, clk);
  dff _52283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _12566_, clk);
  dff _52284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _12567_, clk);
  dff _52285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _12568_, clk);
  dff _52286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _12570_, clk);
  dff _52287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _12571_, clk);
  dff _52288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _12572_, clk);
  dff _52289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _12554_, clk);
  dff _52290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _12555_, clk);
  dff _52291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _12556_, clk);
  dff _52292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _12558_, clk);
  dff _52293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _12559_, clk);
  dff _52294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _12560_, clk);
  dff _52295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _12561_, clk);
  dff _52296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _12563_, clk);
  dff _52297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _12544_, clk);
  dff _52298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _12546_, clk);
  dff _52299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _12547_, clk);
  dff _52300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _12548_, clk);
  dff _52301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _12549_, clk);
  dff _52302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _12551_, clk);
  dff _52303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _12552_, clk);
  dff _52304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _12553_, clk);
  dff _52305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _12535_, clk);
  dff _52306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _12536_, clk);
  dff _52307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _12537_, clk);
  dff _52308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _12539_, clk);
  dff _52309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _12540_, clk);
  dff _52310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _12541_, clk);
  dff _52311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _12542_, clk);
  dff _52312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _12543_, clk);
  dff _52313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _12525_, clk);
  dff _52314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _12527_, clk);
  dff _52315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _12528_, clk);
  dff _52316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _12529_, clk);
  dff _52317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _12530_, clk);
  dff _52318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _12531_, clk);
  dff _52319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _12532_, clk);
  dff _52320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _12533_, clk);
  dff _52321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _12516_, clk);
  dff _52322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _12517_, clk);
  dff _52323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _12518_, clk);
  dff _52324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _12519_, clk);
  dff _52325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _12520_, clk);
  dff _52326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _12522_, clk);
  dff _52327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _12523_, clk);
  dff _52328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _12524_, clk);
  dff _52329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _12505_, clk);
  dff _52330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _12507_, clk);
  dff _52331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _12508_, clk);
  dff _52332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _12509_, clk);
  dff _52333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _12510_, clk);
  dff _52334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _12512_, clk);
  dff _52335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _12513_, clk);
  dff _52336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _12514_, clk);
  dff _52337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _12496_, clk);
  dff _52338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _12497_, clk);
  dff _52339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _12498_, clk);
  dff _52340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _12499_, clk);
  dff _52341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _12500_, clk);
  dff _52342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _12501_, clk);
  dff _52343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _12503_, clk);
  dff _52344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _12504_, clk);
  dff _52345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _12486_, clk);
  dff _52346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _12487_, clk);
  dff _52347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _12488_, clk);
  dff _52348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _12489_, clk);
  dff _52349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _12491_, clk);
  dff _52350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _12492_, clk);
  dff _52351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _12493_, clk);
  dff _52352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _12494_, clk);
  dff _52353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _12476_, clk);
  dff _52354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _12477_, clk);
  dff _52355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _12479_, clk);
  dff _52356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _12480_, clk);
  dff _52357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _12481_, clk);
  dff _52358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _12483_, clk);
  dff _52359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _12484_, clk);
  dff _52360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _12485_, clk);
  dff _52361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _12467_, clk);
  dff _52362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _12468_, clk);
  dff _52363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _12469_, clk);
  dff _52364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _12471_, clk);
  dff _52365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _12472_, clk);
  dff _52366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _12473_, clk);
  dff _52367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _12474_, clk);
  dff _52368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _12475_, clk);
  dff _52369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _12457_, clk);
  dff _52370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _12459_, clk);
  dff _52371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _12460_, clk);
  dff _52372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _12461_, clk);
  dff _52373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _12462_, clk);
  dff _52374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _12463_, clk);
  dff _52375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _12464_, clk);
  dff _52376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _12465_, clk);
  dff _52377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _12448_, clk);
  dff _52378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _12449_, clk);
  dff _52379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _12450_, clk);
  dff _52380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _12451_, clk);
  dff _52381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _12452_, clk);
  dff _52382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _12453_, clk);
  dff _52383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _12455_, clk);
  dff _52384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _12456_, clk);
  dff _52385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _12438_, clk);
  dff _52386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _12439_, clk);
  dff _52387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _12440_, clk);
  dff _52388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _12441_, clk);
  dff _52389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _12443_, clk);
  dff _52390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _12444_, clk);
  dff _52391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _12445_, clk);
  dff _52392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _12446_, clk);
  dff _52393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _12428_, clk);
  dff _52394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _12429_, clk);
  dff _52395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _12431_, clk);
  dff _52396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _12432_, clk);
  dff _52397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _12433_, clk);
  dff _52398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _12435_, clk);
  dff _52399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _12436_, clk);
  dff _52400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _12437_, clk);
  dff _52401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _12419_, clk);
  dff _52402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _12420_, clk);
  dff _52403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _12421_, clk);
  dff _52404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _12423_, clk);
  dff _52405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _12424_, clk);
  dff _52406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _12425_, clk);
  dff _52407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _12426_, clk);
  dff _52408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _12427_, clk);
  dff _52409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _12409_, clk);
  dff _52410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _12411_, clk);
  dff _52411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _12412_, clk);
  dff _52412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _12413_, clk);
  dff _52413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _12414_, clk);
  dff _52414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _12415_, clk);
  dff _52415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _12416_, clk);
  dff _52416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _12417_, clk);
  dff _52417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _12399_, clk);
  dff _52418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _12400_, clk);
  dff _52419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _12401_, clk);
  dff _52420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _12403_, clk);
  dff _52421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _12404_, clk);
  dff _52422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _12405_, clk);
  dff _52423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _12407_, clk);
  dff _52424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _12408_, clk);
  dff _52425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _12389_, clk);
  dff _52426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _12391_, clk);
  dff _52427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _12392_, clk);
  dff _52428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _12393_, clk);
  dff _52429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _12394_, clk);
  dff _52430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _12395_, clk);
  dff _52431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _12396_, clk);
  dff _52432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _12397_, clk);
  dff _52433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _12380_, clk);
  dff _52434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _12381_, clk);
  dff _52435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _12382_, clk);
  dff _52436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _12383_, clk);
  dff _52437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _12384_, clk);
  dff _52438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _12386_, clk);
  dff _52439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _12387_, clk);
  dff _52440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _12388_, clk);
  dff _52441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _12370_, clk);
  dff _52442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _12371_, clk);
  dff _52443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _12372_, clk);
  dff _52444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _12374_, clk);
  dff _52445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _12375_, clk);
  dff _52446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _12376_, clk);
  dff _52447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _12377_, clk);
  dff _52448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _12379_, clk);
  dff _52449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _12360_, clk);
  dff _52450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _12362_, clk);
  dff _52451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _12363_, clk);
  dff _52452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _12364_, clk);
  dff _52453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _12365_, clk);
  dff _52454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _12367_, clk);
  dff _52455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _12368_, clk);
  dff _52456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _12369_, clk);
  dff _52457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _12350_, clk);
  dff _52458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _12352_, clk);
  dff _52459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _12353_, clk);
  dff _52460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _12354_, clk);
  dff _52461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _12356_, clk);
  dff _52462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _12357_, clk);
  dff _52463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _12358_, clk);
  dff _52464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _12359_, clk);
  dff _52465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _12341_, clk);
  dff _52466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _12342_, clk);
  dff _52467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _12344_, clk);
  dff _52468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _12345_, clk);
  dff _52469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _12346_, clk);
  dff _52470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _12347_, clk);
  dff _52471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _12348_, clk);
  dff _52472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _12349_, clk);
  dff _52473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _12331_, clk);
  dff _52474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _12333_, clk);
  dff _52475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _12334_, clk);
  dff _52476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _12335_, clk);
  dff _52477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _12336_, clk);
  dff _52478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _12337_, clk);
  dff _52479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _12338_, clk);
  dff _52480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _12339_, clk);
  dff _52481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _12322_, clk);
  dff _52482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _12323_, clk);
  dff _52483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _12324_, clk);
  dff _52484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _12325_, clk);
  dff _52485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _12326_, clk);
  dff _52486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _12327_, clk);
  dff _52487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _12329_, clk);
  dff _52488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _12330_, clk);
  dff _52489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _12312_, clk);
  dff _52490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _12313_, clk);
  dff _52491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _12314_, clk);
  dff _52492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _12315_, clk);
  dff _52493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _12317_, clk);
  dff _52494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _12318_, clk);
  dff _52495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _12319_, clk);
  dff _52496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _12320_, clk);
  dff _52497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _12302_, clk);
  dff _52498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _12303_, clk);
  dff _52499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _12304_, clk);
  dff _52500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _12306_, clk);
  dff _52501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _12307_, clk);
  dff _52502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _12308_, clk);
  dff _52503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _12310_, clk);
  dff _52504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _12311_, clk);
  dff _52505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _13124_, clk);
  dff _52506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _13125_, clk);
  dff _52507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _13127_, clk);
  dff _52508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _13128_, clk);
  dff _52509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _13129_, clk);
  dff _52510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _13130_, clk);
  dff _52511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _13132_, clk);
  dff _52512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _13133_, clk);
  dff _52513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _14537_, clk);
  dff _52514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _14538_, clk);
  dff _52515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _14539_, clk);
  dff _52516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _14540_, clk);
  dff _52517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _14541_, clk);
  dff _52518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _14542_, clk);
  dff _52519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _14544_, clk);
  dff _52520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _14545_, clk);
  dff _52521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _14527_, clk);
  dff _52522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _14528_, clk);
  dff _52523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _14529_, clk);
  dff _52524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _14530_, clk);
  dff _52525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _14532_, clk);
  dff _52526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _14533_, clk);
  dff _52527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _14534_, clk);
  dff _52528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _14535_, clk);
  dff _52529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _14421_, clk);
  dff _52530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _14422_, clk);
  dff _52531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _14423_, clk);
  dff _52532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _14424_, clk);
  dff _52533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _14425_, clk);
  dff _52534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _14426_, clk);
  dff _52535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _14428_, clk);
  dff _52536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _14429_, clk);
  dff _52537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _14546_, clk);
  dff _52538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _14548_, clk);
  dff _52539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _14549_, clk);
  dff _52540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _14550_, clk);
  dff _52541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _14551_, clk);
  dff _52542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _14552_, clk);
  dff _52543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _14553_, clk);
  dff _52544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _14554_, clk);
  dff _52545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _14430_, clk);
  dff _52546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _14432_, clk);
  dff _52547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _14433_, clk);
  dff _52548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _14434_, clk);
  dff _52549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _14435_, clk);
  dff _52550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _14436_, clk);
  dff _52551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _14437_, clk);
  dff _52552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _14438_, clk);
  dff _52553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _14478_, clk);
  dff _52554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _14480_, clk);
  dff _52555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _14481_, clk);
  dff _52556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _14482_, clk);
  dff _52557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _14483_, clk);
  dff _52558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _14484_, clk);
  dff _52559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _14485_, clk);
  dff _52560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _14486_, clk);
  dff _52561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _14488_, clk);
  dff _52562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _14489_, clk);
  dff _52563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _14490_, clk);
  dff _52564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _14492_, clk);
  dff _52565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _14493_, clk);
  dff _52566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _14494_, clk);
  dff _52567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _14496_, clk);
  dff _52568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _14497_, clk);
  dff _52569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _14150_, clk);
  dff _52570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _14151_, clk);
  dff _52571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _14152_, clk);
  dff _52572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _14153_, clk);
  dff _52573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _14155_, clk);
  dff _52574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _14156_, clk);
  dff _52575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _14157_, clk);
  dff _52576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _14158_, clk);
  dff _52577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _14440_, clk);
  dff _52578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _14441_, clk);
  dff _52579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _14442_, clk);
  dff _52580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _14444_, clk);
  dff _52581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _14445_, clk);
  dff _52582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _14446_, clk);
  dff _52583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _14447_, clk);
  dff _52584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _14448_, clk);
  dff _52585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _14459_, clk);
  dff _52586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _14460_, clk);
  dff _52587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _14461_, clk);
  dff _52588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _14462_, clk);
  dff _52589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _14464_, clk);
  dff _52590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _14465_, clk);
  dff _52591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _14466_, clk);
  dff _52592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _14468_, clk);
  dff _52593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _14469_, clk);
  dff _52594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _14470_, clk);
  dff _52595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _14471_, clk);
  dff _52596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _14472_, clk);
  dff _52597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _14473_, clk);
  dff _52598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _14474_, clk);
  dff _52599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _14476_, clk);
  dff _52600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _14477_, clk);
  dff _52601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _14517_, clk);
  dff _52602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _14518_, clk);
  dff _52603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _14520_, clk);
  dff _52604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _14521_, clk);
  dff _52605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _14522_, clk);
  dff _52606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _14523_, clk);
  dff _52607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _14525_, clk);
  dff _52608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _14526_, clk);
  dff _52609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _14556_, clk);
  dff _52610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _14557_, clk);
  dff _52611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _14558_, clk);
  dff _52612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _14560_, clk);
  dff _52613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _14561_, clk);
  dff _52614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _14562_, clk);
  dff _52615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _14563_, clk);
  dff _52616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _14564_, clk);
  dff _52617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _14605_, clk);
  dff _52618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _14606_, clk);
  dff _52619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _14607_, clk);
  dff _52620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _14608_, clk);
  dff _52621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _14609_, clk);
  dff _52622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _14610_, clk);
  dff _52623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _14611_, clk);
  dff _52624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _14613_, clk);
  dff _52625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _13618_, clk);
  dff _52626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _13619_, clk);
  dff _52627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _13620_, clk);
  dff _52628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _13621_, clk);
  dff _52629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _13622_, clk);
  dff _52630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _13624_, clk);
  dff _52631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _13625_, clk);
  dff _52632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _13626_, clk);
  dff _52633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _13628_, clk);
  dff _52634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _13629_, clk);
  dff _52635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _13630_, clk);
  dff _52636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _13631_, clk);
  dff _52637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _13632_, clk);
  dff _52638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _13633_, clk);
  dff _52639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _13634_, clk);
  dff _52640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _13636_, clk);
  dff _52641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _13646_, clk);
  dff _52642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _13648_, clk);
  dff _52643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _13649_, clk);
  dff _52644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _13650_, clk);
  dff _52645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _13652_, clk);
  dff _52646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _13653_, clk);
  dff _52647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _13654_, clk);
  dff _52648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _13655_, clk);
  dff _52649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _13667_, clk);
  dff _52650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _13668_, clk);
  dff _52651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _13669_, clk);
  dff _52652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _13670_, clk);
  dff _52653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _13671_, clk);
  dff _52654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _13673_, clk);
  dff _52655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _13674_, clk);
  dff _52656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _13675_, clk);
  dff _52657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _13715_, clk);
  dff _52658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _13716_, clk);
  dff _52659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _13717_, clk);
  dff _52660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _13718_, clk);
  dff _52661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _13719_, clk);
  dff _52662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _13721_, clk);
  dff _52663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _13722_, clk);
  dff _52664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _13723_, clk);
  dff _52665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _13734_, clk);
  dff _52666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _13735_, clk);
  dff _52667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _13737_, clk);
  dff _52668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _13738_, clk);
  dff _52669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _13739_, clk);
  dff _52670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _13740_, clk);
  dff _52671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _13741_, clk);
  dff _52672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _13742_, clk);
  dff _52673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _13753_, clk);
  dff _52674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _13754_, clk);
  dff _52675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _13755_, clk);
  dff _52676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _13757_, clk);
  dff _52677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _13758_, clk);
  dff _52678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _13759_, clk);
  dff _52679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _13761_, clk);
  dff _52680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _13762_, clk);
  dff _52681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _13773_, clk);
  dff _52682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _13774_, clk);
  dff _52683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _13775_, clk);
  dff _52684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _13777_, clk);
  dff _52685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _13778_, clk);
  dff _52686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _13779_, clk);
  dff _52687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _13780_, clk);
  dff _52688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _13782_, clk);
  dff _52689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _13792_, clk);
  dff _52690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _13794_, clk);
  dff _52691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _13795_, clk);
  dff _52692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _13796_, clk);
  dff _52693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _13797_, clk);
  dff _52694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _13798_, clk);
  dff _52695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _13799_, clk);
  dff _52696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _13800_, clk);
  dff _52697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _13811_, clk);
  dff _52698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _13813_, clk);
  dff _52699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _13814_, clk);
  dff _52700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _13815_, clk);
  dff _52701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _13816_, clk);
  dff _52702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _13818_, clk);
  dff _52703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _13819_, clk);
  dff _52704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _13820_, clk);
  dff _52705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _13831_, clk);
  dff _52706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _13832_, clk);
  dff _52707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _13833_, clk);
  dff _52708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _13834_, clk);
  dff _52709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _13835_, clk);
  dff _52710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _13837_, clk);
  dff _52711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _13838_, clk);
  dff _52712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _13839_, clk);
  dff _52713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _13850_, clk);
  dff _52714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _13851_, clk);
  dff _52715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _13852_, clk);
  dff _52716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _13854_, clk);
  dff _52717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _13855_, clk);
  dff _52718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _13856_, clk);
  dff _52719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _13857_, clk);
  dff _52720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _13858_, clk);
  dff _52721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _13870_, clk);
  dff _52722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _13871_, clk);
  dff _52723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _13872_, clk);
  dff _52724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _13874_, clk);
  dff _52725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _13875_, clk);
  dff _52726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _13876_, clk);
  dff _52727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _13877_, clk);
  dff _52728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _13878_, clk);
  dff _52729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _13889_, clk);
  dff _52730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _13890_, clk);
  dff _52731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _13891_, clk);
  dff _52732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _13892_, clk);
  dff _52733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _13894_, clk);
  dff _52734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _13895_, clk);
  dff _52735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _13896_, clk);
  dff _52736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _13897_, clk);
  dff _52737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _13908_, clk);
  dff _52738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _13910_, clk);
  dff _52739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _13911_, clk);
  dff _52740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _13912_, clk);
  dff _52741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _13913_, clk);
  dff _52742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _13914_, clk);
  dff _52743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _13915_, clk);
  dff _52744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _13916_, clk);
  dff _52745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _13918_, clk);
  dff _52746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _13919_, clk);
  dff _52747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _13920_, clk);
  dff _52748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _13922_, clk);
  dff _52749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _13923_, clk);
  dff _52750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _13924_, clk);
  dff _52751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _13925_, clk);
  dff _52752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _13926_, clk);
  dff _52753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _13937_, clk);
  dff _52754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _13938_, clk);
  dff _52755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _13939_, clk);
  dff _52756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _13940_, clk);
  dff _52757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _13942_, clk);
  dff _52758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _13943_, clk);
  dff _52759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _13944_, clk);
  dff _52760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _13946_, clk);
  dff _52761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _14005_, clk);
  dff _52762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _14006_, clk);
  dff _52763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _14007_, clk);
  dff _52764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _14008_, clk);
  dff _52765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _14010_, clk);
  dff _52766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _14011_, clk);
  dff _52767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _14012_, clk);
  dff _52768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _14013_, clk);
  dff _52769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _14015_, clk);
  dff _52770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _14016_, clk);
  dff _52771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _14017_, clk);
  dff _52772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _14018_, clk);
  dff _52773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _14019_, clk);
  dff _52774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _14020_, clk);
  dff _52775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _14022_, clk);
  dff _52776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _14023_, clk);
  dff _52777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _14024_, clk);
  dff _52778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _14025_, clk);
  dff _52779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _14027_, clk);
  dff _52780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _14028_, clk);
  dff _52781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _14029_, clk);
  dff _52782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _14030_, clk);
  dff _52783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _14031_, clk);
  dff _52784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _14032_, clk);
  dff _52785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _14034_, clk);
  dff _52786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _14035_, clk);
  dff _52787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _14036_, clk);
  dff _52788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _14037_, clk);
  dff _52789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _14039_, clk);
  dff _52790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _14040_, clk);
  dff _52791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _14041_, clk);
  dff _52792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _14042_, clk);
  dff _52793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _14043_, clk);
  dff _52794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _14044_, clk);
  dff _52795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _14046_, clk);
  dff _52796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _14047_, clk);
  dff _52797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _14048_, clk);
  dff _52798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _14049_, clk);
  dff _52799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _14051_, clk);
  dff _52800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _14052_, clk);
  dff _52801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _14053_, clk);
  dff _52802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _14054_, clk);
  dff _52803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _14055_, clk);
  dff _52804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _14056_, clk);
  dff _52805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _14058_, clk);
  dff _52806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _14059_, clk);
  dff _52807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _14060_, clk);
  dff _52808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _14061_, clk);
  dff _52809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _14063_, clk);
  dff _52810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _14064_, clk);
  dff _52811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _14065_, clk);
  dff _52812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _14066_, clk);
  dff _52813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _14067_, clk);
  dff _52814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _14068_, clk);
  dff _52815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _14070_, clk);
  dff _52816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _14071_, clk);
  dff _52817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _14072_, clk);
  dff _52818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _14074_, clk);
  dff _52819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _14075_, clk);
  dff _52820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _14076_, clk);
  dff _52821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _14078_, clk);
  dff _52822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _14079_, clk);
  dff _52823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _14080_, clk);
  dff _52824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _14081_, clk);
  dff _52825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _14083_, clk);
  dff _52826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _14084_, clk);
  dff _52827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _14085_, clk);
  dff _52828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _14086_, clk);
  dff _52829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _14087_, clk);
  dff _52830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _14088_, clk);
  dff _52831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _14090_, clk);
  dff _52832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _14091_, clk);
  dff _52833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _14092_, clk);
  dff _52834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _14093_, clk);
  dff _52835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _14095_, clk);
  dff _52836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _14096_, clk);
  dff _52837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _14097_, clk);
  dff _52838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _14098_, clk);
  dff _52839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _14099_, clk);
  dff _52840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _14100_, clk);
  dff _52841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _14102_, clk);
  dff _52842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _14103_, clk);
  dff _52843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _14104_, clk);
  dff _52844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _14105_, clk);
  dff _52845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _14107_, clk);
  dff _52846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _14108_, clk);
  dff _52847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _14109_, clk);
  dff _52848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _14110_, clk);
  dff _52849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _14111_, clk);
  dff _52850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _14112_, clk);
  dff _52851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _14114_, clk);
  dff _52852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _14115_, clk);
  dff _52853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _14116_, clk);
  dff _52854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _14117_, clk);
  dff _52855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _14119_, clk);
  dff _52856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _14120_, clk);
  dff _52857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _14121_, clk);
  dff _52858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _14122_, clk);
  dff _52859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _14123_, clk);
  dff _52860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _14124_, clk);
  dff _52861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _14126_, clk);
  dff _52862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _14127_, clk);
  dff _52863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _14128_, clk);
  dff _52864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _14129_, clk);
  dff _52865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _14131_, clk);
  dff _52866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _14132_, clk);
  dff _52867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _14133_, clk);
  dff _52868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _14134_, clk);
  dff _52869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _14135_, clk);
  dff _52870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _14136_, clk);
  dff _52871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _14138_, clk);
  dff _52872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _14139_, clk);
  dff _52873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _14140_, clk);
  dff _52874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _14141_, clk);
  dff _52875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _14143_, clk);
  dff _52876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _14144_, clk);
  dff _52877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _14145_, clk);
  dff _52878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _14146_, clk);
  dff _52879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _14147_, clk);
  dff _52880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _14148_, clk);
  dff _52881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _14159_, clk);
  dff _52882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _14160_, clk);
  dff _52883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _14162_, clk);
  dff _52884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _14163_, clk);
  dff _52885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _14164_, clk);
  dff _52886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _14165_, clk);
  dff _52887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _14167_, clk);
  dff _52888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _14168_, clk);
  dff _52889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _14169_, clk);
  dff _52890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _14170_, clk);
  dff _52891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _14171_, clk);
  dff _52892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _14172_, clk);
  dff _52893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _14174_, clk);
  dff _52894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _14175_, clk);
  dff _52895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _14176_, clk);
  dff _52896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _14177_, clk);
  dff _52897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _14179_, clk);
  dff _52898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _14180_, clk);
  dff _52899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _14181_, clk);
  dff _52900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _14183_, clk);
  dff _52901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _14184_, clk);
  dff _52902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _14185_, clk);
  dff _52903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _14187_, clk);
  dff _52904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _14188_, clk);
  dff _52905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _14189_, clk);
  dff _52906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _14190_, clk);
  dff _52907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _14191_, clk);
  dff _52908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _14192_, clk);
  dff _52909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _14193_, clk);
  dff _52910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _14195_, clk);
  dff _52911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _14196_, clk);
  dff _52912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _14197_, clk);
  dff _52913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _14199_, clk);
  dff _52914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _14200_, clk);
  dff _52915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _14201_, clk);
  dff _52916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _14202_, clk);
  dff _52917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _14203_, clk);
  dff _52918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _14204_, clk);
  dff _52919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _14205_, clk);
  dff _52920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _14207_, clk);
  dff _52921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _14208_, clk);
  dff _52922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _14209_, clk);
  dff _52923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _14211_, clk);
  dff _52924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _14212_, clk);
  dff _52925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _14213_, clk);
  dff _52926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _14214_, clk);
  dff _52927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _14215_, clk);
  dff _52928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _14216_, clk);
  dff _52929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _14217_, clk);
  dff _52930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _14219_, clk);
  dff _52931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _14220_, clk);
  dff _52932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _14221_, clk);
  dff _52933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _14223_, clk);
  dff _52934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _14224_, clk);
  dff _52935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _14225_, clk);
  dff _52936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _14226_, clk);
  dff _52937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _14227_, clk);
  dff _52938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _14228_, clk);
  dff _52939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _14229_, clk);
  dff _52940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _14231_, clk);
  dff _52941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _14232_, clk);
  dff _52942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _14233_, clk);
  dff _52943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _14235_, clk);
  dff _52944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _14236_, clk);
  dff _52945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _14237_, clk);
  dff _52946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _14238_, clk);
  dff _52947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _14239_, clk);
  dff _52948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _14240_, clk);
  dff _52949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _14241_, clk);
  dff _52950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _14243_, clk);
  dff _52951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _14244_, clk);
  dff _52952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _14245_, clk);
  dff _52953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _14247_, clk);
  dff _52954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _14248_, clk);
  dff _52955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _14249_, clk);
  dff _52956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _14250_, clk);
  dff _52957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _14251_, clk);
  dff _52958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _14252_, clk);
  dff _52959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _14253_, clk);
  dff _52960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _14255_, clk);
  dff _52961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _14256_, clk);
  dff _52962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _14257_, clk);
  dff _52963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _14259_, clk);
  dff _52964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _14260_, clk);
  dff _52965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _14261_, clk);
  dff _52966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _14262_, clk);
  dff _52967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _14263_, clk);
  dff _52968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _14264_, clk);
  dff _52969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _14265_, clk);
  dff _52970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _14267_, clk);
  dff _52971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _14268_, clk);
  dff _52972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _14269_, clk);
  dff _52973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _14271_, clk);
  dff _52974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _14272_, clk);
  dff _52975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _14273_, clk);
  dff _52976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _14274_, clk);
  dff _52977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _14275_, clk);
  dff _52978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _14276_, clk);
  dff _52979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _14277_, clk);
  dff _52980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _14279_, clk);
  dff _52981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _14280_, clk);
  dff _52982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _14281_, clk);
  dff _52983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _14283_, clk);
  dff _52984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _14284_, clk);
  dff _52985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _14285_, clk);
  dff _52986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _14287_, clk);
  dff _52987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _14288_, clk);
  dff _52988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _14289_, clk);
  dff _52989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _14290_, clk);
  dff _52990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _14292_, clk);
  dff _52991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _14293_, clk);
  dff _52992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _14294_, clk);
  dff _52993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _14295_, clk);
  dff _52994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _14296_, clk);
  dff _52995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _14297_, clk);
  dff _52996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _14299_, clk);
  dff _52997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _14300_, clk);
  dff _52998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _14301_, clk);
  dff _52999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _14302_, clk);
  dff _53000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _14304_, clk);
  dff _53001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _14305_, clk);
  dff _53002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _14306_, clk);
  dff _53003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _14307_, clk);
  dff _53004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _14308_, clk);
  dff _53005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _14309_, clk);
  dff _53006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _14311_, clk);
  dff _53007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _14312_, clk);
  dff _53008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _14313_, clk);
  dff _53009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _14314_, clk);
  dff _53010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _14316_, clk);
  dff _53011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _14317_, clk);
  dff _53012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _14318_, clk);
  dff _53013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _14319_, clk);
  dff _53014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _14320_, clk);
  dff _53015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _14321_, clk);
  dff _53016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _14322_, clk);
  dff _53017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _14324_, clk);
  dff _53018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _14325_, clk);
  dff _53019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _14326_, clk);
  dff _53020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _14328_, clk);
  dff _53021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _14329_, clk);
  dff _53022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _14330_, clk);
  dff _53023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _14331_, clk);
  dff _53024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _14332_, clk);
  dff _53025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _14333_, clk);
  dff _53026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _14335_, clk);
  dff _53027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _14336_, clk);
  dff _53028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _14337_, clk);
  dff _53029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _14338_, clk);
  dff _53030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _14340_, clk);
  dff _53031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _14341_, clk);
  dff _53032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _14342_, clk);
  dff _53033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _14343_, clk);
  dff _53034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _14344_, clk);
  dff _53035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _14345_, clk);
  dff _53036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _14347_, clk);
  dff _53037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _14348_, clk);
  dff _53038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _14349_, clk);
  dff _53039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _14350_, clk);
  dff _53040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _14352_, clk);
  dff _53041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _14353_, clk);
  dff _53042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _14354_, clk);
  dff _53043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _14355_, clk);
  dff _53044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _14356_, clk);
  dff _53045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _14357_, clk);
  dff _53046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _14359_, clk);
  dff _53047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _14360_, clk);
  dff _53048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _14361_, clk);
  dff _53049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _14362_, clk);
  dff _53050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _14364_, clk);
  dff _53051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _14365_, clk);
  dff _53052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _14366_, clk);
  dff _53053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _14367_, clk);
  dff _53054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _14368_, clk);
  dff _53055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _14369_, clk);
  dff _53056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _14370_, clk);
  dff _53057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _14372_, clk);
  dff _53058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _14373_, clk);
  dff _53059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _14375_, clk);
  dff _53060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _14376_, clk);
  dff _53061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _14377_, clk);
  dff _53062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _14378_, clk);
  dff _53063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _14379_, clk);
  dff _53064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _14380_, clk);
  dff _53065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _14381_, clk);
  dff _53066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _14383_, clk);
  dff _53067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _14384_, clk);
  dff _53068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _14385_, clk);
  dff _53069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _14387_, clk);
  dff _53070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _14388_, clk);
  dff _53071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _14389_, clk);
  dff _53072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _14390_, clk);
  dff _53073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _14392_, clk);
  dff _53074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _14393_, clk);
  dff _53075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _14394_, clk);
  dff _53076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _14396_, clk);
  dff _53077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _14397_, clk);
  dff _53078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _14398_, clk);
  dff _53079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _14399_, clk);
  dff _53080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _14400_, clk);
  dff _53081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _14401_, clk);
  dff _53082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _14402_, clk);
  dff _53083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _14404_, clk);
  dff _53084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _14405_, clk);
  dff _53085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _14406_, clk);
  dff _53086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _14408_, clk);
  dff _53087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _14409_, clk);
  dff _53088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _14410_, clk);
  dff _53089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _14411_, clk);
  dff _53090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _14412_, clk);
  dff _53091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _14413_, clk);
  dff _53092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _14414_, clk);
  dff _53093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _14416_, clk);
  dff _53094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _14417_, clk);
  dff _53095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _14418_, clk);
  dff _53096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _14420_, clk);
  dff _53097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _14449_, clk);
  dff _53098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _14450_, clk);
  dff _53099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _14452_, clk);
  dff _53100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _14453_, clk);
  dff _53101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _14454_, clk);
  dff _53102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _14456_, clk);
  dff _53103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _14457_, clk);
  dff _53104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _14458_, clk);
  dff _53105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _14498_, clk);
  dff _53106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _14499_, clk);
  dff _53107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _14501_, clk);
  dff _53108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _14502_, clk);
  dff _53109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _14503_, clk);
  dff _53110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _14504_, clk);
  dff _53111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _14505_, clk);
  dff _53112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _14506_, clk);
  dff _53113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _14508_, clk);
  dff _53114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _14509_, clk);
  dff _53115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _14510_, clk);
  dff _53116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _14511_, clk);
  dff _53117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _14513_, clk);
  dff _53118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _14514_, clk);
  dff _53119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _14515_, clk);
  dff _53120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _14516_, clk);
  dff _53121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _14565_, clk);
  dff _53122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _14566_, clk);
  dff _53123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _14568_, clk);
  dff _53124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _14569_, clk);
  dff _53125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _14570_, clk);
  dff _53126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _14572_, clk);
  dff _53127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _14573_, clk);
  dff _53128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _14574_, clk);
  dff _53129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0], _14681_, clk);
  dff _53130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1], _14683_, clk);
  dff _53131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2], _14684_, clk);
  dff _53132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3], _14685_, clk);
  dff _53133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4], _14687_, clk);
  dff _53134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5], _14688_, clk);
  dff _53135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6], _14689_, clk);
  dff _53136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7], _02668_, clk);
  dff _53137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _14575_, clk);
  dff _53138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _14576_, clk);
  dff _53139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _14577_, clk);
  dff _53140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _14578_, clk);
  dff _53141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _14580_, clk);
  dff _53142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _14581_, clk);
  dff _53143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _14582_, clk);
  dff _53144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _14583_, clk);
  dff _53145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _14671_, clk);
  dff _53146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _14673_, clk);
  dff _53147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _14674_, clk);
  dff _53148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _14675_, clk);
  dff _53149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _14677_, clk);
  dff _53150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _14678_, clk);
  dff _53151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _14679_, clk);
  dff _53152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _14680_, clk);
  dff _53153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _14662_, clk);
  dff _53154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _14663_, clk);
  dff _53155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _14665_, clk);
  dff _53156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _14666_, clk);
  dff _53157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _14667_, clk);
  dff _53158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _14668_, clk);
  dff _53159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _14669_, clk);
  dff _53160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _14670_, clk);
  dff _53161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _14585_, clk);
  dff _53162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _14586_, clk);
  dff _53163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _14587_, clk);
  dff _53164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _14588_, clk);
  dff _53165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _14589_, clk);
  dff _53166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _14590_, clk);
  dff _53167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _14592_, clk);
  dff _53168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _14593_, clk);
  dff _53169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _14653_, clk);
  dff _53170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _14654_, clk);
  dff _53171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _14655_, clk);
  dff _53172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _14656_, clk);
  dff _53173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _14657_, clk);
  dff _53174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _14658_, clk);
  dff _53175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _14659_, clk);
  dff _53176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _14661_, clk);
  dff _53177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _14594_, clk);
  dff _53178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _14596_, clk);
  dff _53179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _14597_, clk);
  dff _53180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _14598_, clk);
  dff _53181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _14599_, clk);
  dff _53182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _14601_, clk);
  dff _53183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _14602_, clk);
  dff _53184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _14603_, clk);
  dff _53185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _14643_, clk);
  dff _53186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _14644_, clk);
  dff _53187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _14645_, clk);
  dff _53188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _14646_, clk);
  dff _53189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _14647_, clk);
  dff _53190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _14649_, clk);
  dff _53191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _14650_, clk);
  dff _53192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _14651_, clk);
  dff _53193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _14633_, clk);
  dff _53194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _14634_, clk);
  dff _53195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _14635_, clk);
  dff _53196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _14637_, clk);
  dff _53197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _14638_, clk);
  dff _53198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _14639_, clk);
  dff _53199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _14641_, clk);
  dff _53200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _14642_, clk);
  dff _53201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _14614_, clk);
  dff _53202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _14615_, clk);
  dff _53203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _14617_, clk);
  dff _53204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _14618_, clk);
  dff _53205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _14619_, clk);
  dff _53206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _14620_, clk);
  dff _53207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _14621_, clk);
  dff _53208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _14622_, clk);
  dff _53209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _14623_, clk);
  dff _53210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _14625_, clk);
  dff _53211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _14626_, clk);
  dff _53212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _14627_, clk);
  dff _53213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _14629_, clk);
  dff _53214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _14630_, clk);
  dff _53215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _14631_, clk);
  dff _53216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _14632_, clk);
  dff _53217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _14803_, clk);
  dff _53218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _14804_, clk);
  dff _53219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _14805_, clk);
  dff _53220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _14806_, clk);
  dff _53221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _14807_, clk);
  dff _53222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _14808_, clk);
  dff _53223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _14809_, clk);
  dff _53224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02659_, clk);
  dff _53225_ (\oc8051_top_1.oc8051_rom1.data_o [0], 1'b0, clk);
  dff _53226_ (\oc8051_top_1.oc8051_rom1.data_o [1], 1'b0, clk);
  dff _53227_ (\oc8051_top_1.oc8051_rom1.data_o [2], 1'b0, clk);
  dff _53228_ (\oc8051_top_1.oc8051_rom1.data_o [3], 1'b0, clk);
  dff _53229_ (\oc8051_top_1.oc8051_rom1.data_o [4], 1'b0, clk);
  dff _53230_ (\oc8051_top_1.oc8051_rom1.data_o [5], 1'b0, clk);
  dff _53231_ (\oc8051_top_1.oc8051_rom1.data_o [6], 1'b0, clk);
  dff _53232_ (\oc8051_top_1.oc8051_rom1.data_o [7], 1'b0, clk);
  dff _53233_ (\oc8051_top_1.oc8051_rom1.data_o [8], 1'b0, clk);
  dff _53234_ (\oc8051_top_1.oc8051_rom1.data_o [9], 1'b0, clk);
  dff _53235_ (\oc8051_top_1.oc8051_rom1.data_o [10], 1'b0, clk);
  dff _53236_ (\oc8051_top_1.oc8051_rom1.data_o [11], 1'b0, clk);
  dff _53237_ (\oc8051_top_1.oc8051_rom1.data_o [12], 1'b0, clk);
  dff _53238_ (\oc8051_top_1.oc8051_rom1.data_o [13], 1'b0, clk);
  dff _53239_ (\oc8051_top_1.oc8051_rom1.data_o [14], 1'b0, clk);
  dff _53240_ (\oc8051_top_1.oc8051_rom1.data_o [15], 1'b0, clk);
  dff _53241_ (\oc8051_top_1.oc8051_rom1.data_o [16], 1'b0, clk);
  dff _53242_ (\oc8051_top_1.oc8051_rom1.data_o [17], 1'b0, clk);
  dff _53243_ (\oc8051_top_1.oc8051_rom1.data_o [18], 1'b0, clk);
  dff _53244_ (\oc8051_top_1.oc8051_rom1.data_o [19], 1'b0, clk);
  dff _53245_ (\oc8051_top_1.oc8051_rom1.data_o [20], 1'b0, clk);
  dff _53246_ (\oc8051_top_1.oc8051_rom1.data_o [21], 1'b0, clk);
  dff _53247_ (\oc8051_top_1.oc8051_rom1.data_o [22], 1'b0, clk);
  dff _53248_ (\oc8051_top_1.oc8051_rom1.data_o [23], 1'b0, clk);
  dff _53249_ (\oc8051_top_1.oc8051_rom1.data_o [24], 1'b0, clk);
  dff _53250_ (\oc8051_top_1.oc8051_rom1.data_o [25], 1'b0, clk);
  dff _53251_ (\oc8051_top_1.oc8051_rom1.data_o [26], 1'b0, clk);
  dff _53252_ (\oc8051_top_1.oc8051_rom1.data_o [27], 1'b0, clk);
  dff _53253_ (\oc8051_top_1.oc8051_rom1.data_o [28], 1'b0, clk);
  dff _53254_ (\oc8051_top_1.oc8051_rom1.data_o [29], 1'b0, clk);
  dff _53255_ (\oc8051_top_1.oc8051_rom1.data_o [30], 1'b0, clk);
  dff _53256_ (\oc8051_top_1.oc8051_rom1.data_o [31], 1'b0, clk);
  dff _53257_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _53258_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _06501_, clk);
  dff _53259_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _06515_, clk);
  dff _53260_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _06516_, clk);
  dff _53261_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _06517_, clk);
  dff _53262_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _06502_, clk);
  dff _53263_ (\oc8051_top_1.oc8051_sfr1.bit_out , _06503_, clk);
  dff _53264_ (\oc8051_top_1.oc8051_sfr1.wait_data , _06504_, clk);
  dff _53265_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _06518_, clk);
  dff _53266_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _06519_, clk);
  dff _53267_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _06520_, clk);
  dff _53268_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _06521_, clk);
  dff _53269_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _06522_, clk);
  dff _53270_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _06523_, clk);
  dff _53271_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _06524_, clk);
  dff _53272_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _06505_, clk);
  dff _53273_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _06506_, clk);
  dff _53274_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _22204_, clk);
  dff _53275_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _22213_, clk);
  dff _53276_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _22214_, clk);
  dff _53277_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _22222_, clk);
  dff _53278_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _22233_, clk);
  dff _53279_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _22243_, clk);
  dff _53280_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _22254_, clk);
  dff _53281_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _20533_, clk);
  dff _53282_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _10754_, clk);
  dff _53283_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _10762_, clk);
  dff _53284_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _10770_, clk);
  dff _53285_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _10777_, clk);
  dff _53286_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _10786_, clk);
  dff _53287_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _10793_, clk);
  dff _53288_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _10801_, clk);
  dff _53289_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _08893_, clk);
  dff _53290_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _16111_, clk);
  dff _53291_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _16119_, clk);
  dff _53292_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _16127_, clk);
  dff _53293_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _16135_, clk);
  dff _53294_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _16143_, clk);
  dff _53295_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _16150_, clk);
  dff _53296_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _16159_, clk);
  dff _53297_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _15457_, clk);
  dff _53298_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _16166_, clk);
  dff _53299_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _16175_, clk);
  dff _53300_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _16182_, clk);
  dff _53301_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _16190_, clk);
  dff _53302_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _16198_, clk);
  dff _53303_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _16206_, clk);
  dff _53304_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _16214_, clk);
  dff _53305_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _15472_, clk);
  dff _53306_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _25367_, clk);
  dff _53307_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _25366_, clk);
  dff _53308_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _53309_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _25365_, clk);
  dff _53310_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00010_, clk);
  dff _53311_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00012_, clk);
  dff _53312_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00014_, clk);
  dff _53313_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00016_, clk);
  dff _53314_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00017_, clk);
  dff _53315_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00019_, clk);
  dff _53316_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00021_, clk);
  dff _53317_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _25364_, clk);
  dff _53318_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00022_, clk);
  dff _53319_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _25363_, clk);
  dff _53320_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _25362_, clk);
  dff _53321_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00024_, clk);
  dff _53322_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00026_, clk);
  dff _53323_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _25361_, clk);
  dff _53324_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00028_, clk);
  dff _53325_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00030_, clk);
  dff _53326_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _25360_, clk);
  dff _53327_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00032_, clk);
  dff _53328_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _25359_, clk);
  dff _53329_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00034_, clk);
  dff _53330_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _25358_, clk);
  dff _53331_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _25357_, clk);
  dff _53332_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _25356_, clk);
  dff _53333_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _25355_, clk);
  dff _53334_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _25354_, clk);
  dff _53335_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00036_, clk);
  dff _53336_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00038_, clk);
  dff _53337_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00040_, clk);
  dff _53338_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _25353_, clk);
  dff _53339_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00042_, clk);
  dff _53340_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00044_, clk);
  dff _53341_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00046_, clk);
  dff _53342_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00048_, clk);
  dff _53343_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00050_, clk);
  dff _53344_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00052_, clk);
  dff _53345_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00054_, clk);
  dff _53346_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _25352_, clk);
  dff _53347_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00056_, clk);
  dff _53348_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00058_, clk);
  dff _53349_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00060_, clk);
  dff _53350_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00062_, clk);
  dff _53351_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00064_, clk);
  dff _53352_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00066_, clk);
  dff _53353_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00068_, clk);
  dff _53354_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _25351_, clk);
  dff _53355_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _25278_, clk);
  dff _53356_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _25279_, clk);
  dff _53357_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _25280_, clk);
  dff _53358_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _25281_, clk);
  dff _53359_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _25282_, clk);
  dff _53360_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _25283_, clk);
  dff _53361_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _25284_, clk);
  dff _53362_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _25274_, clk);
  dff _53363_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _25285_, clk);
  dff _53364_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _25286_, clk);
  dff _53365_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _25287_, clk);
  dff _53366_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _25288_, clk);
  dff _53367_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _25289_, clk);
  dff _53368_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _25290_, clk);
  dff _53369_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _25291_, clk);
  dff _53370_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _25275_, clk);
  dff _53371_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _25292_, clk);
  dff _53372_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _25293_, clk);
  dff _53373_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _25294_, clk);
  dff _53374_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _25295_, clk);
  dff _53375_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _25296_, clk);
  dff _53376_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _25297_, clk);
  dff _53377_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _25298_, clk);
  dff _53378_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _25276_, clk);
  dff _53379_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _25299_, clk);
  dff _53380_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _25300_, clk);
  dff _53381_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _25301_, clk);
  dff _53382_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _25302_, clk);
  dff _53383_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _25303_, clk);
  dff _53384_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _25304_, clk);
  dff _53385_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _25305_, clk);
  dff _53386_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _25277_, clk);
  dff _53387_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _19908_, clk);
  dff _53388_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _19919_, clk);
  dff _53389_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _19930_, clk);
  dff _53390_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _19941_, clk);
  dff _53391_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _19952_, clk);
  dff _53392_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _19963_, clk);
  dff _53393_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _17600_, clk);
  dff _53394_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _11184_, clk);
  dff _53395_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _11985_, clk);
  dff _53396_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _11994_, clk);
  dff _53397_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _12002_, clk);
  dff _53398_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _12009_, clk);
  dff _53399_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _12018_, clk);
  dff _53400_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _12026_, clk);
  dff _53401_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _12034_, clk);
  dff _53402_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _11198_, clk);
  dff _53403_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _25306_, clk);
  dff _53404_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _25307_, clk);
  dff _53405_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _25316_, clk);
  dff _53406_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _25317_, clk);
  dff _53407_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _25318_, clk);
  dff _53408_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _25319_, clk);
  dff _53409_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _25320_, clk);
  dff _53410_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _25321_, clk);
  dff _53411_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _25322_, clk);
  dff _53412_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _25308_, clk);
  dff _53413_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _25323_, clk);
  dff _53414_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _25324_, clk);
  dff _53415_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _25325_, clk);
  dff _53416_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _25326_, clk);
  dff _53417_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _25327_, clk);
  dff _53418_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _25328_, clk);
  dff _53419_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _25329_, clk);
  dff _53420_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _25309_, clk);
  dff _53421_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _25310_, clk);
  dff _53422_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _25311_, clk);
  dff _53423_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _25330_, clk);
  dff _53424_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _25331_, clk);
  dff _53425_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _25332_, clk);
  dff _53426_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _25333_, clk);
  dff _53427_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _25334_, clk);
  dff _53428_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _25335_, clk);
  dff _53429_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _25336_, clk);
  dff _53430_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _25312_, clk);
  dff _53431_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _25337_, clk);
  dff _53432_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _25338_, clk);
  dff _53433_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _25339_, clk);
  dff _53434_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _25340_, clk);
  dff _53435_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _25341_, clk);
  dff _53436_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _25342_, clk);
  dff _53437_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _25343_, clk);
  dff _53438_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _25313_, clk);
  dff _53439_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _25314_, clk);
  dff _53440_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _25344_, clk);
  dff _53441_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _25345_, clk);
  dff _53442_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _25346_, clk);
  dff _53443_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _25347_, clk);
  dff _53444_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _25348_, clk);
  dff _53445_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _25349_, clk);
  dff _53446_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _25350_, clk);
  dff _53447_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _25315_, clk);
  dff _53448_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01625_, clk);
  dff _53449_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01628_, clk);
  dff _53450_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01631_, clk);
  dff _53451_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01634_, clk);
  dff _53452_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02181_, clk);
  dff _53453_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02183_, clk);
  dff _53454_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02185_, clk);
  dff _53455_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02187_, clk);
  dff _53456_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02189_, clk);
  dff _53457_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02191_, clk);
  dff _53458_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02193_, clk);
  dff _53459_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01637_, clk);
  dff _53460_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02195_, clk);
  dff _53461_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02197_, clk);
  dff _53462_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02199_, clk);
  dff _53463_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02201_, clk);
  dff _53464_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02203_, clk);
  dff _53465_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02205_, clk);
  dff _53466_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02207_, clk);
  dff _53467_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01640_, clk);
  dff _53468_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01643_, clk);
  dff _53469_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02209_, clk);
  dff _53470_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02211_, clk);
  dff _53471_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02213_, clk);
  dff _53472_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02215_, clk);
  dff _53473_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02217_, clk);
  dff _53474_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02219_, clk);
  dff _53475_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02221_, clk);
  dff _53476_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01646_, clk);
  dff _53477_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02223_, clk);
  dff _53478_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02225_, clk);
  dff _53479_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02227_, clk);
  dff _53480_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02229_, clk);
  dff _53481_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02231_, clk);
  dff _53482_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02233_, clk);
  dff _53483_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02235_, clk);
  dff _53484_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01649_, clk);
  dff _53485_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01652_, clk);
  dff _53486_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02237_, clk);
  dff _53487_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02239_, clk);
  dff _53488_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02241_, clk);
  dff _53489_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02243_, clk);
  dff _53490_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02245_, clk);
  dff _53491_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02247_, clk);
  dff _53492_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02249_, clk);
  dff _53493_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01655_, clk);
  dff _53494_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01196_, clk);
  dff _53495_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01198_, clk);
  dff _53496_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01200_, clk);
  dff _53497_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01202_, clk);
  dff _53498_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01204_, clk);
  dff _53499_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01206_, clk);
  dff _53500_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01208_, clk);
  dff _53501_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01210_, clk);
  dff _53502_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01212_, clk);
  dff _53503_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01214_, clk);
  dff _53504_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01216_, clk);
  dff _53505_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00511_, clk);
  dff _53506_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00488_, clk);
  dff _53507_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00491_, clk);
  dff _53508_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00493_, clk);
  dff _53509_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00496_, clk);
  dff _53510_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00498_, clk);
  dff _53511_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00501_, clk);
  dff _53512_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01218_, clk);
  dff _53513_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00503_, clk);
  dff _53514_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01220_, clk);
  dff _53515_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01222_, clk);
  dff _53516_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01224_, clk);
  dff _53517_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00506_, clk);
  dff _53518_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01226_, clk);
  dff _53519_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01228_, clk);
  dff _53520_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01230_, clk);
  dff _53521_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01232_, clk);
  dff _53522_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01234_, clk);
  dff _53523_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01236_, clk);
  dff _53524_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01238_, clk);
  dff _53525_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00509_, clk);
  dff _53526_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00514_, clk);
  dff _53527_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00517_, clk);
  dff _53528_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00519_, clk);
  dff _53529_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00522_, clk);
  dff _53530_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00525_, clk);
  dff _53531_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01240_, clk);
  dff _53532_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01242_, clk);
  dff _53533_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01244_, clk);
  dff _53534_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00527_, clk);
  dff _53535_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01246_, clk);
  dff _53536_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01248_, clk);
  dff _53537_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01250_, clk);
  dff _53538_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01252_, clk);
  dff _53539_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01254_, clk);
  dff _53540_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01256_, clk);
  dff _53541_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01258_, clk);
  dff _53542_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01260_, clk);
  dff _53543_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01262_, clk);
  dff _53544_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01264_, clk);
  dff _53545_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00530_, clk);
  dff _53546_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01266_, clk);
  dff _53547_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01268_, clk);
  dff _53548_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01270_, clk);
  dff _53549_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01272_, clk);
  dff _53550_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01274_, clk);
  dff _53551_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01276_, clk);
  dff _53552_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01278_, clk);
  dff _53553_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00532_, clk);
  dff _53554_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01280_, clk);
  dff _53555_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01282_, clk);
  dff _53556_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01284_, clk);
  dff _53557_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01286_, clk);
  dff _53558_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01288_, clk);
  dff _53559_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01290_, clk);
  dff _53560_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01292_, clk);
  dff _53561_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00535_, clk);
  dff _53562_ (\uc8051golden_1.IRAM[0] [0], _06726_, clk);
  dff _53563_ (\uc8051golden_1.IRAM[0] [1], _06727_, clk);
  dff _53564_ (\uc8051golden_1.IRAM[0] [2], _06728_, clk);
  dff _53565_ (\uc8051golden_1.IRAM[0] [3], _06729_, clk);
  dff _53566_ (\uc8051golden_1.IRAM[0] [4], _06730_, clk);
  dff _53567_ (\uc8051golden_1.IRAM[0] [5], _06731_, clk);
  dff _53568_ (\uc8051golden_1.IRAM[0] [6], _06732_, clk);
  dff _53569_ (\uc8051golden_1.IRAM[0] [7], _06733_, clk);
  dff _53570_ (\uc8051golden_1.B [0], _09277_, clk);
  dff _53571_ (\uc8051golden_1.B [1], _09278_, clk);
  dff _53572_ (\uc8051golden_1.B [2], _09279_, clk);
  dff _53573_ (\uc8051golden_1.B [3], _09280_, clk);
  dff _53574_ (\uc8051golden_1.B [4], _09281_, clk);
  dff _53575_ (\uc8051golden_1.B [5], _09282_, clk);
  dff _53576_ (\uc8051golden_1.B [6], _09283_, clk);
  dff _53577_ (\uc8051golden_1.B [7], _06584_, clk);
  dff _53578_ (\uc8051golden_1.ACC [0], _09284_, clk);
  dff _53579_ (\uc8051golden_1.ACC [1], _09285_, clk);
  dff _53580_ (\uc8051golden_1.ACC [2], _09286_, clk);
  dff _53581_ (\uc8051golden_1.ACC [3], _09287_, clk);
  dff _53582_ (\uc8051golden_1.ACC [4], _09288_, clk);
  dff _53583_ (\uc8051golden_1.ACC [5], _09289_, clk);
  dff _53584_ (\uc8051golden_1.ACC [6], _09290_, clk);
  dff _53585_ (\uc8051golden_1.ACC [7], _06585_, clk);
  dff _53586_ (\uc8051golden_1.PCON [0], _09291_, clk);
  dff _53587_ (\uc8051golden_1.PCON [1], _09292_, clk);
  dff _53588_ (\uc8051golden_1.PCON [2], _09293_, clk);
  dff _53589_ (\uc8051golden_1.PCON [3], _09294_, clk);
  dff _53590_ (\uc8051golden_1.PCON [4], _09295_, clk);
  dff _53591_ (\uc8051golden_1.PCON [5], _09296_, clk);
  dff _53592_ (\uc8051golden_1.PCON [6], _09297_, clk);
  dff _53593_ (\uc8051golden_1.PCON [7], _06586_, clk);
  dff _53594_ (\uc8051golden_1.TMOD [0], _09298_, clk);
  dff _53595_ (\uc8051golden_1.TMOD [1], _09299_, clk);
  dff _53596_ (\uc8051golden_1.TMOD [2], _09300_, clk);
  dff _53597_ (\uc8051golden_1.TMOD [3], _09301_, clk);
  dff _53598_ (\uc8051golden_1.TMOD [4], _09302_, clk);
  dff _53599_ (\uc8051golden_1.TMOD [5], _09303_, clk);
  dff _53600_ (\uc8051golden_1.TMOD [6], _09304_, clk);
  dff _53601_ (\uc8051golden_1.TMOD [7], _06587_, clk);
  dff _53602_ (\uc8051golden_1.DPL [0], _09305_, clk);
  dff _53603_ (\uc8051golden_1.DPL [1], _09306_, clk);
  dff _53604_ (\uc8051golden_1.DPL [2], _09307_, clk);
  dff _53605_ (\uc8051golden_1.DPL [3], _09309_, clk);
  dff _53606_ (\uc8051golden_1.DPL [4], _09310_, clk);
  dff _53607_ (\uc8051golden_1.DPL [5], _09311_, clk);
  dff _53608_ (\uc8051golden_1.DPL [6], _09312_, clk);
  dff _53609_ (\uc8051golden_1.DPL [7], _06588_, clk);
  dff _53610_ (\uc8051golden_1.DPH [0], _09313_, clk);
  dff _53611_ (\uc8051golden_1.DPH [1], _09314_, clk);
  dff _53612_ (\uc8051golden_1.DPH [2], _09315_, clk);
  dff _53613_ (\uc8051golden_1.DPH [3], _09316_, clk);
  dff _53614_ (\uc8051golden_1.DPH [4], _09317_, clk);
  dff _53615_ (\uc8051golden_1.DPH [5], _09318_, clk);
  dff _53616_ (\uc8051golden_1.DPH [6], _09319_, clk);
  dff _53617_ (\uc8051golden_1.DPH [7], _06590_, clk);
  dff _53618_ (\uc8051golden_1.TL1 [0], _09320_, clk);
  dff _53619_ (\uc8051golden_1.TL1 [1], _09321_, clk);
  dff _53620_ (\uc8051golden_1.TL1 [2], _09322_, clk);
  dff _53621_ (\uc8051golden_1.TL1 [3], _09323_, clk);
  dff _53622_ (\uc8051golden_1.TL1 [4], _09324_, clk);
  dff _53623_ (\uc8051golden_1.TL1 [5], _09325_, clk);
  dff _53624_ (\uc8051golden_1.TL1 [6], _09326_, clk);
  dff _53625_ (\uc8051golden_1.TL1 [7], _06591_, clk);
  dff _53626_ (\uc8051golden_1.TL0 [0], _09327_, clk);
  dff _53627_ (\uc8051golden_1.TL0 [1], _09328_, clk);
  dff _53628_ (\uc8051golden_1.TL0 [2], _09329_, clk);
  dff _53629_ (\uc8051golden_1.TL0 [3], _09330_, clk);
  dff _53630_ (\uc8051golden_1.TL0 [4], _09331_, clk);
  dff _53631_ (\uc8051golden_1.TL0 [5], _09332_, clk);
  dff _53632_ (\uc8051golden_1.TL0 [6], _09333_, clk);
  dff _53633_ (\uc8051golden_1.TL0 [7], _06592_, clk);
  dff _53634_ (\uc8051golden_1.TCON [0], _09335_, clk);
  dff _53635_ (\uc8051golden_1.TCON [1], _09336_, clk);
  dff _53636_ (\uc8051golden_1.TCON [2], _09337_, clk);
  dff _53637_ (\uc8051golden_1.TCON [3], _09338_, clk);
  dff _53638_ (\uc8051golden_1.TCON [4], _09339_, clk);
  dff _53639_ (\uc8051golden_1.TCON [5], _09340_, clk);
  dff _53640_ (\uc8051golden_1.TCON [6], _09341_, clk);
  dff _53641_ (\uc8051golden_1.TCON [7], _06593_, clk);
  dff _53642_ (\uc8051golden_1.TH1 [0], _09342_, clk);
  dff _53643_ (\uc8051golden_1.TH1 [1], _09343_, clk);
  dff _53644_ (\uc8051golden_1.TH1 [2], _09344_, clk);
  dff _53645_ (\uc8051golden_1.TH1 [3], _09345_, clk);
  dff _53646_ (\uc8051golden_1.TH1 [4], _09346_, clk);
  dff _53647_ (\uc8051golden_1.TH1 [5], _09347_, clk);
  dff _53648_ (\uc8051golden_1.TH1 [6], _09348_, clk);
  dff _53649_ (\uc8051golden_1.TH1 [7], _06594_, clk);
  dff _53650_ (\uc8051golden_1.TH0 [0], _09349_, clk);
  dff _53651_ (\uc8051golden_1.TH0 [1], _09350_, clk);
  dff _53652_ (\uc8051golden_1.TH0 [2], _09351_, clk);
  dff _53653_ (\uc8051golden_1.TH0 [3], _09352_, clk);
  dff _53654_ (\uc8051golden_1.TH0 [4], _09353_, clk);
  dff _53655_ (\uc8051golden_1.TH0 [5], _09354_, clk);
  dff _53656_ (\uc8051golden_1.TH0 [6], _09355_, clk);
  dff _53657_ (\uc8051golden_1.TH0 [7], _06595_, clk);
  dff _53658_ (\uc8051golden_1.PC [0], _09357_, clk);
  dff _53659_ (\uc8051golden_1.PC [1], _09358_, clk);
  dff _53660_ (\uc8051golden_1.PC [2], _09359_, clk);
  dff _53661_ (\uc8051golden_1.PC [3], _09360_, clk);
  dff _53662_ (\uc8051golden_1.PC [4], _09361_, clk);
  dff _53663_ (\uc8051golden_1.PC [5], _09362_, clk);
  dff _53664_ (\uc8051golden_1.PC [6], _09363_, clk);
  dff _53665_ (\uc8051golden_1.PC [7], _09364_, clk);
  dff _53666_ (\uc8051golden_1.PC [8], _09365_, clk);
  dff _53667_ (\uc8051golden_1.PC [9], _09366_, clk);
  dff _53668_ (\uc8051golden_1.PC [10], _09367_, clk);
  dff _53669_ (\uc8051golden_1.PC [11], _09368_, clk);
  dff _53670_ (\uc8051golden_1.PC [12], _09369_, clk);
  dff _53671_ (\uc8051golden_1.PC [13], _09370_, clk);
  dff _53672_ (\uc8051golden_1.PC [14], _09371_, clk);
  dff _53673_ (\uc8051golden_1.PC [15], _06596_, clk);
  dff _53674_ (\uc8051golden_1.P2 [0], _09372_, clk);
  dff _53675_ (\uc8051golden_1.P2 [1], _09373_, clk);
  dff _53676_ (\uc8051golden_1.P2 [2], _09374_, clk);
  dff _53677_ (\uc8051golden_1.P2 [3], _09375_, clk);
  dff _53678_ (\uc8051golden_1.P2 [4], _09376_, clk);
  dff _53679_ (\uc8051golden_1.P2 [5], _09377_, clk);
  dff _53680_ (\uc8051golden_1.P2 [6], _09378_, clk);
  dff _53681_ (\uc8051golden_1.P2 [7], _06597_, clk);
  dff _53682_ (\uc8051golden_1.P3 [0], _09379_, clk);
  dff _53683_ (\uc8051golden_1.P3 [1], _09380_, clk);
  dff _53684_ (\uc8051golden_1.P3 [2], _09381_, clk);
  dff _53685_ (\uc8051golden_1.P3 [3], _09382_, clk);
  dff _53686_ (\uc8051golden_1.P3 [4], _09383_, clk);
  dff _53687_ (\uc8051golden_1.P3 [5], _09384_, clk);
  dff _53688_ (\uc8051golden_1.P3 [6], _09385_, clk);
  dff _53689_ (\uc8051golden_1.P3 [7], _06598_, clk);
  dff _53690_ (\uc8051golden_1.P0 [0], _09386_, clk);
  dff _53691_ (\uc8051golden_1.P0 [1], _09387_, clk);
  dff _53692_ (\uc8051golden_1.P0 [2], _09388_, clk);
  dff _53693_ (\uc8051golden_1.P0 [3], _09389_, clk);
  dff _53694_ (\uc8051golden_1.P0 [4], _09390_, clk);
  dff _53695_ (\uc8051golden_1.P0 [5], _09391_, clk);
  dff _53696_ (\uc8051golden_1.P0 [6], _09392_, clk);
  dff _53697_ (\uc8051golden_1.P0 [7], _06599_, clk);
  dff _53698_ (\uc8051golden_1.P1 [0], _09393_, clk);
  dff _53699_ (\uc8051golden_1.P1 [1], _09394_, clk);
  dff _53700_ (\uc8051golden_1.P1 [2], _09395_, clk);
  dff _53701_ (\uc8051golden_1.P1 [3], _09396_, clk);
  dff _53702_ (\uc8051golden_1.P1 [4], _09397_, clk);
  dff _53703_ (\uc8051golden_1.P1 [5], _09398_, clk);
  dff _53704_ (\uc8051golden_1.P1 [6], _09399_, clk);
  dff _53705_ (\uc8051golden_1.P1 [7], _06600_, clk);
  dff _53706_ (\uc8051golden_1.IP [0], _09400_, clk);
  dff _53707_ (\uc8051golden_1.IP [1], _09401_, clk);
  dff _53708_ (\uc8051golden_1.IP [2], _09402_, clk);
  dff _53709_ (\uc8051golden_1.IP [3], _09403_, clk);
  dff _53710_ (\uc8051golden_1.IP [4], _09404_, clk);
  dff _53711_ (\uc8051golden_1.IP [5], _09405_, clk);
  dff _53712_ (\uc8051golden_1.IP [6], _09406_, clk);
  dff _53713_ (\uc8051golden_1.IP [7], _06601_, clk);
  dff _53714_ (\uc8051golden_1.IE [0], _09407_, clk);
  dff _53715_ (\uc8051golden_1.IE [1], _09408_, clk);
  dff _53716_ (\uc8051golden_1.IE [2], _09409_, clk);
  dff _53717_ (\uc8051golden_1.IE [3], _09410_, clk);
  dff _53718_ (\uc8051golden_1.IE [4], _09411_, clk);
  dff _53719_ (\uc8051golden_1.IE [5], _09412_, clk);
  dff _53720_ (\uc8051golden_1.IE [6], _09413_, clk);
  dff _53721_ (\uc8051golden_1.IE [7], _06602_, clk);
  dff _53722_ (\uc8051golden_1.SCON [0], _09414_, clk);
  dff _53723_ (\uc8051golden_1.SCON [1], _09415_, clk);
  dff _53724_ (\uc8051golden_1.SCON [2], _09417_, clk);
  dff _53725_ (\uc8051golden_1.SCON [3], _09418_, clk);
  dff _53726_ (\uc8051golden_1.SCON [4], _09419_, clk);
  dff _53727_ (\uc8051golden_1.SCON [5], _09420_, clk);
  dff _53728_ (\uc8051golden_1.SCON [6], _09421_, clk);
  dff _53729_ (\uc8051golden_1.SCON [7], _06603_, clk);
  dff _53730_ (\uc8051golden_1.SP [0], _09422_, clk);
  dff _53731_ (\uc8051golden_1.SP [1], _09423_, clk);
  dff _53732_ (\uc8051golden_1.SP [2], _09424_, clk);
  dff _53733_ (\uc8051golden_1.SP [3], _09425_, clk);
  dff _53734_ (\uc8051golden_1.SP [4], _09426_, clk);
  dff _53735_ (\uc8051golden_1.SP [5], _09427_, clk);
  dff _53736_ (\uc8051golden_1.SP [6], _09428_, clk);
  dff _53737_ (\uc8051golden_1.SP [7], _06604_, clk);
  dff _53738_ (\uc8051golden_1.SBUF [0], _09429_, clk);
  dff _53739_ (\uc8051golden_1.SBUF [1], _09430_, clk);
  dff _53740_ (\uc8051golden_1.SBUF [2], _09431_, clk);
  dff _53741_ (\uc8051golden_1.SBUF [3], _09432_, clk);
  dff _53742_ (\uc8051golden_1.SBUF [4], _09433_, clk);
  dff _53743_ (\uc8051golden_1.SBUF [5], _09434_, clk);
  dff _53744_ (\uc8051golden_1.SBUF [6], _09435_, clk);
  dff _53745_ (\uc8051golden_1.SBUF [7], _06605_, clk);
  dff _53746_ (\uc8051golden_1.PSW [0], _09436_, clk);
  dff _53747_ (\uc8051golden_1.PSW [1], _09437_, clk);
  dff _53748_ (\uc8051golden_1.PSW [2], _09438_, clk);
  dff _53749_ (\uc8051golden_1.PSW [3], _09439_, clk);
  dff _53750_ (\uc8051golden_1.PSW [4], _09440_, clk);
  dff _53751_ (\uc8051golden_1.PSW [5], _09441_, clk);
  dff _53752_ (\uc8051golden_1.PSW [6], _09442_, clk);
  dff _53753_ (\uc8051golden_1.PSW [7], _06606_, clk);
  dff _53754_ (\uc8051golden_1.IRAM[1] [0], _06734_, clk);
  dff _53755_ (\uc8051golden_1.IRAM[1] [1], _06735_, clk);
  dff _53756_ (\uc8051golden_1.IRAM[1] [2], _06736_, clk);
  dff _53757_ (\uc8051golden_1.IRAM[1] [3], _06737_, clk);
  dff _53758_ (\uc8051golden_1.IRAM[1] [4], _06738_, clk);
  dff _53759_ (\uc8051golden_1.IRAM[1] [5], _06739_, clk);
  dff _53760_ (\uc8051golden_1.IRAM[1] [6], _06740_, clk);
  dff _53761_ (\uc8051golden_1.IRAM[1] [7], _06741_, clk);
  dff _53762_ (\uc8051golden_1.IRAM[2] [0], _06742_, clk);
  dff _53763_ (\uc8051golden_1.IRAM[2] [1], _06743_, clk);
  dff _53764_ (\uc8051golden_1.IRAM[2] [2], _06744_, clk);
  dff _53765_ (\uc8051golden_1.IRAM[2] [3], _06746_, clk);
  dff _53766_ (\uc8051golden_1.IRAM[2] [4], _06747_, clk);
  dff _53767_ (\uc8051golden_1.IRAM[2] [5], _06748_, clk);
  dff _53768_ (\uc8051golden_1.IRAM[2] [6], _06749_, clk);
  dff _53769_ (\uc8051golden_1.IRAM[2] [7], _06750_, clk);
  dff _53770_ (\uc8051golden_1.IRAM[3] [0], _06751_, clk);
  dff _53771_ (\uc8051golden_1.IRAM[3] [1], _06752_, clk);
  dff _53772_ (\uc8051golden_1.IRAM[3] [2], _06753_, clk);
  dff _53773_ (\uc8051golden_1.IRAM[3] [3], _06754_, clk);
  dff _53774_ (\uc8051golden_1.IRAM[3] [4], _06755_, clk);
  dff _53775_ (\uc8051golden_1.IRAM[3] [5], _06756_, clk);
  dff _53776_ (\uc8051golden_1.IRAM[3] [6], _06757_, clk);
  dff _53777_ (\uc8051golden_1.IRAM[3] [7], _06758_, clk);
  dff _53778_ (\uc8051golden_1.IRAM[4] [0], _06759_, clk);
  dff _53779_ (\uc8051golden_1.IRAM[4] [1], _06760_, clk);
  dff _53780_ (\uc8051golden_1.IRAM[4] [2], _06761_, clk);
  dff _53781_ (\uc8051golden_1.IRAM[4] [3], _06762_, clk);
  dff _53782_ (\uc8051golden_1.IRAM[4] [4], _06763_, clk);
  dff _53783_ (\uc8051golden_1.IRAM[4] [5], _06764_, clk);
  dff _53784_ (\uc8051golden_1.IRAM[4] [6], _06765_, clk);
  dff _53785_ (\uc8051golden_1.IRAM[4] [7], _06766_, clk);
  dff _53786_ (\uc8051golden_1.IRAM[5] [0], _06767_, clk);
  dff _53787_ (\uc8051golden_1.IRAM[5] [1], _06768_, clk);
  dff _53788_ (\uc8051golden_1.IRAM[5] [2], _06769_, clk);
  dff _53789_ (\uc8051golden_1.IRAM[5] [3], _06770_, clk);
  dff _53790_ (\uc8051golden_1.IRAM[5] [4], _06771_, clk);
  dff _53791_ (\uc8051golden_1.IRAM[5] [5], _06772_, clk);
  dff _53792_ (\uc8051golden_1.IRAM[5] [6], _06773_, clk);
  dff _53793_ (\uc8051golden_1.IRAM[5] [7], _06774_, clk);
  dff _53794_ (\uc8051golden_1.IRAM[6] [0], _06775_, clk);
  dff _53795_ (\uc8051golden_1.IRAM[6] [1], _06776_, clk);
  dff _53796_ (\uc8051golden_1.IRAM[6] [2], _06778_, clk);
  dff _53797_ (\uc8051golden_1.IRAM[6] [3], _06779_, clk);
  dff _53798_ (\uc8051golden_1.IRAM[6] [4], _06780_, clk);
  dff _53799_ (\uc8051golden_1.IRAM[6] [5], _06781_, clk);
  dff _53800_ (\uc8051golden_1.IRAM[6] [6], _06782_, clk);
  dff _53801_ (\uc8051golden_1.IRAM[6] [7], _06783_, clk);
  dff _53802_ (\uc8051golden_1.IRAM[7] [0], _06784_, clk);
  dff _53803_ (\uc8051golden_1.IRAM[7] [1], _06785_, clk);
  dff _53804_ (\uc8051golden_1.IRAM[7] [2], _06786_, clk);
  dff _53805_ (\uc8051golden_1.IRAM[7] [3], _06787_, clk);
  dff _53806_ (\uc8051golden_1.IRAM[7] [4], _06788_, clk);
  dff _53807_ (\uc8051golden_1.IRAM[7] [5], _06789_, clk);
  dff _53808_ (\uc8051golden_1.IRAM[7] [6], _06790_, clk);
  dff _53809_ (\uc8051golden_1.IRAM[7] [7], _06791_, clk);
  dff _53810_ (\uc8051golden_1.IRAM[8] [0], _06792_, clk);
  dff _53811_ (\uc8051golden_1.IRAM[8] [1], _06793_, clk);
  dff _53812_ (\uc8051golden_1.IRAM[8] [2], _06794_, clk);
  dff _53813_ (\uc8051golden_1.IRAM[8] [3], _06795_, clk);
  dff _53814_ (\uc8051golden_1.IRAM[8] [4], _06796_, clk);
  dff _53815_ (\uc8051golden_1.IRAM[8] [5], _06797_, clk);
  dff _53816_ (\uc8051golden_1.IRAM[8] [6], _06798_, clk);
  dff _53817_ (\uc8051golden_1.IRAM[8] [7], _06799_, clk);
  dff _53818_ (\uc8051golden_1.IRAM[9] [0], _06800_, clk);
  dff _53819_ (\uc8051golden_1.IRAM[9] [1], _06801_, clk);
  dff _53820_ (\uc8051golden_1.IRAM[9] [2], _06802_, clk);
  dff _53821_ (\uc8051golden_1.IRAM[9] [3], _06803_, clk);
  dff _53822_ (\uc8051golden_1.IRAM[9] [4], _06804_, clk);
  dff _53823_ (\uc8051golden_1.IRAM[9] [5], _06805_, clk);
  dff _53824_ (\uc8051golden_1.IRAM[9] [6], _06806_, clk);
  dff _53825_ (\uc8051golden_1.IRAM[9] [7], _06807_, clk);
  dff _53826_ (\uc8051golden_1.IRAM[10] [0], _06808_, clk);
  dff _53827_ (\uc8051golden_1.IRAM[10] [1], _06810_, clk);
  dff _53828_ (\uc8051golden_1.IRAM[10] [2], _06811_, clk);
  dff _53829_ (\uc8051golden_1.IRAM[10] [3], _06812_, clk);
  dff _53830_ (\uc8051golden_1.IRAM[10] [4], _06813_, clk);
  dff _53831_ (\uc8051golden_1.IRAM[10] [5], _06814_, clk);
  dff _53832_ (\uc8051golden_1.IRAM[10] [6], _06815_, clk);
  dff _53833_ (\uc8051golden_1.IRAM[10] [7], _06816_, clk);
  dff _53834_ (\uc8051golden_1.IRAM[11] [0], _06817_, clk);
  dff _53835_ (\uc8051golden_1.IRAM[11] [1], _06818_, clk);
  dff _53836_ (\uc8051golden_1.IRAM[11] [2], _06819_, clk);
  dff _53837_ (\uc8051golden_1.IRAM[11] [3], _06820_, clk);
  dff _53838_ (\uc8051golden_1.IRAM[11] [4], _06821_, clk);
  dff _53839_ (\uc8051golden_1.IRAM[11] [5], _06822_, clk);
  dff _53840_ (\uc8051golden_1.IRAM[11] [6], _06823_, clk);
  dff _53841_ (\uc8051golden_1.IRAM[11] [7], _06824_, clk);
  dff _53842_ (\uc8051golden_1.IRAM[12] [0], _06825_, clk);
  dff _53843_ (\uc8051golden_1.IRAM[12] [1], _06826_, clk);
  dff _53844_ (\uc8051golden_1.IRAM[12] [2], _06827_, clk);
  dff _53845_ (\uc8051golden_1.IRAM[12] [3], _06828_, clk);
  dff _53846_ (\uc8051golden_1.IRAM[12] [4], _06829_, clk);
  dff _53847_ (\uc8051golden_1.IRAM[12] [5], _06830_, clk);
  dff _53848_ (\uc8051golden_1.IRAM[12] [6], _06831_, clk);
  dff _53849_ (\uc8051golden_1.IRAM[12] [7], _06832_, clk);
  dff _53850_ (\uc8051golden_1.IRAM[13] [0], _06833_, clk);
  dff _53851_ (\uc8051golden_1.IRAM[13] [1], _06834_, clk);
  dff _53852_ (\uc8051golden_1.IRAM[13] [2], _06835_, clk);
  dff _53853_ (\uc8051golden_1.IRAM[13] [3], _06836_, clk);
  dff _53854_ (\uc8051golden_1.IRAM[13] [4], _06837_, clk);
  dff _53855_ (\uc8051golden_1.IRAM[13] [5], _06838_, clk);
  dff _53856_ (\uc8051golden_1.IRAM[13] [6], _06839_, clk);
  dff _53857_ (\uc8051golden_1.IRAM[13] [7], _06840_, clk);
  dff _53858_ (\uc8051golden_1.IRAM[14] [0], _06841_, clk);
  dff _53859_ (\uc8051golden_1.IRAM[14] [1], _06843_, clk);
  dff _53860_ (\uc8051golden_1.IRAM[14] [2], _06844_, clk);
  dff _53861_ (\uc8051golden_1.IRAM[14] [3], _06845_, clk);
  dff _53862_ (\uc8051golden_1.IRAM[14] [4], _06846_, clk);
  dff _53863_ (\uc8051golden_1.IRAM[14] [5], _06847_, clk);
  dff _53864_ (\uc8051golden_1.IRAM[14] [6], _06848_, clk);
  dff _53865_ (\uc8051golden_1.IRAM[14] [7], _06849_, clk);
  dff _53866_ (\uc8051golden_1.IRAM[15] [0], _06850_, clk);
  dff _53867_ (\uc8051golden_1.IRAM[15] [1], _06851_, clk);
  dff _53868_ (\uc8051golden_1.IRAM[15] [2], _06852_, clk);
  dff _53869_ (\uc8051golden_1.IRAM[15] [3], _06853_, clk);
  dff _53870_ (\uc8051golden_1.IRAM[15] [4], _06854_, clk);
  dff _53871_ (\uc8051golden_1.IRAM[15] [5], _06855_, clk);
  dff _53872_ (\uc8051golden_1.IRAM[15] [6], _06856_, clk);
  dff _53873_ (\uc8051golden_1.IRAM[15] [7], _06857_, clk);
  dff _53874_ (\uc8051golden_1.IRAM[16] [0], _06858_, clk);
  dff _53875_ (\uc8051golden_1.IRAM[16] [1], _06859_, clk);
  dff _53876_ (\uc8051golden_1.IRAM[16] [2], _06860_, clk);
  dff _53877_ (\uc8051golden_1.IRAM[16] [3], _06861_, clk);
  dff _53878_ (\uc8051golden_1.IRAM[16] [4], _06862_, clk);
  dff _53879_ (\uc8051golden_1.IRAM[16] [5], _06863_, clk);
  dff _53880_ (\uc8051golden_1.IRAM[16] [6], _06864_, clk);
  dff _53881_ (\uc8051golden_1.IRAM[16] [7], _06865_, clk);
  dff _53882_ (\uc8051golden_1.IRAM[17] [0], _06866_, clk);
  dff _53883_ (\uc8051golden_1.IRAM[17] [1], _06867_, clk);
  dff _53884_ (\uc8051golden_1.IRAM[17] [2], _06868_, clk);
  dff _53885_ (\uc8051golden_1.IRAM[17] [3], _06869_, clk);
  dff _53886_ (\uc8051golden_1.IRAM[17] [4], _06870_, clk);
  dff _53887_ (\uc8051golden_1.IRAM[17] [5], _06871_, clk);
  dff _53888_ (\uc8051golden_1.IRAM[17] [6], _06872_, clk);
  dff _53889_ (\uc8051golden_1.IRAM[17] [7], _06873_, clk);
  dff _53890_ (\uc8051golden_1.IRAM[18] [0], _06875_, clk);
  dff _53891_ (\uc8051golden_1.IRAM[18] [1], _06876_, clk);
  dff _53892_ (\uc8051golden_1.IRAM[18] [2], _06877_, clk);
  dff _53893_ (\uc8051golden_1.IRAM[18] [3], _06878_, clk);
  dff _53894_ (\uc8051golden_1.IRAM[18] [4], _06879_, clk);
  dff _53895_ (\uc8051golden_1.IRAM[18] [5], _06880_, clk);
  dff _53896_ (\uc8051golden_1.IRAM[18] [6], _06881_, clk);
  dff _53897_ (\uc8051golden_1.IRAM[18] [7], _06882_, clk);
  dff _53898_ (\uc8051golden_1.IRAM[19] [0], _06883_, clk);
  dff _53899_ (\uc8051golden_1.IRAM[19] [1], _06884_, clk);
  dff _53900_ (\uc8051golden_1.IRAM[19] [2], _06885_, clk);
  dff _53901_ (\uc8051golden_1.IRAM[19] [3], _06886_, clk);
  dff _53902_ (\uc8051golden_1.IRAM[19] [4], _06887_, clk);
  dff _53903_ (\uc8051golden_1.IRAM[19] [5], _06888_, clk);
  dff _53904_ (\uc8051golden_1.IRAM[19] [6], _06889_, clk);
  dff _53905_ (\uc8051golden_1.IRAM[19] [7], _06890_, clk);
  dff _53906_ (\uc8051golden_1.IRAM[20] [0], _06891_, clk);
  dff _53907_ (\uc8051golden_1.IRAM[20] [1], _06892_, clk);
  dff _53908_ (\uc8051golden_1.IRAM[20] [2], _06893_, clk);
  dff _53909_ (\uc8051golden_1.IRAM[20] [3], _06894_, clk);
  dff _53910_ (\uc8051golden_1.IRAM[20] [4], _06895_, clk);
  dff _53911_ (\uc8051golden_1.IRAM[20] [5], _06896_, clk);
  dff _53912_ (\uc8051golden_1.IRAM[20] [6], _06897_, clk);
  dff _53913_ (\uc8051golden_1.IRAM[20] [7], _06898_, clk);
  dff _53914_ (\uc8051golden_1.IRAM[21] [0], _06899_, clk);
  dff _53915_ (\uc8051golden_1.IRAM[21] [1], _06900_, clk);
  dff _53916_ (\uc8051golden_1.IRAM[21] [2], _06901_, clk);
  dff _53917_ (\uc8051golden_1.IRAM[21] [3], _06902_, clk);
  dff _53918_ (\uc8051golden_1.IRAM[21] [4], _06903_, clk);
  dff _53919_ (\uc8051golden_1.IRAM[21] [5], _06904_, clk);
  dff _53920_ (\uc8051golden_1.IRAM[21] [6], _06905_, clk);
  dff _53921_ (\uc8051golden_1.IRAM[21] [7], _06906_, clk);
  dff _53922_ (\uc8051golden_1.IRAM[22] [0], _06907_, clk);
  dff _53923_ (\uc8051golden_1.IRAM[22] [1], _06908_, clk);
  dff _53924_ (\uc8051golden_1.IRAM[22] [2], _06910_, clk);
  dff _53925_ (\uc8051golden_1.IRAM[22] [3], _06911_, clk);
  dff _53926_ (\uc8051golden_1.IRAM[22] [4], _06912_, clk);
  dff _53927_ (\uc8051golden_1.IRAM[22] [5], _06913_, clk);
  dff _53928_ (\uc8051golden_1.IRAM[22] [6], _06914_, clk);
  dff _53929_ (\uc8051golden_1.IRAM[22] [7], _06915_, clk);
  dff _53930_ (\uc8051golden_1.IRAM[23] [0], _06916_, clk);
  dff _53931_ (\uc8051golden_1.IRAM[23] [1], _06917_, clk);
  dff _53932_ (\uc8051golden_1.IRAM[23] [2], _06918_, clk);
  dff _53933_ (\uc8051golden_1.IRAM[23] [3], _06919_, clk);
  dff _53934_ (\uc8051golden_1.IRAM[23] [4], _06920_, clk);
  dff _53935_ (\uc8051golden_1.IRAM[23] [5], _06921_, clk);
  dff _53936_ (\uc8051golden_1.IRAM[23] [6], _06922_, clk);
  dff _53937_ (\uc8051golden_1.IRAM[23] [7], _06923_, clk);
  dff _53938_ (\uc8051golden_1.IRAM[24] [0], _06924_, clk);
  dff _53939_ (\uc8051golden_1.IRAM[24] [1], _06925_, clk);
  dff _53940_ (\uc8051golden_1.IRAM[24] [2], _06926_, clk);
  dff _53941_ (\uc8051golden_1.IRAM[24] [3], _06927_, clk);
  dff _53942_ (\uc8051golden_1.IRAM[24] [4], _06928_, clk);
  dff _53943_ (\uc8051golden_1.IRAM[24] [5], _06929_, clk);
  dff _53944_ (\uc8051golden_1.IRAM[24] [6], _06930_, clk);
  dff _53945_ (\uc8051golden_1.IRAM[24] [7], _06931_, clk);
  dff _53946_ (\uc8051golden_1.IRAM[25] [0], _06932_, clk);
  dff _53947_ (\uc8051golden_1.IRAM[25] [1], _06933_, clk);
  dff _53948_ (\uc8051golden_1.IRAM[25] [2], _06934_, clk);
  dff _53949_ (\uc8051golden_1.IRAM[25] [3], _06935_, clk);
  dff _53950_ (\uc8051golden_1.IRAM[25] [4], _06936_, clk);
  dff _53951_ (\uc8051golden_1.IRAM[25] [5], _06937_, clk);
  dff _53952_ (\uc8051golden_1.IRAM[25] [6], _06938_, clk);
  dff _53953_ (\uc8051golden_1.IRAM[25] [7], _06939_, clk);
  dff _53954_ (\uc8051golden_1.IRAM[26] [0], _06940_, clk);
  dff _53955_ (\uc8051golden_1.IRAM[26] [1], _06941_, clk);
  dff _53956_ (\uc8051golden_1.IRAM[26] [2], _06942_, clk);
  dff _53957_ (\uc8051golden_1.IRAM[26] [3], _06944_, clk);
  dff _53958_ (\uc8051golden_1.IRAM[26] [4], _06945_, clk);
  dff _53959_ (\uc8051golden_1.IRAM[26] [5], _06946_, clk);
  dff _53960_ (\uc8051golden_1.IRAM[26] [6], _06947_, clk);
  dff _53961_ (\uc8051golden_1.IRAM[26] [7], _06948_, clk);
  dff _53962_ (\uc8051golden_1.IRAM[27] [0], _06949_, clk);
  dff _53963_ (\uc8051golden_1.IRAM[27] [1], _06950_, clk);
  dff _53964_ (\uc8051golden_1.IRAM[27] [2], _06951_, clk);
  dff _53965_ (\uc8051golden_1.IRAM[27] [3], _06952_, clk);
  dff _53966_ (\uc8051golden_1.IRAM[27] [4], _06953_, clk);
  dff _53967_ (\uc8051golden_1.IRAM[27] [5], _06954_, clk);
  dff _53968_ (\uc8051golden_1.IRAM[27] [6], _06955_, clk);
  dff _53969_ (\uc8051golden_1.IRAM[27] [7], _06956_, clk);
  dff _53970_ (\uc8051golden_1.IRAM[28] [0], _06957_, clk);
  dff _53971_ (\uc8051golden_1.IRAM[28] [1], _06958_, clk);
  dff _53972_ (\uc8051golden_1.IRAM[28] [2], _06959_, clk);
  dff _53973_ (\uc8051golden_1.IRAM[28] [3], _06960_, clk);
  dff _53974_ (\uc8051golden_1.IRAM[28] [4], _06961_, clk);
  dff _53975_ (\uc8051golden_1.IRAM[28] [5], _06962_, clk);
  dff _53976_ (\uc8051golden_1.IRAM[28] [6], _06963_, clk);
  dff _53977_ (\uc8051golden_1.IRAM[28] [7], _06964_, clk);
  dff _53978_ (\uc8051golden_1.IRAM[29] [0], _06965_, clk);
  dff _53979_ (\uc8051golden_1.IRAM[29] [1], _06966_, clk);
  dff _53980_ (\uc8051golden_1.IRAM[29] [2], _06967_, clk);
  dff _53981_ (\uc8051golden_1.IRAM[29] [3], _06968_, clk);
  dff _53982_ (\uc8051golden_1.IRAM[29] [4], _06969_, clk);
  dff _53983_ (\uc8051golden_1.IRAM[29] [5], _06970_, clk);
  dff _53984_ (\uc8051golden_1.IRAM[29] [6], _06971_, clk);
  dff _53985_ (\uc8051golden_1.IRAM[29] [7], _06972_, clk);
  dff _53986_ (\uc8051golden_1.IRAM[30] [0], _06973_, clk);
  dff _53987_ (\uc8051golden_1.IRAM[30] [1], _06974_, clk);
  dff _53988_ (\uc8051golden_1.IRAM[30] [2], _06975_, clk);
  dff _53989_ (\uc8051golden_1.IRAM[30] [3], _06976_, clk);
  dff _53990_ (\uc8051golden_1.IRAM[30] [4], _06978_, clk);
  dff _53991_ (\uc8051golden_1.IRAM[30] [5], _06979_, clk);
  dff _53992_ (\uc8051golden_1.IRAM[30] [6], _06980_, clk);
  dff _53993_ (\uc8051golden_1.IRAM[30] [7], _06981_, clk);
  dff _53994_ (\uc8051golden_1.IRAM[31] [0], _06982_, clk);
  dff _53995_ (\uc8051golden_1.IRAM[31] [1], _06983_, clk);
  dff _53996_ (\uc8051golden_1.IRAM[31] [2], _06984_, clk);
  dff _53997_ (\uc8051golden_1.IRAM[31] [3], _06985_, clk);
  dff _53998_ (\uc8051golden_1.IRAM[31] [4], _06986_, clk);
  dff _53999_ (\uc8051golden_1.IRAM[31] [5], _06987_, clk);
  dff _54000_ (\uc8051golden_1.IRAM[31] [6], _06988_, clk);
  dff _54001_ (\uc8051golden_1.IRAM[31] [7], _06989_, clk);
  dff _54002_ (\uc8051golden_1.IRAM[32] [0], _06990_, clk);
  dff _54003_ (\uc8051golden_1.IRAM[32] [1], _06991_, clk);
  dff _54004_ (\uc8051golden_1.IRAM[32] [2], _06992_, clk);
  dff _54005_ (\uc8051golden_1.IRAM[32] [3], _06993_, clk);
  dff _54006_ (\uc8051golden_1.IRAM[32] [4], _06994_, clk);
  dff _54007_ (\uc8051golden_1.IRAM[32] [5], _06995_, clk);
  dff _54008_ (\uc8051golden_1.IRAM[32] [6], _06996_, clk);
  dff _54009_ (\uc8051golden_1.IRAM[32] [7], _06997_, clk);
  dff _54010_ (\uc8051golden_1.IRAM[33] [0], _06998_, clk);
  dff _54011_ (\uc8051golden_1.IRAM[33] [1], _06999_, clk);
  dff _54012_ (\uc8051golden_1.IRAM[33] [2], _07000_, clk);
  dff _54013_ (\uc8051golden_1.IRAM[33] [3], _07001_, clk);
  dff _54014_ (\uc8051golden_1.IRAM[33] [4], _07002_, clk);
  dff _54015_ (\uc8051golden_1.IRAM[33] [5], _07003_, clk);
  dff _54016_ (\uc8051golden_1.IRAM[33] [6], _07004_, clk);
  dff _54017_ (\uc8051golden_1.IRAM[33] [7], _07005_, clk);
  dff _54018_ (\uc8051golden_1.IRAM[34] [0], _07006_, clk);
  dff _54019_ (\uc8051golden_1.IRAM[34] [1], _07007_, clk);
  dff _54020_ (\uc8051golden_1.IRAM[34] [2], _07008_, clk);
  dff _54021_ (\uc8051golden_1.IRAM[34] [3], _07009_, clk);
  dff _54022_ (\uc8051golden_1.IRAM[34] [4], _07011_, clk);
  dff _54023_ (\uc8051golden_1.IRAM[34] [5], _07012_, clk);
  dff _54024_ (\uc8051golden_1.IRAM[34] [6], _07013_, clk);
  dff _54025_ (\uc8051golden_1.IRAM[34] [7], _07014_, clk);
  dff _54026_ (\uc8051golden_1.IRAM[35] [0], _07015_, clk);
  dff _54027_ (\uc8051golden_1.IRAM[35] [1], _07016_, clk);
  dff _54028_ (\uc8051golden_1.IRAM[35] [2], _07017_, clk);
  dff _54029_ (\uc8051golden_1.IRAM[35] [3], _07018_, clk);
  dff _54030_ (\uc8051golden_1.IRAM[35] [4], _07019_, clk);
  dff _54031_ (\uc8051golden_1.IRAM[35] [5], _07020_, clk);
  dff _54032_ (\uc8051golden_1.IRAM[35] [6], _07021_, clk);
  dff _54033_ (\uc8051golden_1.IRAM[35] [7], _07022_, clk);
  dff _54034_ (\uc8051golden_1.IRAM[36] [0], _07023_, clk);
  dff _54035_ (\uc8051golden_1.IRAM[36] [1], _07024_, clk);
  dff _54036_ (\uc8051golden_1.IRAM[36] [2], _07025_, clk);
  dff _54037_ (\uc8051golden_1.IRAM[36] [3], _07026_, clk);
  dff _54038_ (\uc8051golden_1.IRAM[36] [4], _07027_, clk);
  dff _54039_ (\uc8051golden_1.IRAM[36] [5], _07028_, clk);
  dff _54040_ (\uc8051golden_1.IRAM[36] [6], _07029_, clk);
  dff _54041_ (\uc8051golden_1.IRAM[36] [7], _07030_, clk);
  dff _54042_ (\uc8051golden_1.IRAM[37] [0], _07031_, clk);
  dff _54043_ (\uc8051golden_1.IRAM[37] [1], _07032_, clk);
  dff _54044_ (\uc8051golden_1.IRAM[37] [2], _07033_, clk);
  dff _54045_ (\uc8051golden_1.IRAM[37] [3], _07034_, clk);
  dff _54046_ (\uc8051golden_1.IRAM[37] [4], _07035_, clk);
  dff _54047_ (\uc8051golden_1.IRAM[37] [5], _07036_, clk);
  dff _54048_ (\uc8051golden_1.IRAM[37] [6], _07037_, clk);
  dff _54049_ (\uc8051golden_1.IRAM[37] [7], _07038_, clk);
  dff _54050_ (\uc8051golden_1.IRAM[38] [0], _07039_, clk);
  dff _54051_ (\uc8051golden_1.IRAM[38] [1], _07040_, clk);
  dff _54052_ (\uc8051golden_1.IRAM[38] [2], _07041_, clk);
  dff _54053_ (\uc8051golden_1.IRAM[38] [3], _07042_, clk);
  dff _54054_ (\uc8051golden_1.IRAM[38] [4], _07043_, clk);
  dff _54055_ (\uc8051golden_1.IRAM[38] [5], _07044_, clk);
  dff _54056_ (\uc8051golden_1.IRAM[38] [6], _07046_, clk);
  dff _54057_ (\uc8051golden_1.IRAM[38] [7], _07047_, clk);
  dff _54058_ (\uc8051golden_1.IRAM[39] [0], _07048_, clk);
  dff _54059_ (\uc8051golden_1.IRAM[39] [1], _07049_, clk);
  dff _54060_ (\uc8051golden_1.IRAM[39] [2], _07050_, clk);
  dff _54061_ (\uc8051golden_1.IRAM[39] [3], _07051_, clk);
  dff _54062_ (\uc8051golden_1.IRAM[39] [4], _07052_, clk);
  dff _54063_ (\uc8051golden_1.IRAM[39] [5], _07053_, clk);
  dff _54064_ (\uc8051golden_1.IRAM[39] [6], _07054_, clk);
  dff _54065_ (\uc8051golden_1.IRAM[39] [7], _07055_, clk);
  dff _54066_ (\uc8051golden_1.IRAM[40] [0], _07056_, clk);
  dff _54067_ (\uc8051golden_1.IRAM[40] [1], _07057_, clk);
  dff _54068_ (\uc8051golden_1.IRAM[40] [2], _07058_, clk);
  dff _54069_ (\uc8051golden_1.IRAM[40] [3], _07059_, clk);
  dff _54070_ (\uc8051golden_1.IRAM[40] [4], _07060_, clk);
  dff _54071_ (\uc8051golden_1.IRAM[40] [5], _07061_, clk);
  dff _54072_ (\uc8051golden_1.IRAM[40] [6], _07062_, clk);
  dff _54073_ (\uc8051golden_1.IRAM[40] [7], _07063_, clk);
  dff _54074_ (\uc8051golden_1.IRAM[41] [0], _07064_, clk);
  dff _54075_ (\uc8051golden_1.IRAM[41] [1], _07065_, clk);
  dff _54076_ (\uc8051golden_1.IRAM[41] [2], _07066_, clk);
  dff _54077_ (\uc8051golden_1.IRAM[41] [3], _07067_, clk);
  dff _54078_ (\uc8051golden_1.IRAM[41] [4], _07068_, clk);
  dff _54079_ (\uc8051golden_1.IRAM[41] [5], _07069_, clk);
  dff _54080_ (\uc8051golden_1.IRAM[41] [6], _07070_, clk);
  dff _54081_ (\uc8051golden_1.IRAM[41] [7], _07071_, clk);
  dff _54082_ (\uc8051golden_1.IRAM[42] [0], _07072_, clk);
  dff _54083_ (\uc8051golden_1.IRAM[42] [1], _07073_, clk);
  dff _54084_ (\uc8051golden_1.IRAM[42] [2], _07074_, clk);
  dff _54085_ (\uc8051golden_1.IRAM[42] [3], _07075_, clk);
  dff _54086_ (\uc8051golden_1.IRAM[42] [4], _07076_, clk);
  dff _54087_ (\uc8051golden_1.IRAM[42] [5], _07077_, clk);
  dff _54088_ (\uc8051golden_1.IRAM[42] [6], _07078_, clk);
  dff _54089_ (\uc8051golden_1.IRAM[42] [7], _07080_, clk);
  dff _54090_ (\uc8051golden_1.IRAM[43] [0], _07081_, clk);
  dff _54091_ (\uc8051golden_1.IRAM[43] [1], _07082_, clk);
  dff _54092_ (\uc8051golden_1.IRAM[43] [2], _07083_, clk);
  dff _54093_ (\uc8051golden_1.IRAM[43] [3], _07084_, clk);
  dff _54094_ (\uc8051golden_1.IRAM[43] [4], _07085_, clk);
  dff _54095_ (\uc8051golden_1.IRAM[43] [5], _07086_, clk);
  dff _54096_ (\uc8051golden_1.IRAM[43] [6], _07087_, clk);
  dff _54097_ (\uc8051golden_1.IRAM[43] [7], _07088_, clk);
  dff _54098_ (\uc8051golden_1.IRAM[44] [0], _07089_, clk);
  dff _54099_ (\uc8051golden_1.IRAM[44] [1], _07090_, clk);
  dff _54100_ (\uc8051golden_1.IRAM[44] [2], _07091_, clk);
  dff _54101_ (\uc8051golden_1.IRAM[44] [3], _07092_, clk);
  dff _54102_ (\uc8051golden_1.IRAM[44] [4], _07093_, clk);
  dff _54103_ (\uc8051golden_1.IRAM[44] [5], _07094_, clk);
  dff _54104_ (\uc8051golden_1.IRAM[44] [6], _07095_, clk);
  dff _54105_ (\uc8051golden_1.IRAM[44] [7], _07096_, clk);
  dff _54106_ (\uc8051golden_1.IRAM[45] [0], _07097_, clk);
  dff _54107_ (\uc8051golden_1.IRAM[45] [1], _07098_, clk);
  dff _54108_ (\uc8051golden_1.IRAM[45] [2], _07099_, clk);
  dff _54109_ (\uc8051golden_1.IRAM[45] [3], _07100_, clk);
  dff _54110_ (\uc8051golden_1.IRAM[45] [4], _07101_, clk);
  dff _54111_ (\uc8051golden_1.IRAM[45] [5], _07102_, clk);
  dff _54112_ (\uc8051golden_1.IRAM[45] [6], _07103_, clk);
  dff _54113_ (\uc8051golden_1.IRAM[45] [7], _07104_, clk);
  dff _54114_ (\uc8051golden_1.IRAM[46] [0], _07105_, clk);
  dff _54115_ (\uc8051golden_1.IRAM[46] [1], _07106_, clk);
  dff _54116_ (\uc8051golden_1.IRAM[46] [2], _07107_, clk);
  dff _54117_ (\uc8051golden_1.IRAM[46] [3], _07108_, clk);
  dff _54118_ (\uc8051golden_1.IRAM[46] [4], _07109_, clk);
  dff _54119_ (\uc8051golden_1.IRAM[46] [5], _07110_, clk);
  dff _54120_ (\uc8051golden_1.IRAM[46] [6], _07111_, clk);
  dff _54121_ (\uc8051golden_1.IRAM[46] [7], _07112_, clk);
  dff _54122_ (\uc8051golden_1.IRAM[47] [0], _07114_, clk);
  dff _54123_ (\uc8051golden_1.IRAM[47] [1], _07115_, clk);
  dff _54124_ (\uc8051golden_1.IRAM[47] [2], _07116_, clk);
  dff _54125_ (\uc8051golden_1.IRAM[47] [3], _07117_, clk);
  dff _54126_ (\uc8051golden_1.IRAM[47] [4], _07118_, clk);
  dff _54127_ (\uc8051golden_1.IRAM[47] [5], _07119_, clk);
  dff _54128_ (\uc8051golden_1.IRAM[47] [6], _07120_, clk);
  dff _54129_ (\uc8051golden_1.IRAM[47] [7], _07121_, clk);
  dff _54130_ (\uc8051golden_1.IRAM[48] [0], _07122_, clk);
  dff _54131_ (\uc8051golden_1.IRAM[48] [1], _07123_, clk);
  dff _54132_ (\uc8051golden_1.IRAM[48] [2], _07124_, clk);
  dff _54133_ (\uc8051golden_1.IRAM[48] [3], _07125_, clk);
  dff _54134_ (\uc8051golden_1.IRAM[48] [4], _07126_, clk);
  dff _54135_ (\uc8051golden_1.IRAM[48] [5], _07127_, clk);
  dff _54136_ (\uc8051golden_1.IRAM[48] [6], _07128_, clk);
  dff _54137_ (\uc8051golden_1.IRAM[48] [7], _07129_, clk);
  dff _54138_ (\uc8051golden_1.IRAM[49] [0], _07130_, clk);
  dff _54139_ (\uc8051golden_1.IRAM[49] [1], _07131_, clk);
  dff _54140_ (\uc8051golden_1.IRAM[49] [2], _07132_, clk);
  dff _54141_ (\uc8051golden_1.IRAM[49] [3], _07133_, clk);
  dff _54142_ (\uc8051golden_1.IRAM[49] [4], _07134_, clk);
  dff _54143_ (\uc8051golden_1.IRAM[49] [5], _07135_, clk);
  dff _54144_ (\uc8051golden_1.IRAM[49] [6], _07136_, clk);
  dff _54145_ (\uc8051golden_1.IRAM[49] [7], _07137_, clk);
  dff _54146_ (\uc8051golden_1.IRAM[50] [0], _07138_, clk);
  dff _54147_ (\uc8051golden_1.IRAM[50] [1], _07139_, clk);
  dff _54148_ (\uc8051golden_1.IRAM[50] [2], _07140_, clk);
  dff _54149_ (\uc8051golden_1.IRAM[50] [3], _07141_, clk);
  dff _54150_ (\uc8051golden_1.IRAM[50] [4], _07142_, clk);
  dff _54151_ (\uc8051golden_1.IRAM[50] [5], _07143_, clk);
  dff _54152_ (\uc8051golden_1.IRAM[50] [6], _07144_, clk);
  dff _54153_ (\uc8051golden_1.IRAM[50] [7], _07145_, clk);
  dff _54154_ (\uc8051golden_1.IRAM[51] [0], _07146_, clk);
  dff _54155_ (\uc8051golden_1.IRAM[51] [1], _07148_, clk);
  dff _54156_ (\uc8051golden_1.IRAM[51] [2], _07149_, clk);
  dff _54157_ (\uc8051golden_1.IRAM[51] [3], _07150_, clk);
  dff _54158_ (\uc8051golden_1.IRAM[51] [4], _07151_, clk);
  dff _54159_ (\uc8051golden_1.IRAM[51] [5], _07152_, clk);
  dff _54160_ (\uc8051golden_1.IRAM[51] [6], _07153_, clk);
  dff _54161_ (\uc8051golden_1.IRAM[51] [7], _07154_, clk);
  dff _54162_ (\uc8051golden_1.IRAM[52] [0], _07155_, clk);
  dff _54163_ (\uc8051golden_1.IRAM[52] [1], _07156_, clk);
  dff _54164_ (\uc8051golden_1.IRAM[52] [2], _07157_, clk);
  dff _54165_ (\uc8051golden_1.IRAM[52] [3], _07158_, clk);
  dff _54166_ (\uc8051golden_1.IRAM[52] [4], _07159_, clk);
  dff _54167_ (\uc8051golden_1.IRAM[52] [5], _07160_, clk);
  dff _54168_ (\uc8051golden_1.IRAM[52] [6], _07161_, clk);
  dff _54169_ (\uc8051golden_1.IRAM[52] [7], _07162_, clk);
  dff _54170_ (\uc8051golden_1.IRAM[53] [0], _07163_, clk);
  dff _54171_ (\uc8051golden_1.IRAM[53] [1], _07164_, clk);
  dff _54172_ (\uc8051golden_1.IRAM[53] [2], _07165_, clk);
  dff _54173_ (\uc8051golden_1.IRAM[53] [3], _07166_, clk);
  dff _54174_ (\uc8051golden_1.IRAM[53] [4], _07167_, clk);
  dff _54175_ (\uc8051golden_1.IRAM[53] [5], _07168_, clk);
  dff _54176_ (\uc8051golden_1.IRAM[53] [6], _07169_, clk);
  dff _54177_ (\uc8051golden_1.IRAM[53] [7], _07170_, clk);
  dff _54178_ (\uc8051golden_1.IRAM[54] [0], _07171_, clk);
  dff _54179_ (\uc8051golden_1.IRAM[54] [1], _07172_, clk);
  dff _54180_ (\uc8051golden_1.IRAM[54] [2], _07173_, clk);
  dff _54181_ (\uc8051golden_1.IRAM[54] [3], _07174_, clk);
  dff _54182_ (\uc8051golden_1.IRAM[54] [4], _07175_, clk);
  dff _54183_ (\uc8051golden_1.IRAM[54] [5], _07176_, clk);
  dff _54184_ (\uc8051golden_1.IRAM[54] [6], _07177_, clk);
  dff _54185_ (\uc8051golden_1.IRAM[54] [7], _07178_, clk);
  dff _54186_ (\uc8051golden_1.IRAM[55] [0], _07179_, clk);
  dff _54187_ (\uc8051golden_1.IRAM[55] [1], _07180_, clk);
  dff _54188_ (\uc8051golden_1.IRAM[55] [2], _07182_, clk);
  dff _54189_ (\uc8051golden_1.IRAM[55] [3], _07183_, clk);
  dff _54190_ (\uc8051golden_1.IRAM[55] [4], _07184_, clk);
  dff _54191_ (\uc8051golden_1.IRAM[55] [5], _07185_, clk);
  dff _54192_ (\uc8051golden_1.IRAM[55] [6], _07186_, clk);
  dff _54193_ (\uc8051golden_1.IRAM[55] [7], _07187_, clk);
  dff _54194_ (\uc8051golden_1.IRAM[56] [0], _07188_, clk);
  dff _54195_ (\uc8051golden_1.IRAM[56] [1], _07189_, clk);
  dff _54196_ (\uc8051golden_1.IRAM[56] [2], _07190_, clk);
  dff _54197_ (\uc8051golden_1.IRAM[56] [3], _07191_, clk);
  dff _54198_ (\uc8051golden_1.IRAM[56] [4], _07192_, clk);
  dff _54199_ (\uc8051golden_1.IRAM[56] [5], _07193_, clk);
  dff _54200_ (\uc8051golden_1.IRAM[56] [6], _07194_, clk);
  dff _54201_ (\uc8051golden_1.IRAM[56] [7], _07195_, clk);
  dff _54202_ (\uc8051golden_1.IRAM[57] [0], _07196_, clk);
  dff _54203_ (\uc8051golden_1.IRAM[57] [1], _07197_, clk);
  dff _54204_ (\uc8051golden_1.IRAM[57] [2], _07198_, clk);
  dff _54205_ (\uc8051golden_1.IRAM[57] [3], _07199_, clk);
  dff _54206_ (\uc8051golden_1.IRAM[57] [4], _07200_, clk);
  dff _54207_ (\uc8051golden_1.IRAM[57] [5], _07201_, clk);
  dff _54208_ (\uc8051golden_1.IRAM[57] [6], _07202_, clk);
  dff _54209_ (\uc8051golden_1.IRAM[57] [7], _07203_, clk);
  dff _54210_ (\uc8051golden_1.IRAM[58] [0], _07204_, clk);
  dff _54211_ (\uc8051golden_1.IRAM[58] [1], _07205_, clk);
  dff _54212_ (\uc8051golden_1.IRAM[58] [2], _07206_, clk);
  dff _54213_ (\uc8051golden_1.IRAM[58] [3], _07207_, clk);
  dff _54214_ (\uc8051golden_1.IRAM[58] [4], _07208_, clk);
  dff _54215_ (\uc8051golden_1.IRAM[58] [5], _07209_, clk);
  dff _54216_ (\uc8051golden_1.IRAM[58] [6], _07210_, clk);
  dff _54217_ (\uc8051golden_1.IRAM[58] [7], _07211_, clk);
  dff _54218_ (\uc8051golden_1.IRAM[59] [0], _07212_, clk);
  dff _54219_ (\uc8051golden_1.IRAM[59] [1], _07213_, clk);
  dff _54220_ (\uc8051golden_1.IRAM[59] [2], _07214_, clk);
  dff _54221_ (\uc8051golden_1.IRAM[59] [3], _07215_, clk);
  dff _54222_ (\uc8051golden_1.IRAM[59] [4], _07217_, clk);
  dff _54223_ (\uc8051golden_1.IRAM[59] [5], _07218_, clk);
  dff _54224_ (\uc8051golden_1.IRAM[59] [6], _07219_, clk);
  dff _54225_ (\uc8051golden_1.IRAM[59] [7], _07220_, clk);
  dff _54226_ (\uc8051golden_1.IRAM[60] [0], _07221_, clk);
  dff _54227_ (\uc8051golden_1.IRAM[60] [1], _07222_, clk);
  dff _54228_ (\uc8051golden_1.IRAM[60] [2], _07223_, clk);
  dff _54229_ (\uc8051golden_1.IRAM[60] [3], _07224_, clk);
  dff _54230_ (\uc8051golden_1.IRAM[60] [4], _07225_, clk);
  dff _54231_ (\uc8051golden_1.IRAM[60] [5], _07226_, clk);
  dff _54232_ (\uc8051golden_1.IRAM[60] [6], _07227_, clk);
  dff _54233_ (\uc8051golden_1.IRAM[60] [7], _07228_, clk);
  dff _54234_ (\uc8051golden_1.IRAM[61] [0], _07229_, clk);
  dff _54235_ (\uc8051golden_1.IRAM[61] [1], _07230_, clk);
  dff _54236_ (\uc8051golden_1.IRAM[61] [2], _07231_, clk);
  dff _54237_ (\uc8051golden_1.IRAM[61] [3], _07232_, clk);
  dff _54238_ (\uc8051golden_1.IRAM[61] [4], _07233_, clk);
  dff _54239_ (\uc8051golden_1.IRAM[61] [5], _07234_, clk);
  dff _54240_ (\uc8051golden_1.IRAM[61] [6], _07235_, clk);
  dff _54241_ (\uc8051golden_1.IRAM[61] [7], _07236_, clk);
  dff _54242_ (\uc8051golden_1.IRAM[62] [0], _07237_, clk);
  dff _54243_ (\uc8051golden_1.IRAM[62] [1], _07238_, clk);
  dff _54244_ (\uc8051golden_1.IRAM[62] [2], _07239_, clk);
  dff _54245_ (\uc8051golden_1.IRAM[62] [3], _07240_, clk);
  dff _54246_ (\uc8051golden_1.IRAM[62] [4], _07241_, clk);
  dff _54247_ (\uc8051golden_1.IRAM[62] [5], _07242_, clk);
  dff _54248_ (\uc8051golden_1.IRAM[62] [6], _07243_, clk);
  dff _54249_ (\uc8051golden_1.IRAM[62] [7], _07244_, clk);
  dff _54250_ (\uc8051golden_1.IRAM[63] [0], _07245_, clk);
  dff _54251_ (\uc8051golden_1.IRAM[63] [1], _07246_, clk);
  dff _54252_ (\uc8051golden_1.IRAM[63] [2], _07247_, clk);
  dff _54253_ (\uc8051golden_1.IRAM[63] [3], _07248_, clk);
  dff _54254_ (\uc8051golden_1.IRAM[63] [4], _07249_, clk);
  dff _54255_ (\uc8051golden_1.IRAM[63] [5], _07251_, clk);
  dff _54256_ (\uc8051golden_1.IRAM[63] [6], _07252_, clk);
  dff _54257_ (\uc8051golden_1.IRAM[63] [7], _07253_, clk);
  dff _54258_ (\uc8051golden_1.IRAM[64] [0], _07254_, clk);
  dff _54259_ (\uc8051golden_1.IRAM[64] [1], _07255_, clk);
  dff _54260_ (\uc8051golden_1.IRAM[64] [2], _07256_, clk);
  dff _54261_ (\uc8051golden_1.IRAM[64] [3], _07257_, clk);
  dff _54262_ (\uc8051golden_1.IRAM[64] [4], _07258_, clk);
  dff _54263_ (\uc8051golden_1.IRAM[64] [5], _07259_, clk);
  dff _54264_ (\uc8051golden_1.IRAM[64] [6], _07260_, clk);
  dff _54265_ (\uc8051golden_1.IRAM[64] [7], _07261_, clk);
  dff _54266_ (\uc8051golden_1.IRAM[65] [0], _07262_, clk);
  dff _54267_ (\uc8051golden_1.IRAM[65] [1], _07263_, clk);
  dff _54268_ (\uc8051golden_1.IRAM[65] [2], _07264_, clk);
  dff _54269_ (\uc8051golden_1.IRAM[65] [3], _07265_, clk);
  dff _54270_ (\uc8051golden_1.IRAM[65] [4], _07266_, clk);
  dff _54271_ (\uc8051golden_1.IRAM[65] [5], _07267_, clk);
  dff _54272_ (\uc8051golden_1.IRAM[65] [6], _07268_, clk);
  dff _54273_ (\uc8051golden_1.IRAM[65] [7], _07269_, clk);
  dff _54274_ (\uc8051golden_1.IRAM[66] [0], _07270_, clk);
  dff _54275_ (\uc8051golden_1.IRAM[66] [1], _07271_, clk);
  dff _54276_ (\uc8051golden_1.IRAM[66] [2], _07272_, clk);
  dff _54277_ (\uc8051golden_1.IRAM[66] [3], _07273_, clk);
  dff _54278_ (\uc8051golden_1.IRAM[66] [4], _07274_, clk);
  dff _54279_ (\uc8051golden_1.IRAM[66] [5], _07275_, clk);
  dff _54280_ (\uc8051golden_1.IRAM[66] [6], _07276_, clk);
  dff _54281_ (\uc8051golden_1.IRAM[66] [7], _07277_, clk);
  dff _54282_ (\uc8051golden_1.IRAM[67] [0], _07278_, clk);
  dff _54283_ (\uc8051golden_1.IRAM[67] [1], _07279_, clk);
  dff _54284_ (\uc8051golden_1.IRAM[67] [2], _07280_, clk);
  dff _54285_ (\uc8051golden_1.IRAM[67] [3], _07281_, clk);
  dff _54286_ (\uc8051golden_1.IRAM[67] [4], _07282_, clk);
  dff _54287_ (\uc8051golden_1.IRAM[67] [5], _07284_, clk);
  dff _54288_ (\uc8051golden_1.IRAM[67] [6], _07285_, clk);
  dff _54289_ (\uc8051golden_1.IRAM[67] [7], _07286_, clk);
  dff _54290_ (\uc8051golden_1.IRAM[68] [0], _07287_, clk);
  dff _54291_ (\uc8051golden_1.IRAM[68] [1], _07288_, clk);
  dff _54292_ (\uc8051golden_1.IRAM[68] [2], _07289_, clk);
  dff _54293_ (\uc8051golden_1.IRAM[68] [3], _07290_, clk);
  dff _54294_ (\uc8051golden_1.IRAM[68] [4], _07291_, clk);
  dff _54295_ (\uc8051golden_1.IRAM[68] [5], _07292_, clk);
  dff _54296_ (\uc8051golden_1.IRAM[68] [6], _07293_, clk);
  dff _54297_ (\uc8051golden_1.IRAM[68] [7], _07294_, clk);
  dff _54298_ (\uc8051golden_1.IRAM[69] [0], _07295_, clk);
  dff _54299_ (\uc8051golden_1.IRAM[69] [1], _07296_, clk);
  dff _54300_ (\uc8051golden_1.IRAM[69] [2], _07297_, clk);
  dff _54301_ (\uc8051golden_1.IRAM[69] [3], _07298_, clk);
  dff _54302_ (\uc8051golden_1.IRAM[69] [4], _07299_, clk);
  dff _54303_ (\uc8051golden_1.IRAM[69] [5], _07300_, clk);
  dff _54304_ (\uc8051golden_1.IRAM[69] [6], _07301_, clk);
  dff _54305_ (\uc8051golden_1.IRAM[69] [7], _07302_, clk);
  dff _54306_ (\uc8051golden_1.IRAM[70] [0], _07303_, clk);
  dff _54307_ (\uc8051golden_1.IRAM[70] [1], _07304_, clk);
  dff _54308_ (\uc8051golden_1.IRAM[70] [2], _07305_, clk);
  dff _54309_ (\uc8051golden_1.IRAM[70] [3], _07306_, clk);
  dff _54310_ (\uc8051golden_1.IRAM[70] [4], _07307_, clk);
  dff _54311_ (\uc8051golden_1.IRAM[70] [5], _07308_, clk);
  dff _54312_ (\uc8051golden_1.IRAM[70] [6], _07309_, clk);
  dff _54313_ (\uc8051golden_1.IRAM[70] [7], _07310_, clk);
  dff _54314_ (\uc8051golden_1.IRAM[71] [0], _07311_, clk);
  dff _54315_ (\uc8051golden_1.IRAM[71] [1], _07312_, clk);
  dff _54316_ (\uc8051golden_1.IRAM[71] [2], _07313_, clk);
  dff _54317_ (\uc8051golden_1.IRAM[71] [3], _07314_, clk);
  dff _54318_ (\uc8051golden_1.IRAM[71] [4], _07315_, clk);
  dff _54319_ (\uc8051golden_1.IRAM[71] [5], _07316_, clk);
  dff _54320_ (\uc8051golden_1.IRAM[71] [6], _07318_, clk);
  dff _54321_ (\uc8051golden_1.IRAM[71] [7], _07319_, clk);
  dff _54322_ (\uc8051golden_1.IRAM[72] [0], _07320_, clk);
  dff _54323_ (\uc8051golden_1.IRAM[72] [1], _07321_, clk);
  dff _54324_ (\uc8051golden_1.IRAM[72] [2], _07322_, clk);
  dff _54325_ (\uc8051golden_1.IRAM[72] [3], _07323_, clk);
  dff _54326_ (\uc8051golden_1.IRAM[72] [4], _07324_, clk);
  dff _54327_ (\uc8051golden_1.IRAM[72] [5], _07325_, clk);
  dff _54328_ (\uc8051golden_1.IRAM[72] [6], _07326_, clk);
  dff _54329_ (\uc8051golden_1.IRAM[72] [7], _07327_, clk);
  dff _54330_ (\uc8051golden_1.IRAM[73] [0], _07328_, clk);
  dff _54331_ (\uc8051golden_1.IRAM[73] [1], _07329_, clk);
  dff _54332_ (\uc8051golden_1.IRAM[73] [2], _07330_, clk);
  dff _54333_ (\uc8051golden_1.IRAM[73] [3], _07331_, clk);
  dff _54334_ (\uc8051golden_1.IRAM[73] [4], _07332_, clk);
  dff _54335_ (\uc8051golden_1.IRAM[73] [5], _07333_, clk);
  dff _54336_ (\uc8051golden_1.IRAM[73] [6], _07334_, clk);
  dff _54337_ (\uc8051golden_1.IRAM[73] [7], _07335_, clk);
  dff _54338_ (\uc8051golden_1.IRAM[74] [0], _07336_, clk);
  dff _54339_ (\uc8051golden_1.IRAM[74] [1], _07337_, clk);
  dff _54340_ (\uc8051golden_1.IRAM[74] [2], _07338_, clk);
  dff _54341_ (\uc8051golden_1.IRAM[74] [3], _07339_, clk);
  dff _54342_ (\uc8051golden_1.IRAM[74] [4], _07340_, clk);
  dff _54343_ (\uc8051golden_1.IRAM[74] [5], _07341_, clk);
  dff _54344_ (\uc8051golden_1.IRAM[74] [6], _07342_, clk);
  dff _54345_ (\uc8051golden_1.IRAM[74] [7], _07343_, clk);
  dff _54346_ (\uc8051golden_1.IRAM[75] [0], _07344_, clk);
  dff _54347_ (\uc8051golden_1.IRAM[75] [1], _07345_, clk);
  dff _54348_ (\uc8051golden_1.IRAM[75] [2], _07346_, clk);
  dff _54349_ (\uc8051golden_1.IRAM[75] [3], _07347_, clk);
  dff _54350_ (\uc8051golden_1.IRAM[75] [4], _07348_, clk);
  dff _54351_ (\uc8051golden_1.IRAM[75] [5], _07349_, clk);
  dff _54352_ (\uc8051golden_1.IRAM[75] [6], _07350_, clk);
  dff _54353_ (\uc8051golden_1.IRAM[75] [7], _07351_, clk);
  dff _54354_ (\uc8051golden_1.IRAM[76] [0], _07353_, clk);
  dff _54355_ (\uc8051golden_1.IRAM[76] [1], _07354_, clk);
  dff _54356_ (\uc8051golden_1.IRAM[76] [2], _07355_, clk);
  dff _54357_ (\uc8051golden_1.IRAM[76] [3], _07356_, clk);
  dff _54358_ (\uc8051golden_1.IRAM[76] [4], _07357_, clk);
  dff _54359_ (\uc8051golden_1.IRAM[76] [5], _07358_, clk);
  dff _54360_ (\uc8051golden_1.IRAM[76] [6], _07359_, clk);
  dff _54361_ (\uc8051golden_1.IRAM[76] [7], _07360_, clk);
  dff _54362_ (\uc8051golden_1.IRAM[77] [0], _07361_, clk);
  dff _54363_ (\uc8051golden_1.IRAM[77] [1], _07362_, clk);
  dff _54364_ (\uc8051golden_1.IRAM[77] [2], _07363_, clk);
  dff _54365_ (\uc8051golden_1.IRAM[77] [3], _07364_, clk);
  dff _54366_ (\uc8051golden_1.IRAM[77] [4], _07365_, clk);
  dff _54367_ (\uc8051golden_1.IRAM[77] [5], _07366_, clk);
  dff _54368_ (\uc8051golden_1.IRAM[77] [6], _07367_, clk);
  dff _54369_ (\uc8051golden_1.IRAM[77] [7], _07368_, clk);
  dff _54370_ (\uc8051golden_1.IRAM[78] [0], _07369_, clk);
  dff _54371_ (\uc8051golden_1.IRAM[78] [1], _07370_, clk);
  dff _54372_ (\uc8051golden_1.IRAM[78] [2], _07371_, clk);
  dff _54373_ (\uc8051golden_1.IRAM[78] [3], _07372_, clk);
  dff _54374_ (\uc8051golden_1.IRAM[78] [4], _07373_, clk);
  dff _54375_ (\uc8051golden_1.IRAM[78] [5], _07374_, clk);
  dff _54376_ (\uc8051golden_1.IRAM[78] [6], _07375_, clk);
  dff _54377_ (\uc8051golden_1.IRAM[78] [7], _07376_, clk);
  dff _54378_ (\uc8051golden_1.IRAM[79] [0], _07377_, clk);
  dff _54379_ (\uc8051golden_1.IRAM[79] [1], _07378_, clk);
  dff _54380_ (\uc8051golden_1.IRAM[79] [2], _07379_, clk);
  dff _54381_ (\uc8051golden_1.IRAM[79] [3], _07380_, clk);
  dff _54382_ (\uc8051golden_1.IRAM[79] [4], _07381_, clk);
  dff _54383_ (\uc8051golden_1.IRAM[79] [5], _07382_, clk);
  dff _54384_ (\uc8051golden_1.IRAM[79] [6], _07383_, clk);
  dff _54385_ (\uc8051golden_1.IRAM[79] [7], _07384_, clk);
  dff _54386_ (\uc8051golden_1.IRAM[80] [0], _07385_, clk);
  dff _54387_ (\uc8051golden_1.IRAM[80] [1], _07387_, clk);
  dff _54388_ (\uc8051golden_1.IRAM[80] [2], _07388_, clk);
  dff _54389_ (\uc8051golden_1.IRAM[80] [3], _07389_, clk);
  dff _54390_ (\uc8051golden_1.IRAM[80] [4], _07390_, clk);
  dff _54391_ (\uc8051golden_1.IRAM[80] [5], _07391_, clk);
  dff _54392_ (\uc8051golden_1.IRAM[80] [6], _07392_, clk);
  dff _54393_ (\uc8051golden_1.IRAM[80] [7], _07393_, clk);
  dff _54394_ (\uc8051golden_1.IRAM[81] [0], _07394_, clk);
  dff _54395_ (\uc8051golden_1.IRAM[81] [1], _07395_, clk);
  dff _54396_ (\uc8051golden_1.IRAM[81] [2], _07396_, clk);
  dff _54397_ (\uc8051golden_1.IRAM[81] [3], _07397_, clk);
  dff _54398_ (\uc8051golden_1.IRAM[81] [4], _07398_, clk);
  dff _54399_ (\uc8051golden_1.IRAM[81] [5], _07399_, clk);
  dff _54400_ (\uc8051golden_1.IRAM[81] [6], _07400_, clk);
  dff _54401_ (\uc8051golden_1.IRAM[81] [7], _07401_, clk);
  dff _54402_ (\uc8051golden_1.IRAM[82] [0], _07402_, clk);
  dff _54403_ (\uc8051golden_1.IRAM[82] [1], _07403_, clk);
  dff _54404_ (\uc8051golden_1.IRAM[82] [2], _07404_, clk);
  dff _54405_ (\uc8051golden_1.IRAM[82] [3], _07405_, clk);
  dff _54406_ (\uc8051golden_1.IRAM[82] [4], _07406_, clk);
  dff _54407_ (\uc8051golden_1.IRAM[82] [5], _07407_, clk);
  dff _54408_ (\uc8051golden_1.IRAM[82] [6], _07408_, clk);
  dff _54409_ (\uc8051golden_1.IRAM[82] [7], _07409_, clk);
  dff _54410_ (\uc8051golden_1.IRAM[83] [0], _07410_, clk);
  dff _54411_ (\uc8051golden_1.IRAM[83] [1], _07411_, clk);
  dff _54412_ (\uc8051golden_1.IRAM[83] [2], _07412_, clk);
  dff _54413_ (\uc8051golden_1.IRAM[83] [3], _07413_, clk);
  dff _54414_ (\uc8051golden_1.IRAM[83] [4], _07414_, clk);
  dff _54415_ (\uc8051golden_1.IRAM[83] [5], _07415_, clk);
  dff _54416_ (\uc8051golden_1.IRAM[83] [6], _07416_, clk);
  dff _54417_ (\uc8051golden_1.IRAM[83] [7], _07417_, clk);
  dff _54418_ (\uc8051golden_1.IRAM[84] [0], _07418_, clk);
  dff _54419_ (\uc8051golden_1.IRAM[84] [1], _07419_, clk);
  dff _54420_ (\uc8051golden_1.IRAM[84] [2], _07421_, clk);
  dff _54421_ (\uc8051golden_1.IRAM[84] [3], _07422_, clk);
  dff _54422_ (\uc8051golden_1.IRAM[84] [4], _07423_, clk);
  dff _54423_ (\uc8051golden_1.IRAM[84] [5], _07424_, clk);
  dff _54424_ (\uc8051golden_1.IRAM[84] [6], _07425_, clk);
  dff _54425_ (\uc8051golden_1.IRAM[84] [7], _07426_, clk);
  dff _54426_ (\uc8051golden_1.IRAM[85] [0], _07427_, clk);
  dff _54427_ (\uc8051golden_1.IRAM[85] [1], _07428_, clk);
  dff _54428_ (\uc8051golden_1.IRAM[85] [2], _07429_, clk);
  dff _54429_ (\uc8051golden_1.IRAM[85] [3], _07430_, clk);
  dff _54430_ (\uc8051golden_1.IRAM[85] [4], _07431_, clk);
  dff _54431_ (\uc8051golden_1.IRAM[85] [5], _07432_, clk);
  dff _54432_ (\uc8051golden_1.IRAM[85] [6], _07433_, clk);
  dff _54433_ (\uc8051golden_1.IRAM[85] [7], _07434_, clk);
  dff _54434_ (\uc8051golden_1.IRAM[86] [0], _07435_, clk);
  dff _54435_ (\uc8051golden_1.IRAM[86] [1], _07436_, clk);
  dff _54436_ (\uc8051golden_1.IRAM[86] [2], _07437_, clk);
  dff _54437_ (\uc8051golden_1.IRAM[86] [3], _07438_, clk);
  dff _54438_ (\uc8051golden_1.IRAM[86] [4], _07439_, clk);
  dff _54439_ (\uc8051golden_1.IRAM[86] [5], _07440_, clk);
  dff _54440_ (\uc8051golden_1.IRAM[86] [6], _07441_, clk);
  dff _54441_ (\uc8051golden_1.IRAM[86] [7], _07442_, clk);
  dff _54442_ (\uc8051golden_1.IRAM[87] [0], _07443_, clk);
  dff _54443_ (\uc8051golden_1.IRAM[87] [1], _07444_, clk);
  dff _54444_ (\uc8051golden_1.IRAM[87] [2], _07445_, clk);
  dff _54445_ (\uc8051golden_1.IRAM[87] [3], _07446_, clk);
  dff _54446_ (\uc8051golden_1.IRAM[87] [4], _07447_, clk);
  dff _54447_ (\uc8051golden_1.IRAM[87] [5], _07448_, clk);
  dff _54448_ (\uc8051golden_1.IRAM[87] [6], _07449_, clk);
  dff _54449_ (\uc8051golden_1.IRAM[87] [7], _07450_, clk);
  dff _54450_ (\uc8051golden_1.IRAM[88] [0], _07451_, clk);
  dff _54451_ (\uc8051golden_1.IRAM[88] [1], _07452_, clk);
  dff _54452_ (\uc8051golden_1.IRAM[88] [2], _07453_, clk);
  dff _54453_ (\uc8051golden_1.IRAM[88] [3], _07455_, clk);
  dff _54454_ (\uc8051golden_1.IRAM[88] [4], _07456_, clk);
  dff _54455_ (\uc8051golden_1.IRAM[88] [5], _07457_, clk);
  dff _54456_ (\uc8051golden_1.IRAM[88] [6], _07458_, clk);
  dff _54457_ (\uc8051golden_1.IRAM[88] [7], _07459_, clk);
  dff _54458_ (\uc8051golden_1.IRAM[89] [0], _07460_, clk);
  dff _54459_ (\uc8051golden_1.IRAM[89] [1], _07461_, clk);
  dff _54460_ (\uc8051golden_1.IRAM[89] [2], _07462_, clk);
  dff _54461_ (\uc8051golden_1.IRAM[89] [3], _07463_, clk);
  dff _54462_ (\uc8051golden_1.IRAM[89] [4], _07464_, clk);
  dff _54463_ (\uc8051golden_1.IRAM[89] [5], _07465_, clk);
  dff _54464_ (\uc8051golden_1.IRAM[89] [6], _07466_, clk);
  dff _54465_ (\uc8051golden_1.IRAM[89] [7], _07467_, clk);
  dff _54466_ (\uc8051golden_1.IRAM[90] [0], _07468_, clk);
  dff _54467_ (\uc8051golden_1.IRAM[90] [1], _07469_, clk);
  dff _54468_ (\uc8051golden_1.IRAM[90] [2], _07470_, clk);
  dff _54469_ (\uc8051golden_1.IRAM[90] [3], _07471_, clk);
  dff _54470_ (\uc8051golden_1.IRAM[90] [4], _07472_, clk);
  dff _54471_ (\uc8051golden_1.IRAM[90] [5], _07473_, clk);
  dff _54472_ (\uc8051golden_1.IRAM[90] [6], _07474_, clk);
  dff _54473_ (\uc8051golden_1.IRAM[90] [7], _07475_, clk);
  dff _54474_ (\uc8051golden_1.IRAM[91] [0], _07476_, clk);
  dff _54475_ (\uc8051golden_1.IRAM[91] [1], _07477_, clk);
  dff _54476_ (\uc8051golden_1.IRAM[91] [2], _07478_, clk);
  dff _54477_ (\uc8051golden_1.IRAM[91] [3], _07479_, clk);
  dff _54478_ (\uc8051golden_1.IRAM[91] [4], _07480_, clk);
  dff _54479_ (\uc8051golden_1.IRAM[91] [5], _07481_, clk);
  dff _54480_ (\uc8051golden_1.IRAM[91] [6], _07482_, clk);
  dff _54481_ (\uc8051golden_1.IRAM[91] [7], _07483_, clk);
  dff _54482_ (\uc8051golden_1.IRAM[92] [0], _07484_, clk);
  dff _54483_ (\uc8051golden_1.IRAM[92] [1], _07485_, clk);
  dff _54484_ (\uc8051golden_1.IRAM[92] [2], _07486_, clk);
  dff _54485_ (\uc8051golden_1.IRAM[92] [3], _07487_, clk);
  dff _54486_ (\uc8051golden_1.IRAM[92] [4], _07488_, clk);
  dff _54487_ (\uc8051golden_1.IRAM[92] [5], _07490_, clk);
  dff _54488_ (\uc8051golden_1.IRAM[92] [6], _07491_, clk);
  dff _54489_ (\uc8051golden_1.IRAM[92] [7], _07492_, clk);
  dff _54490_ (\uc8051golden_1.IRAM[93] [0], _07493_, clk);
  dff _54491_ (\uc8051golden_1.IRAM[93] [1], _07494_, clk);
  dff _54492_ (\uc8051golden_1.IRAM[93] [2], _07495_, clk);
  dff _54493_ (\uc8051golden_1.IRAM[93] [3], _07496_, clk);
  dff _54494_ (\uc8051golden_1.IRAM[93] [4], _07497_, clk);
  dff _54495_ (\uc8051golden_1.IRAM[93] [5], _07498_, clk);
  dff _54496_ (\uc8051golden_1.IRAM[93] [6], _07499_, clk);
  dff _54497_ (\uc8051golden_1.IRAM[93] [7], _07500_, clk);
  dff _54498_ (\uc8051golden_1.IRAM[94] [0], _07501_, clk);
  dff _54499_ (\uc8051golden_1.IRAM[94] [1], _07502_, clk);
  dff _54500_ (\uc8051golden_1.IRAM[94] [2], _07503_, clk);
  dff _54501_ (\uc8051golden_1.IRAM[94] [3], _07504_, clk);
  dff _54502_ (\uc8051golden_1.IRAM[94] [4], _07505_, clk);
  dff _54503_ (\uc8051golden_1.IRAM[94] [5], _07506_, clk);
  dff _54504_ (\uc8051golden_1.IRAM[94] [6], _07507_, clk);
  dff _54505_ (\uc8051golden_1.IRAM[94] [7], _07508_, clk);
  dff _54506_ (\uc8051golden_1.IRAM[95] [0], _07509_, clk);
  dff _54507_ (\uc8051golden_1.IRAM[95] [1], _07510_, clk);
  dff _54508_ (\uc8051golden_1.IRAM[95] [2], _07511_, clk);
  dff _54509_ (\uc8051golden_1.IRAM[95] [3], _07512_, clk);
  dff _54510_ (\uc8051golden_1.IRAM[95] [4], _07513_, clk);
  dff _54511_ (\uc8051golden_1.IRAM[95] [5], _07514_, clk);
  dff _54512_ (\uc8051golden_1.IRAM[95] [6], _07515_, clk);
  dff _54513_ (\uc8051golden_1.IRAM[95] [7], _07516_, clk);
  dff _54514_ (\uc8051golden_1.IRAM[96] [0], _07517_, clk);
  dff _54515_ (\uc8051golden_1.IRAM[96] [1], _07518_, clk);
  dff _54516_ (\uc8051golden_1.IRAM[96] [2], _07519_, clk);
  dff _54517_ (\uc8051golden_1.IRAM[96] [3], _07520_, clk);
  dff _54518_ (\uc8051golden_1.IRAM[96] [4], _07521_, clk);
  dff _54519_ (\uc8051golden_1.IRAM[96] [5], _07522_, clk);
  dff _54520_ (\uc8051golden_1.IRAM[96] [6], _07524_, clk);
  dff _54521_ (\uc8051golden_1.IRAM[96] [7], _07525_, clk);
  dff _54522_ (\uc8051golden_1.IRAM[97] [0], _07526_, clk);
  dff _54523_ (\uc8051golden_1.IRAM[97] [1], _07527_, clk);
  dff _54524_ (\uc8051golden_1.IRAM[97] [2], _07528_, clk);
  dff _54525_ (\uc8051golden_1.IRAM[97] [3], _07529_, clk);
  dff _54526_ (\uc8051golden_1.IRAM[97] [4], _07530_, clk);
  dff _54527_ (\uc8051golden_1.IRAM[97] [5], _07531_, clk);
  dff _54528_ (\uc8051golden_1.IRAM[97] [6], _07532_, clk);
  dff _54529_ (\uc8051golden_1.IRAM[97] [7], _07533_, clk);
  dff _54530_ (\uc8051golden_1.IRAM[98] [0], _07534_, clk);
  dff _54531_ (\uc8051golden_1.IRAM[98] [1], _07535_, clk);
  dff _54532_ (\uc8051golden_1.IRAM[98] [2], _07536_, clk);
  dff _54533_ (\uc8051golden_1.IRAM[98] [3], _07537_, clk);
  dff _54534_ (\uc8051golden_1.IRAM[98] [4], _07538_, clk);
  dff _54535_ (\uc8051golden_1.IRAM[98] [5], _07539_, clk);
  dff _54536_ (\uc8051golden_1.IRAM[98] [6], _07540_, clk);
  dff _54537_ (\uc8051golden_1.IRAM[98] [7], _07541_, clk);
  dff _54538_ (\uc8051golden_1.IRAM[99] [0], _07542_, clk);
  dff _54539_ (\uc8051golden_1.IRAM[99] [1], _07543_, clk);
  dff _54540_ (\uc8051golden_1.IRAM[99] [2], _07544_, clk);
  dff _54541_ (\uc8051golden_1.IRAM[99] [3], _07545_, clk);
  dff _54542_ (\uc8051golden_1.IRAM[99] [4], _07546_, clk);
  dff _54543_ (\uc8051golden_1.IRAM[99] [5], _07547_, clk);
  dff _54544_ (\uc8051golden_1.IRAM[99] [6], _07548_, clk);
  dff _54545_ (\uc8051golden_1.IRAM[99] [7], _07549_, clk);
  dff _54546_ (\uc8051golden_1.IRAM[100] [0], _07550_, clk);
  dff _54547_ (\uc8051golden_1.IRAM[100] [1], _07551_, clk);
  dff _54548_ (\uc8051golden_1.IRAM[100] [2], _07552_, clk);
  dff _54549_ (\uc8051golden_1.IRAM[100] [3], _07553_, clk);
  dff _54550_ (\uc8051golden_1.IRAM[100] [4], _07554_, clk);
  dff _54551_ (\uc8051golden_1.IRAM[100] [5], _07555_, clk);
  dff _54552_ (\uc8051golden_1.IRAM[100] [6], _07556_, clk);
  dff _54553_ (\uc8051golden_1.IRAM[100] [7], _07558_, clk);
  dff _54554_ (\uc8051golden_1.IRAM[101] [0], _07559_, clk);
  dff _54555_ (\uc8051golden_1.IRAM[101] [1], _07560_, clk);
  dff _54556_ (\uc8051golden_1.IRAM[101] [2], _07561_, clk);
  dff _54557_ (\uc8051golden_1.IRAM[101] [3], _07562_, clk);
  dff _54558_ (\uc8051golden_1.IRAM[101] [4], _07563_, clk);
  dff _54559_ (\uc8051golden_1.IRAM[101] [5], _07564_, clk);
  dff _54560_ (\uc8051golden_1.IRAM[101] [6], _07565_, clk);
  dff _54561_ (\uc8051golden_1.IRAM[101] [7], _07566_, clk);
  dff _54562_ (\uc8051golden_1.IRAM[102] [0], _07567_, clk);
  dff _54563_ (\uc8051golden_1.IRAM[102] [1], _07568_, clk);
  dff _54564_ (\uc8051golden_1.IRAM[102] [2], _07569_, clk);
  dff _54565_ (\uc8051golden_1.IRAM[102] [3], _07570_, clk);
  dff _54566_ (\uc8051golden_1.IRAM[102] [4], _07571_, clk);
  dff _54567_ (\uc8051golden_1.IRAM[102] [5], _07572_, clk);
  dff _54568_ (\uc8051golden_1.IRAM[102] [6], _07573_, clk);
  dff _54569_ (\uc8051golden_1.IRAM[102] [7], _07574_, clk);
  dff _54570_ (\uc8051golden_1.IRAM[103] [0], _07575_, clk);
  dff _54571_ (\uc8051golden_1.IRAM[103] [1], _07576_, clk);
  dff _54572_ (\uc8051golden_1.IRAM[103] [2], _07577_, clk);
  dff _54573_ (\uc8051golden_1.IRAM[103] [3], _07578_, clk);
  dff _54574_ (\uc8051golden_1.IRAM[103] [4], _07579_, clk);
  dff _54575_ (\uc8051golden_1.IRAM[103] [5], _07580_, clk);
  dff _54576_ (\uc8051golden_1.IRAM[103] [6], _07581_, clk);
  dff _54577_ (\uc8051golden_1.IRAM[103] [7], _07582_, clk);
  dff _54578_ (\uc8051golden_1.IRAM[104] [0], _07583_, clk);
  dff _54579_ (\uc8051golden_1.IRAM[104] [1], _07584_, clk);
  dff _54580_ (\uc8051golden_1.IRAM[104] [2], _07585_, clk);
  dff _54581_ (\uc8051golden_1.IRAM[104] [3], _07586_, clk);
  dff _54582_ (\uc8051golden_1.IRAM[104] [4], _07587_, clk);
  dff _54583_ (\uc8051golden_1.IRAM[104] [5], _07588_, clk);
  dff _54584_ (\uc8051golden_1.IRAM[104] [6], _07589_, clk);
  dff _54585_ (\uc8051golden_1.IRAM[104] [7], _07590_, clk);
  dff _54586_ (\uc8051golden_1.IRAM[105] [0], _07592_, clk);
  dff _54587_ (\uc8051golden_1.IRAM[105] [1], _07593_, clk);
  dff _54588_ (\uc8051golden_1.IRAM[105] [2], _07594_, clk);
  dff _54589_ (\uc8051golden_1.IRAM[105] [3], _07595_, clk);
  dff _54590_ (\uc8051golden_1.IRAM[105] [4], _07596_, clk);
  dff _54591_ (\uc8051golden_1.IRAM[105] [5], _07597_, clk);
  dff _54592_ (\uc8051golden_1.IRAM[105] [6], _07598_, clk);
  dff _54593_ (\uc8051golden_1.IRAM[105] [7], _07599_, clk);
  dff _54594_ (\uc8051golden_1.IRAM[106] [0], _07600_, clk);
  dff _54595_ (\uc8051golden_1.IRAM[106] [1], _07601_, clk);
  dff _54596_ (\uc8051golden_1.IRAM[106] [2], _07602_, clk);
  dff _54597_ (\uc8051golden_1.IRAM[106] [3], _07603_, clk);
  dff _54598_ (\uc8051golden_1.IRAM[106] [4], _07604_, clk);
  dff _54599_ (\uc8051golden_1.IRAM[106] [5], _07605_, clk);
  dff _54600_ (\uc8051golden_1.IRAM[106] [6], _07606_, clk);
  dff _54601_ (\uc8051golden_1.IRAM[106] [7], _07607_, clk);
  dff _54602_ (\uc8051golden_1.IRAM[107] [0], _07608_, clk);
  dff _54603_ (\uc8051golden_1.IRAM[107] [1], _07609_, clk);
  dff _54604_ (\uc8051golden_1.IRAM[107] [2], _07610_, clk);
  dff _54605_ (\uc8051golden_1.IRAM[107] [3], _07611_, clk);
  dff _54606_ (\uc8051golden_1.IRAM[107] [4], _07612_, clk);
  dff _54607_ (\uc8051golden_1.IRAM[107] [5], _07613_, clk);
  dff _54608_ (\uc8051golden_1.IRAM[107] [6], _07614_, clk);
  dff _54609_ (\uc8051golden_1.IRAM[107] [7], _07615_, clk);
  dff _54610_ (\uc8051golden_1.IRAM[108] [0], _07616_, clk);
  dff _54611_ (\uc8051golden_1.IRAM[108] [1], _07617_, clk);
  dff _54612_ (\uc8051golden_1.IRAM[108] [2], _07618_, clk);
  dff _54613_ (\uc8051golden_1.IRAM[108] [3], _07619_, clk);
  dff _54614_ (\uc8051golden_1.IRAM[108] [4], _07620_, clk);
  dff _54615_ (\uc8051golden_1.IRAM[108] [5], _07621_, clk);
  dff _54616_ (\uc8051golden_1.IRAM[108] [6], _07622_, clk);
  dff _54617_ (\uc8051golden_1.IRAM[108] [7], _07623_, clk);
  dff _54618_ (\uc8051golden_1.IRAM[109] [0], _07624_, clk);
  dff _54619_ (\uc8051golden_1.IRAM[109] [1], _07625_, clk);
  dff _54620_ (\uc8051golden_1.IRAM[109] [2], _07627_, clk);
  dff _54621_ (\uc8051golden_1.IRAM[109] [3], _07628_, clk);
  dff _54622_ (\uc8051golden_1.IRAM[109] [4], _07629_, clk);
  dff _54623_ (\uc8051golden_1.IRAM[109] [5], _07630_, clk);
  dff _54624_ (\uc8051golden_1.IRAM[109] [6], _07631_, clk);
  dff _54625_ (\uc8051golden_1.IRAM[109] [7], _07632_, clk);
  dff _54626_ (\uc8051golden_1.IRAM[110] [0], _07633_, clk);
  dff _54627_ (\uc8051golden_1.IRAM[110] [1], _07634_, clk);
  dff _54628_ (\uc8051golden_1.IRAM[110] [2], _07635_, clk);
  dff _54629_ (\uc8051golden_1.IRAM[110] [3], _07636_, clk);
  dff _54630_ (\uc8051golden_1.IRAM[110] [4], _07637_, clk);
  dff _54631_ (\uc8051golden_1.IRAM[110] [5], _07638_, clk);
  dff _54632_ (\uc8051golden_1.IRAM[110] [6], _07639_, clk);
  dff _54633_ (\uc8051golden_1.IRAM[110] [7], _07640_, clk);
  dff _54634_ (\uc8051golden_1.IRAM[111] [0], _07641_, clk);
  dff _54635_ (\uc8051golden_1.IRAM[111] [1], _07642_, clk);
  dff _54636_ (\uc8051golden_1.IRAM[111] [2], _07643_, clk);
  dff _54637_ (\uc8051golden_1.IRAM[111] [3], _07644_, clk);
  dff _54638_ (\uc8051golden_1.IRAM[111] [4], _07645_, clk);
  dff _54639_ (\uc8051golden_1.IRAM[111] [5], _07646_, clk);
  dff _54640_ (\uc8051golden_1.IRAM[111] [6], _07647_, clk);
  dff _54641_ (\uc8051golden_1.IRAM[111] [7], _07648_, clk);
  dff _54642_ (\uc8051golden_1.IRAM[112] [0], _07649_, clk);
  dff _54643_ (\uc8051golden_1.IRAM[112] [1], _07650_, clk);
  dff _54644_ (\uc8051golden_1.IRAM[112] [2], _07651_, clk);
  dff _54645_ (\uc8051golden_1.IRAM[112] [3], _07652_, clk);
  dff _54646_ (\uc8051golden_1.IRAM[112] [4], _07653_, clk);
  dff _54647_ (\uc8051golden_1.IRAM[112] [5], _07654_, clk);
  dff _54648_ (\uc8051golden_1.IRAM[112] [6], _07655_, clk);
  dff _54649_ (\uc8051golden_1.IRAM[112] [7], _07656_, clk);
  dff _54650_ (\uc8051golden_1.IRAM[113] [0], _07657_, clk);
  dff _54651_ (\uc8051golden_1.IRAM[113] [1], _07658_, clk);
  dff _54652_ (\uc8051golden_1.IRAM[113] [2], _07659_, clk);
  dff _54653_ (\uc8051golden_1.IRAM[113] [3], _07661_, clk);
  dff _54654_ (\uc8051golden_1.IRAM[113] [4], _07662_, clk);
  dff _54655_ (\uc8051golden_1.IRAM[113] [5], _07663_, clk);
  dff _54656_ (\uc8051golden_1.IRAM[113] [6], _07664_, clk);
  dff _54657_ (\uc8051golden_1.IRAM[113] [7], _07665_, clk);
  dff _54658_ (\uc8051golden_1.IRAM[114] [0], _07666_, clk);
  dff _54659_ (\uc8051golden_1.IRAM[114] [1], _07667_, clk);
  dff _54660_ (\uc8051golden_1.IRAM[114] [2], _07668_, clk);
  dff _54661_ (\uc8051golden_1.IRAM[114] [3], _07669_, clk);
  dff _54662_ (\uc8051golden_1.IRAM[114] [4], _07670_, clk);
  dff _54663_ (\uc8051golden_1.IRAM[114] [5], _07671_, clk);
  dff _54664_ (\uc8051golden_1.IRAM[114] [6], _07672_, clk);
  dff _54665_ (\uc8051golden_1.IRAM[114] [7], _07673_, clk);
  dff _54666_ (\uc8051golden_1.IRAM[115] [0], _07674_, clk);
  dff _54667_ (\uc8051golden_1.IRAM[115] [1], _07675_, clk);
  dff _54668_ (\uc8051golden_1.IRAM[115] [2], _07676_, clk);
  dff _54669_ (\uc8051golden_1.IRAM[115] [3], _07677_, clk);
  dff _54670_ (\uc8051golden_1.IRAM[115] [4], _07678_, clk);
  dff _54671_ (\uc8051golden_1.IRAM[115] [5], _07679_, clk);
  dff _54672_ (\uc8051golden_1.IRAM[115] [6], _07680_, clk);
  dff _54673_ (\uc8051golden_1.IRAM[115] [7], _07681_, clk);
  dff _54674_ (\uc8051golden_1.IRAM[116] [0], _07682_, clk);
  dff _54675_ (\uc8051golden_1.IRAM[116] [1], _07683_, clk);
  dff _54676_ (\uc8051golden_1.IRAM[116] [2], _07684_, clk);
  dff _54677_ (\uc8051golden_1.IRAM[116] [3], _07685_, clk);
  dff _54678_ (\uc8051golden_1.IRAM[116] [4], _07686_, clk);
  dff _54679_ (\uc8051golden_1.IRAM[116] [5], _07687_, clk);
  dff _54680_ (\uc8051golden_1.IRAM[116] [6], _07688_, clk);
  dff _54681_ (\uc8051golden_1.IRAM[116] [7], _07689_, clk);
  dff _54682_ (\uc8051golden_1.IRAM[117] [0], _07690_, clk);
  dff _54683_ (\uc8051golden_1.IRAM[117] [1], _07691_, clk);
  dff _54684_ (\uc8051golden_1.IRAM[117] [2], _07692_, clk);
  dff _54685_ (\uc8051golden_1.IRAM[117] [3], _07693_, clk);
  dff _54686_ (\uc8051golden_1.IRAM[117] [4], _07695_, clk);
  dff _54687_ (\uc8051golden_1.IRAM[117] [5], _07696_, clk);
  dff _54688_ (\uc8051golden_1.IRAM[117] [6], _07697_, clk);
  dff _54689_ (\uc8051golden_1.IRAM[117] [7], _07698_, clk);
  dff _54690_ (\uc8051golden_1.IRAM[118] [0], _07699_, clk);
  dff _54691_ (\uc8051golden_1.IRAM[118] [1], _07700_, clk);
  dff _54692_ (\uc8051golden_1.IRAM[118] [2], _07701_, clk);
  dff _54693_ (\uc8051golden_1.IRAM[118] [3], _07702_, clk);
  dff _54694_ (\uc8051golden_1.IRAM[118] [4], _07703_, clk);
  dff _54695_ (\uc8051golden_1.IRAM[118] [5], _07704_, clk);
  dff _54696_ (\uc8051golden_1.IRAM[118] [6], _07705_, clk);
  dff _54697_ (\uc8051golden_1.IRAM[118] [7], _07706_, clk);
  dff _54698_ (\uc8051golden_1.IRAM[119] [0], _07707_, clk);
  dff _54699_ (\uc8051golden_1.IRAM[119] [1], _07708_, clk);
  dff _54700_ (\uc8051golden_1.IRAM[119] [2], _07709_, clk);
  dff _54701_ (\uc8051golden_1.IRAM[119] [3], _07710_, clk);
  dff _54702_ (\uc8051golden_1.IRAM[119] [4], _07711_, clk);
  dff _54703_ (\uc8051golden_1.IRAM[119] [5], _07712_, clk);
  dff _54704_ (\uc8051golden_1.IRAM[119] [6], _07713_, clk);
  dff _54705_ (\uc8051golden_1.IRAM[119] [7], _07714_, clk);
  dff _54706_ (\uc8051golden_1.IRAM[120] [0], _07715_, clk);
  dff _54707_ (\uc8051golden_1.IRAM[120] [1], _07716_, clk);
  dff _54708_ (\uc8051golden_1.IRAM[120] [2], _07717_, clk);
  dff _54709_ (\uc8051golden_1.IRAM[120] [3], _07718_, clk);
  dff _54710_ (\uc8051golden_1.IRAM[120] [4], _07719_, clk);
  dff _54711_ (\uc8051golden_1.IRAM[120] [5], _07720_, clk);
  dff _54712_ (\uc8051golden_1.IRAM[120] [6], _07721_, clk);
  dff _54713_ (\uc8051golden_1.IRAM[120] [7], _07722_, clk);
  dff _54714_ (\uc8051golden_1.IRAM[121] [0], _07723_, clk);
  dff _54715_ (\uc8051golden_1.IRAM[121] [1], _07724_, clk);
  dff _54716_ (\uc8051golden_1.IRAM[121] [2], _07725_, clk);
  dff _54717_ (\uc8051golden_1.IRAM[121] [3], _07726_, clk);
  dff _54718_ (\uc8051golden_1.IRAM[121] [4], _07727_, clk);
  dff _54719_ (\uc8051golden_1.IRAM[121] [5], _07729_, clk);
  dff _54720_ (\uc8051golden_1.IRAM[121] [6], _07730_, clk);
  dff _54721_ (\uc8051golden_1.IRAM[121] [7], _07731_, clk);
  dff _54722_ (\uc8051golden_1.IRAM[122] [0], _07732_, clk);
  dff _54723_ (\uc8051golden_1.IRAM[122] [1], _07733_, clk);
  dff _54724_ (\uc8051golden_1.IRAM[122] [2], _07734_, clk);
  dff _54725_ (\uc8051golden_1.IRAM[122] [3], _07735_, clk);
  dff _54726_ (\uc8051golden_1.IRAM[122] [4], _07736_, clk);
  dff _54727_ (\uc8051golden_1.IRAM[122] [5], _07737_, clk);
  dff _54728_ (\uc8051golden_1.IRAM[122] [6], _07738_, clk);
  dff _54729_ (\uc8051golden_1.IRAM[122] [7], _07739_, clk);
  dff _54730_ (\uc8051golden_1.IRAM[123] [0], _07740_, clk);
  dff _54731_ (\uc8051golden_1.IRAM[123] [1], _07741_, clk);
  dff _54732_ (\uc8051golden_1.IRAM[123] [2], _07742_, clk);
  dff _54733_ (\uc8051golden_1.IRAM[123] [3], _07743_, clk);
  dff _54734_ (\uc8051golden_1.IRAM[123] [4], _07744_, clk);
  dff _54735_ (\uc8051golden_1.IRAM[123] [5], _07745_, clk);
  dff _54736_ (\uc8051golden_1.IRAM[123] [6], _07746_, clk);
  dff _54737_ (\uc8051golden_1.IRAM[123] [7], _07747_, clk);
  dff _54738_ (\uc8051golden_1.IRAM[124] [0], _07748_, clk);
  dff _54739_ (\uc8051golden_1.IRAM[124] [1], _07749_, clk);
  dff _54740_ (\uc8051golden_1.IRAM[124] [2], _07750_, clk);
  dff _54741_ (\uc8051golden_1.IRAM[124] [3], _07751_, clk);
  dff _54742_ (\uc8051golden_1.IRAM[124] [4], _07752_, clk);
  dff _54743_ (\uc8051golden_1.IRAM[124] [5], _07753_, clk);
  dff _54744_ (\uc8051golden_1.IRAM[124] [6], _07754_, clk);
  dff _54745_ (\uc8051golden_1.IRAM[124] [7], _07755_, clk);
  dff _54746_ (\uc8051golden_1.IRAM[125] [0], _07756_, clk);
  dff _54747_ (\uc8051golden_1.IRAM[125] [1], _07757_, clk);
  dff _54748_ (\uc8051golden_1.IRAM[125] [2], _07758_, clk);
  dff _54749_ (\uc8051golden_1.IRAM[125] [3], _07759_, clk);
  dff _54750_ (\uc8051golden_1.IRAM[125] [4], _07760_, clk);
  dff _54751_ (\uc8051golden_1.IRAM[125] [5], _07761_, clk);
  dff _54752_ (\uc8051golden_1.IRAM[125] [6], _07762_, clk);
  dff _54753_ (\uc8051golden_1.IRAM[125] [7], _07764_, clk);
  dff _54754_ (\uc8051golden_1.IRAM[126] [0], _07765_, clk);
  dff _54755_ (\uc8051golden_1.IRAM[126] [1], _07766_, clk);
  dff _54756_ (\uc8051golden_1.IRAM[126] [2], _07767_, clk);
  dff _54757_ (\uc8051golden_1.IRAM[126] [3], _07768_, clk);
  dff _54758_ (\uc8051golden_1.IRAM[126] [4], _07769_, clk);
  dff _54759_ (\uc8051golden_1.IRAM[126] [5], _07770_, clk);
  dff _54760_ (\uc8051golden_1.IRAM[126] [6], _07771_, clk);
  dff _54761_ (\uc8051golden_1.IRAM[126] [7], _07772_, clk);
  dff _54762_ (\uc8051golden_1.IRAM[127] [0], _07773_, clk);
  dff _54763_ (\uc8051golden_1.IRAM[127] [1], _07774_, clk);
  dff _54764_ (\uc8051golden_1.IRAM[127] [2], _07775_, clk);
  dff _54765_ (\uc8051golden_1.IRAM[127] [3], _07776_, clk);
  dff _54766_ (\uc8051golden_1.IRAM[127] [4], _07777_, clk);
  dff _54767_ (\uc8051golden_1.IRAM[127] [5], _07778_, clk);
  dff _54768_ (\uc8051golden_1.IRAM[127] [6], _07779_, clk);
  dff _54769_ (\uc8051golden_1.IRAM[127] [7], _07780_, clk);
  dff _54770_ (\uc8051golden_1.IRAM[128] [0], _07781_, clk);
  dff _54771_ (\uc8051golden_1.IRAM[128] [1], _07782_, clk);
  dff _54772_ (\uc8051golden_1.IRAM[128] [2], _07783_, clk);
  dff _54773_ (\uc8051golden_1.IRAM[128] [3], _07784_, clk);
  dff _54774_ (\uc8051golden_1.IRAM[128] [4], _07785_, clk);
  dff _54775_ (\uc8051golden_1.IRAM[128] [5], _07786_, clk);
  dff _54776_ (\uc8051golden_1.IRAM[128] [6], _07787_, clk);
  dff _54777_ (\uc8051golden_1.IRAM[128] [7], _07788_, clk);
  dff _54778_ (\uc8051golden_1.IRAM[129] [0], _07789_, clk);
  dff _54779_ (\uc8051golden_1.IRAM[129] [1], _07790_, clk);
  dff _54780_ (\uc8051golden_1.IRAM[129] [2], _07791_, clk);
  dff _54781_ (\uc8051golden_1.IRAM[129] [3], _07792_, clk);
  dff _54782_ (\uc8051golden_1.IRAM[129] [4], _07793_, clk);
  dff _54783_ (\uc8051golden_1.IRAM[129] [5], _07794_, clk);
  dff _54784_ (\uc8051golden_1.IRAM[129] [6], _07795_, clk);
  dff _54785_ (\uc8051golden_1.IRAM[129] [7], _07797_, clk);
  dff _54786_ (\uc8051golden_1.IRAM[130] [0], _07798_, clk);
  dff _54787_ (\uc8051golden_1.IRAM[130] [1], _07799_, clk);
  dff _54788_ (\uc8051golden_1.IRAM[130] [2], _07800_, clk);
  dff _54789_ (\uc8051golden_1.IRAM[130] [3], _07801_, clk);
  dff _54790_ (\uc8051golden_1.IRAM[130] [4], _07802_, clk);
  dff _54791_ (\uc8051golden_1.IRAM[130] [5], _07803_, clk);
  dff _54792_ (\uc8051golden_1.IRAM[130] [6], _07804_, clk);
  dff _54793_ (\uc8051golden_1.IRAM[130] [7], _07805_, clk);
  dff _54794_ (\uc8051golden_1.IRAM[131] [0], _07806_, clk);
  dff _54795_ (\uc8051golden_1.IRAM[131] [1], _07807_, clk);
  dff _54796_ (\uc8051golden_1.IRAM[131] [2], _07808_, clk);
  dff _54797_ (\uc8051golden_1.IRAM[131] [3], _07809_, clk);
  dff _54798_ (\uc8051golden_1.IRAM[131] [4], _07810_, clk);
  dff _54799_ (\uc8051golden_1.IRAM[131] [5], _07811_, clk);
  dff _54800_ (\uc8051golden_1.IRAM[131] [6], _07812_, clk);
  dff _54801_ (\uc8051golden_1.IRAM[131] [7], _07813_, clk);
  dff _54802_ (\uc8051golden_1.IRAM[132] [0], _07814_, clk);
  dff _54803_ (\uc8051golden_1.IRAM[132] [1], _07815_, clk);
  dff _54804_ (\uc8051golden_1.IRAM[132] [2], _07816_, clk);
  dff _54805_ (\uc8051golden_1.IRAM[132] [3], _07817_, clk);
  dff _54806_ (\uc8051golden_1.IRAM[132] [4], _07818_, clk);
  dff _54807_ (\uc8051golden_1.IRAM[132] [5], _07819_, clk);
  dff _54808_ (\uc8051golden_1.IRAM[132] [6], _07820_, clk);
  dff _54809_ (\uc8051golden_1.IRAM[132] [7], _07821_, clk);
  dff _54810_ (\uc8051golden_1.IRAM[133] [0], _07822_, clk);
  dff _54811_ (\uc8051golden_1.IRAM[133] [1], _07823_, clk);
  dff _54812_ (\uc8051golden_1.IRAM[133] [2], _07824_, clk);
  dff _54813_ (\uc8051golden_1.IRAM[133] [3], _07825_, clk);
  dff _54814_ (\uc8051golden_1.IRAM[133] [4], _07826_, clk);
  dff _54815_ (\uc8051golden_1.IRAM[133] [5], _07827_, clk);
  dff _54816_ (\uc8051golden_1.IRAM[133] [6], _07828_, clk);
  dff _54817_ (\uc8051golden_1.IRAM[133] [7], _07829_, clk);
  dff _54818_ (\uc8051golden_1.IRAM[134] [0], _07831_, clk);
  dff _54819_ (\uc8051golden_1.IRAM[134] [1], _07832_, clk);
  dff _54820_ (\uc8051golden_1.IRAM[134] [2], _07833_, clk);
  dff _54821_ (\uc8051golden_1.IRAM[134] [3], _07834_, clk);
  dff _54822_ (\uc8051golden_1.IRAM[134] [4], _07835_, clk);
  dff _54823_ (\uc8051golden_1.IRAM[134] [5], _07836_, clk);
  dff _54824_ (\uc8051golden_1.IRAM[134] [6], _07837_, clk);
  dff _54825_ (\uc8051golden_1.IRAM[134] [7], _07838_, clk);
  dff _54826_ (\uc8051golden_1.IRAM[135] [0], _07839_, clk);
  dff _54827_ (\uc8051golden_1.IRAM[135] [1], _07840_, clk);
  dff _54828_ (\uc8051golden_1.IRAM[135] [2], _07841_, clk);
  dff _54829_ (\uc8051golden_1.IRAM[135] [3], _07842_, clk);
  dff _54830_ (\uc8051golden_1.IRAM[135] [4], _07843_, clk);
  dff _54831_ (\uc8051golden_1.IRAM[135] [5], _07844_, clk);
  dff _54832_ (\uc8051golden_1.IRAM[135] [6], _07845_, clk);
  dff _54833_ (\uc8051golden_1.IRAM[135] [7], _07846_, clk);
  dff _54834_ (\uc8051golden_1.IRAM[136] [0], _07847_, clk);
  dff _54835_ (\uc8051golden_1.IRAM[136] [1], _07848_, clk);
  dff _54836_ (\uc8051golden_1.IRAM[136] [2], _07849_, clk);
  dff _54837_ (\uc8051golden_1.IRAM[136] [3], _07850_, clk);
  dff _54838_ (\uc8051golden_1.IRAM[136] [4], _07851_, clk);
  dff _54839_ (\uc8051golden_1.IRAM[136] [5], _07852_, clk);
  dff _54840_ (\uc8051golden_1.IRAM[136] [6], _07853_, clk);
  dff _54841_ (\uc8051golden_1.IRAM[136] [7], _07854_, clk);
  dff _54842_ (\uc8051golden_1.IRAM[137] [0], _07855_, clk);
  dff _54843_ (\uc8051golden_1.IRAM[137] [1], _07856_, clk);
  dff _54844_ (\uc8051golden_1.IRAM[137] [2], _07857_, clk);
  dff _54845_ (\uc8051golden_1.IRAM[137] [3], _07858_, clk);
  dff _54846_ (\uc8051golden_1.IRAM[137] [4], _07859_, clk);
  dff _54847_ (\uc8051golden_1.IRAM[137] [5], _07860_, clk);
  dff _54848_ (\uc8051golden_1.IRAM[137] [6], _07861_, clk);
  dff _54849_ (\uc8051golden_1.IRAM[137] [7], _07862_, clk);
  dff _54850_ (\uc8051golden_1.IRAM[138] [0], _07863_, clk);
  dff _54851_ (\uc8051golden_1.IRAM[138] [1], _07865_, clk);
  dff _54852_ (\uc8051golden_1.IRAM[138] [2], _07866_, clk);
  dff _54853_ (\uc8051golden_1.IRAM[138] [3], _07867_, clk);
  dff _54854_ (\uc8051golden_1.IRAM[138] [4], _07868_, clk);
  dff _54855_ (\uc8051golden_1.IRAM[138] [5], _07869_, clk);
  dff _54856_ (\uc8051golden_1.IRAM[138] [6], _07870_, clk);
  dff _54857_ (\uc8051golden_1.IRAM[138] [7], _07871_, clk);
  dff _54858_ (\uc8051golden_1.IRAM[139] [0], _07872_, clk);
  dff _54859_ (\uc8051golden_1.IRAM[139] [1], _07873_, clk);
  dff _54860_ (\uc8051golden_1.IRAM[139] [2], _07874_, clk);
  dff _54861_ (\uc8051golden_1.IRAM[139] [3], _07875_, clk);
  dff _54862_ (\uc8051golden_1.IRAM[139] [4], _07876_, clk);
  dff _54863_ (\uc8051golden_1.IRAM[139] [5], _07877_, clk);
  dff _54864_ (\uc8051golden_1.IRAM[139] [6], _07878_, clk);
  dff _54865_ (\uc8051golden_1.IRAM[139] [7], _07879_, clk);
  dff _54866_ (\uc8051golden_1.IRAM[140] [0], _07880_, clk);
  dff _54867_ (\uc8051golden_1.IRAM[140] [1], _07881_, clk);
  dff _54868_ (\uc8051golden_1.IRAM[140] [2], _07882_, clk);
  dff _54869_ (\uc8051golden_1.IRAM[140] [3], _07883_, clk);
  dff _54870_ (\uc8051golden_1.IRAM[140] [4], _07884_, clk);
  dff _54871_ (\uc8051golden_1.IRAM[140] [5], _07885_, clk);
  dff _54872_ (\uc8051golden_1.IRAM[140] [6], _07886_, clk);
  dff _54873_ (\uc8051golden_1.IRAM[140] [7], _07887_, clk);
  dff _54874_ (\uc8051golden_1.IRAM[141] [0], _07888_, clk);
  dff _54875_ (\uc8051golden_1.IRAM[141] [1], _07889_, clk);
  dff _54876_ (\uc8051golden_1.IRAM[141] [2], _07890_, clk);
  dff _54877_ (\uc8051golden_1.IRAM[141] [3], _07891_, clk);
  dff _54878_ (\uc8051golden_1.IRAM[141] [4], _07892_, clk);
  dff _54879_ (\uc8051golden_1.IRAM[141] [5], _07893_, clk);
  dff _54880_ (\uc8051golden_1.IRAM[141] [6], _07894_, clk);
  dff _54881_ (\uc8051golden_1.IRAM[141] [7], _07895_, clk);
  dff _54882_ (\uc8051golden_1.IRAM[142] [0], _07896_, clk);
  dff _54883_ (\uc8051golden_1.IRAM[142] [1], _07897_, clk);
  dff _54884_ (\uc8051golden_1.IRAM[142] [2], _07898_, clk);
  dff _54885_ (\uc8051golden_1.IRAM[142] [3], _07900_, clk);
  dff _54886_ (\uc8051golden_1.IRAM[142] [4], _07901_, clk);
  dff _54887_ (\uc8051golden_1.IRAM[142] [5], _07902_, clk);
  dff _54888_ (\uc8051golden_1.IRAM[142] [6], _07903_, clk);
  dff _54889_ (\uc8051golden_1.IRAM[142] [7], _07904_, clk);
  dff _54890_ (\uc8051golden_1.IRAM[143] [0], _07905_, clk);
  dff _54891_ (\uc8051golden_1.IRAM[143] [1], _07906_, clk);
  dff _54892_ (\uc8051golden_1.IRAM[143] [2], _07907_, clk);
  dff _54893_ (\uc8051golden_1.IRAM[143] [3], _07908_, clk);
  dff _54894_ (\uc8051golden_1.IRAM[143] [4], _07909_, clk);
  dff _54895_ (\uc8051golden_1.IRAM[143] [5], _07910_, clk);
  dff _54896_ (\uc8051golden_1.IRAM[143] [6], _07911_, clk);
  dff _54897_ (\uc8051golden_1.IRAM[143] [7], _07912_, clk);
  dff _54898_ (\uc8051golden_1.IRAM[144] [0], _07913_, clk);
  dff _54899_ (\uc8051golden_1.IRAM[144] [1], _07914_, clk);
  dff _54900_ (\uc8051golden_1.IRAM[144] [2], _07915_, clk);
  dff _54901_ (\uc8051golden_1.IRAM[144] [3], _07916_, clk);
  dff _54902_ (\uc8051golden_1.IRAM[144] [4], _07917_, clk);
  dff _54903_ (\uc8051golden_1.IRAM[144] [5], _07918_, clk);
  dff _54904_ (\uc8051golden_1.IRAM[144] [6], _07919_, clk);
  dff _54905_ (\uc8051golden_1.IRAM[144] [7], _07920_, clk);
  dff _54906_ (\uc8051golden_1.IRAM[145] [0], _07921_, clk);
  dff _54907_ (\uc8051golden_1.IRAM[145] [1], _07922_, clk);
  dff _54908_ (\uc8051golden_1.IRAM[145] [2], _07923_, clk);
  dff _54909_ (\uc8051golden_1.IRAM[145] [3], _07924_, clk);
  dff _54910_ (\uc8051golden_1.IRAM[145] [4], _07925_, clk);
  dff _54911_ (\uc8051golden_1.IRAM[145] [5], _07926_, clk);
  dff _54912_ (\uc8051golden_1.IRAM[145] [6], _07927_, clk);
  dff _54913_ (\uc8051golden_1.IRAM[145] [7], _07928_, clk);
  dff _54914_ (\uc8051golden_1.IRAM[146] [0], _07929_, clk);
  dff _54915_ (\uc8051golden_1.IRAM[146] [1], _07930_, clk);
  dff _54916_ (\uc8051golden_1.IRAM[146] [2], _07931_, clk);
  dff _54917_ (\uc8051golden_1.IRAM[146] [3], _07932_, clk);
  dff _54918_ (\uc8051golden_1.IRAM[146] [4], _07934_, clk);
  dff _54919_ (\uc8051golden_1.IRAM[146] [5], _07935_, clk);
  dff _54920_ (\uc8051golden_1.IRAM[146] [6], _07936_, clk);
  dff _54921_ (\uc8051golden_1.IRAM[146] [7], _07937_, clk);
  dff _54922_ (\uc8051golden_1.IRAM[147] [0], _07938_, clk);
  dff _54923_ (\uc8051golden_1.IRAM[147] [1], _07939_, clk);
  dff _54924_ (\uc8051golden_1.IRAM[147] [2], _07940_, clk);
  dff _54925_ (\uc8051golden_1.IRAM[147] [3], _07941_, clk);
  dff _54926_ (\uc8051golden_1.IRAM[147] [4], _07942_, clk);
  dff _54927_ (\uc8051golden_1.IRAM[147] [5], _07943_, clk);
  dff _54928_ (\uc8051golden_1.IRAM[147] [6], _07944_, clk);
  dff _54929_ (\uc8051golden_1.IRAM[147] [7], _07945_, clk);
  dff _54930_ (\uc8051golden_1.IRAM[148] [0], _07946_, clk);
  dff _54931_ (\uc8051golden_1.IRAM[148] [1], _07947_, clk);
  dff _54932_ (\uc8051golden_1.IRAM[148] [2], _07948_, clk);
  dff _54933_ (\uc8051golden_1.IRAM[148] [3], _07949_, clk);
  dff _54934_ (\uc8051golden_1.IRAM[148] [4], _07950_, clk);
  dff _54935_ (\uc8051golden_1.IRAM[148] [5], _07951_, clk);
  dff _54936_ (\uc8051golden_1.IRAM[148] [6], _07952_, clk);
  dff _54937_ (\uc8051golden_1.IRAM[148] [7], _07953_, clk);
  dff _54938_ (\uc8051golden_1.IRAM[149] [0], _07954_, clk);
  dff _54939_ (\uc8051golden_1.IRAM[149] [1], _07955_, clk);
  dff _54940_ (\uc8051golden_1.IRAM[149] [2], _07956_, clk);
  dff _54941_ (\uc8051golden_1.IRAM[149] [3], _07957_, clk);
  dff _54942_ (\uc8051golden_1.IRAM[149] [4], _07958_, clk);
  dff _54943_ (\uc8051golden_1.IRAM[149] [5], _07959_, clk);
  dff _54944_ (\uc8051golden_1.IRAM[149] [6], _07960_, clk);
  dff _54945_ (\uc8051golden_1.IRAM[149] [7], _07961_, clk);
  dff _54946_ (\uc8051golden_1.IRAM[150] [0], _07962_, clk);
  dff _54947_ (\uc8051golden_1.IRAM[150] [1], _07963_, clk);
  dff _54948_ (\uc8051golden_1.IRAM[150] [2], _07964_, clk);
  dff _54949_ (\uc8051golden_1.IRAM[150] [3], _07965_, clk);
  dff _54950_ (\uc8051golden_1.IRAM[150] [4], _07966_, clk);
  dff _54951_ (\uc8051golden_1.IRAM[150] [5], _07968_, clk);
  dff _54952_ (\uc8051golden_1.IRAM[150] [6], _07969_, clk);
  dff _54953_ (\uc8051golden_1.IRAM[150] [7], _07970_, clk);
  dff _54954_ (\uc8051golden_1.IRAM[151] [0], _07971_, clk);
  dff _54955_ (\uc8051golden_1.IRAM[151] [1], _07972_, clk);
  dff _54956_ (\uc8051golden_1.IRAM[151] [2], _07973_, clk);
  dff _54957_ (\uc8051golden_1.IRAM[151] [3], _07974_, clk);
  dff _54958_ (\uc8051golden_1.IRAM[151] [4], _07975_, clk);
  dff _54959_ (\uc8051golden_1.IRAM[151] [5], _07976_, clk);
  dff _54960_ (\uc8051golden_1.IRAM[151] [6], _07977_, clk);
  dff _54961_ (\uc8051golden_1.IRAM[151] [7], _07978_, clk);
  dff _54962_ (\uc8051golden_1.IRAM[152] [0], _07979_, clk);
  dff _54963_ (\uc8051golden_1.IRAM[152] [1], _07980_, clk);
  dff _54964_ (\uc8051golden_1.IRAM[152] [2], _07981_, clk);
  dff _54965_ (\uc8051golden_1.IRAM[152] [3], _07982_, clk);
  dff _54966_ (\uc8051golden_1.IRAM[152] [4], _07983_, clk);
  dff _54967_ (\uc8051golden_1.IRAM[152] [5], _07984_, clk);
  dff _54968_ (\uc8051golden_1.IRAM[152] [6], _07985_, clk);
  dff _54969_ (\uc8051golden_1.IRAM[152] [7], _07986_, clk);
  dff _54970_ (\uc8051golden_1.IRAM[153] [0], _07987_, clk);
  dff _54971_ (\uc8051golden_1.IRAM[153] [1], _07988_, clk);
  dff _54972_ (\uc8051golden_1.IRAM[153] [2], _07989_, clk);
  dff _54973_ (\uc8051golden_1.IRAM[153] [3], _07990_, clk);
  dff _54974_ (\uc8051golden_1.IRAM[153] [4], _07991_, clk);
  dff _54975_ (\uc8051golden_1.IRAM[153] [5], _07992_, clk);
  dff _54976_ (\uc8051golden_1.IRAM[153] [6], _07993_, clk);
  dff _54977_ (\uc8051golden_1.IRAM[153] [7], _07994_, clk);
  dff _54978_ (\uc8051golden_1.IRAM[154] [0], _07995_, clk);
  dff _54979_ (\uc8051golden_1.IRAM[154] [1], _07996_, clk);
  dff _54980_ (\uc8051golden_1.IRAM[154] [2], _07997_, clk);
  dff _54981_ (\uc8051golden_1.IRAM[154] [3], _07998_, clk);
  dff _54982_ (\uc8051golden_1.IRAM[154] [4], _07999_, clk);
  dff _54983_ (\uc8051golden_1.IRAM[154] [5], _08000_, clk);
  dff _54984_ (\uc8051golden_1.IRAM[154] [6], _08002_, clk);
  dff _54985_ (\uc8051golden_1.IRAM[154] [7], _08003_, clk);
  dff _54986_ (\uc8051golden_1.IRAM[155] [0], _08004_, clk);
  dff _54987_ (\uc8051golden_1.IRAM[155] [1], _08005_, clk);
  dff _54988_ (\uc8051golden_1.IRAM[155] [2], _08006_, clk);
  dff _54989_ (\uc8051golden_1.IRAM[155] [3], _08007_, clk);
  dff _54990_ (\uc8051golden_1.IRAM[155] [4], _08008_, clk);
  dff _54991_ (\uc8051golden_1.IRAM[155] [5], _08009_, clk);
  dff _54992_ (\uc8051golden_1.IRAM[155] [6], _08010_, clk);
  dff _54993_ (\uc8051golden_1.IRAM[155] [7], _08011_, clk);
  dff _54994_ (\uc8051golden_1.IRAM[156] [0], _08012_, clk);
  dff _54995_ (\uc8051golden_1.IRAM[156] [1], _08013_, clk);
  dff _54996_ (\uc8051golden_1.IRAM[156] [2], _08014_, clk);
  dff _54997_ (\uc8051golden_1.IRAM[156] [3], _08015_, clk);
  dff _54998_ (\uc8051golden_1.IRAM[156] [4], _08016_, clk);
  dff _54999_ (\uc8051golden_1.IRAM[156] [5], _08017_, clk);
  dff _55000_ (\uc8051golden_1.IRAM[156] [6], _08018_, clk);
  dff _55001_ (\uc8051golden_1.IRAM[156] [7], _08019_, clk);
  dff _55002_ (\uc8051golden_1.IRAM[157] [0], _08020_, clk);
  dff _55003_ (\uc8051golden_1.IRAM[157] [1], _08021_, clk);
  dff _55004_ (\uc8051golden_1.IRAM[157] [2], _08022_, clk);
  dff _55005_ (\uc8051golden_1.IRAM[157] [3], _08023_, clk);
  dff _55006_ (\uc8051golden_1.IRAM[157] [4], _08024_, clk);
  dff _55007_ (\uc8051golden_1.IRAM[157] [5], _08025_, clk);
  dff _55008_ (\uc8051golden_1.IRAM[157] [6], _08026_, clk);
  dff _55009_ (\uc8051golden_1.IRAM[157] [7], _08027_, clk);
  dff _55010_ (\uc8051golden_1.IRAM[158] [0], _08028_, clk);
  dff _55011_ (\uc8051golden_1.IRAM[158] [1], _08029_, clk);
  dff _55012_ (\uc8051golden_1.IRAM[158] [2], _08030_, clk);
  dff _55013_ (\uc8051golden_1.IRAM[158] [3], _08031_, clk);
  dff _55014_ (\uc8051golden_1.IRAM[158] [4], _08032_, clk);
  dff _55015_ (\uc8051golden_1.IRAM[158] [5], _08033_, clk);
  dff _55016_ (\uc8051golden_1.IRAM[158] [6], _08034_, clk);
  dff _55017_ (\uc8051golden_1.IRAM[158] [7], _08035_, clk);
  dff _55018_ (\uc8051golden_1.IRAM[159] [0], _08037_, clk);
  dff _55019_ (\uc8051golden_1.IRAM[159] [1], _08038_, clk);
  dff _55020_ (\uc8051golden_1.IRAM[159] [2], _08039_, clk);
  dff _55021_ (\uc8051golden_1.IRAM[159] [3], _08040_, clk);
  dff _55022_ (\uc8051golden_1.IRAM[159] [4], _08041_, clk);
  dff _55023_ (\uc8051golden_1.IRAM[159] [5], _08042_, clk);
  dff _55024_ (\uc8051golden_1.IRAM[159] [6], _08043_, clk);
  dff _55025_ (\uc8051golden_1.IRAM[159] [7], _08044_, clk);
  dff _55026_ (\uc8051golden_1.IRAM[160] [0], _08045_, clk);
  dff _55027_ (\uc8051golden_1.IRAM[160] [1], _08046_, clk);
  dff _55028_ (\uc8051golden_1.IRAM[160] [2], _08047_, clk);
  dff _55029_ (\uc8051golden_1.IRAM[160] [3], _08048_, clk);
  dff _55030_ (\uc8051golden_1.IRAM[160] [4], _08049_, clk);
  dff _55031_ (\uc8051golden_1.IRAM[160] [5], _08050_, clk);
  dff _55032_ (\uc8051golden_1.IRAM[160] [6], _08051_, clk);
  dff _55033_ (\uc8051golden_1.IRAM[160] [7], _08052_, clk);
  dff _55034_ (\uc8051golden_1.IRAM[161] [0], _08053_, clk);
  dff _55035_ (\uc8051golden_1.IRAM[161] [1], _08054_, clk);
  dff _55036_ (\uc8051golden_1.IRAM[161] [2], _08055_, clk);
  dff _55037_ (\uc8051golden_1.IRAM[161] [3], _08056_, clk);
  dff _55038_ (\uc8051golden_1.IRAM[161] [4], _08057_, clk);
  dff _55039_ (\uc8051golden_1.IRAM[161] [5], _08058_, clk);
  dff _55040_ (\uc8051golden_1.IRAM[161] [6], _08059_, clk);
  dff _55041_ (\uc8051golden_1.IRAM[161] [7], _08060_, clk);
  dff _55042_ (\uc8051golden_1.IRAM[162] [0], _08061_, clk);
  dff _55043_ (\uc8051golden_1.IRAM[162] [1], _08062_, clk);
  dff _55044_ (\uc8051golden_1.IRAM[162] [2], _08063_, clk);
  dff _55045_ (\uc8051golden_1.IRAM[162] [3], _08064_, clk);
  dff _55046_ (\uc8051golden_1.IRAM[162] [4], _08065_, clk);
  dff _55047_ (\uc8051golden_1.IRAM[162] [5], _08066_, clk);
  dff _55048_ (\uc8051golden_1.IRAM[162] [6], _08067_, clk);
  dff _55049_ (\uc8051golden_1.IRAM[162] [7], _08068_, clk);
  dff _55050_ (\uc8051golden_1.IRAM[163] [0], _08069_, clk);
  dff _55051_ (\uc8051golden_1.IRAM[163] [1], _08071_, clk);
  dff _55052_ (\uc8051golden_1.IRAM[163] [2], _08072_, clk);
  dff _55053_ (\uc8051golden_1.IRAM[163] [3], _08073_, clk);
  dff _55054_ (\uc8051golden_1.IRAM[163] [4], _08074_, clk);
  dff _55055_ (\uc8051golden_1.IRAM[163] [5], _08075_, clk);
  dff _55056_ (\uc8051golden_1.IRAM[163] [6], _08076_, clk);
  dff _55057_ (\uc8051golden_1.IRAM[163] [7], _08077_, clk);
  dff _55058_ (\uc8051golden_1.IRAM[164] [0], _08078_, clk);
  dff _55059_ (\uc8051golden_1.IRAM[164] [1], _08079_, clk);
  dff _55060_ (\uc8051golden_1.IRAM[164] [2], _08080_, clk);
  dff _55061_ (\uc8051golden_1.IRAM[164] [3], _08081_, clk);
  dff _55062_ (\uc8051golden_1.IRAM[164] [4], _08082_, clk);
  dff _55063_ (\uc8051golden_1.IRAM[164] [5], _08083_, clk);
  dff _55064_ (\uc8051golden_1.IRAM[164] [6], _08084_, clk);
  dff _55065_ (\uc8051golden_1.IRAM[164] [7], _08085_, clk);
  dff _55066_ (\uc8051golden_1.IRAM[165] [0], _08086_, clk);
  dff _55067_ (\uc8051golden_1.IRAM[165] [1], _08087_, clk);
  dff _55068_ (\uc8051golden_1.IRAM[165] [2], _08088_, clk);
  dff _55069_ (\uc8051golden_1.IRAM[165] [3], _08089_, clk);
  dff _55070_ (\uc8051golden_1.IRAM[165] [4], _08090_, clk);
  dff _55071_ (\uc8051golden_1.IRAM[165] [5], _08091_, clk);
  dff _55072_ (\uc8051golden_1.IRAM[165] [6], _08092_, clk);
  dff _55073_ (\uc8051golden_1.IRAM[165] [7], _08093_, clk);
  dff _55074_ (\uc8051golden_1.IRAM[166] [0], _08094_, clk);
  dff _55075_ (\uc8051golden_1.IRAM[166] [1], _08095_, clk);
  dff _55076_ (\uc8051golden_1.IRAM[166] [2], _08096_, clk);
  dff _55077_ (\uc8051golden_1.IRAM[166] [3], _08097_, clk);
  dff _55078_ (\uc8051golden_1.IRAM[166] [4], _08098_, clk);
  dff _55079_ (\uc8051golden_1.IRAM[166] [5], _08099_, clk);
  dff _55080_ (\uc8051golden_1.IRAM[166] [6], _08100_, clk);
  dff _55081_ (\uc8051golden_1.IRAM[166] [7], _08101_, clk);
  dff _55082_ (\uc8051golden_1.IRAM[167] [0], _08102_, clk);
  dff _55083_ (\uc8051golden_1.IRAM[167] [1], _08103_, clk);
  dff _55084_ (\uc8051golden_1.IRAM[167] [2], _08105_, clk);
  dff _55085_ (\uc8051golden_1.IRAM[167] [3], _08106_, clk);
  dff _55086_ (\uc8051golden_1.IRAM[167] [4], _08107_, clk);
  dff _55087_ (\uc8051golden_1.IRAM[167] [5], _08108_, clk);
  dff _55088_ (\uc8051golden_1.IRAM[167] [6], _08109_, clk);
  dff _55089_ (\uc8051golden_1.IRAM[167] [7], _08110_, clk);
  dff _55090_ (\uc8051golden_1.IRAM[168] [0], _08111_, clk);
  dff _55091_ (\uc8051golden_1.IRAM[168] [1], _08112_, clk);
  dff _55092_ (\uc8051golden_1.IRAM[168] [2], _08113_, clk);
  dff _55093_ (\uc8051golden_1.IRAM[168] [3], _08114_, clk);
  dff _55094_ (\uc8051golden_1.IRAM[168] [4], _08115_, clk);
  dff _55095_ (\uc8051golden_1.IRAM[168] [5], _08116_, clk);
  dff _55096_ (\uc8051golden_1.IRAM[168] [6], _08117_, clk);
  dff _55097_ (\uc8051golden_1.IRAM[168] [7], _08118_, clk);
  dff _55098_ (\uc8051golden_1.IRAM[169] [0], _08119_, clk);
  dff _55099_ (\uc8051golden_1.IRAM[169] [1], _08120_, clk);
  dff _55100_ (\uc8051golden_1.IRAM[169] [2], _08121_, clk);
  dff _55101_ (\uc8051golden_1.IRAM[169] [3], _08122_, clk);
  dff _55102_ (\uc8051golden_1.IRAM[169] [4], _08123_, clk);
  dff _55103_ (\uc8051golden_1.IRAM[169] [5], _08124_, clk);
  dff _55104_ (\uc8051golden_1.IRAM[169] [6], _08125_, clk);
  dff _55105_ (\uc8051golden_1.IRAM[169] [7], _08126_, clk);
  dff _55106_ (\uc8051golden_1.IRAM[170] [0], _08127_, clk);
  dff _55107_ (\uc8051golden_1.IRAM[170] [1], _08128_, clk);
  dff _55108_ (\uc8051golden_1.IRAM[170] [2], _08129_, clk);
  dff _55109_ (\uc8051golden_1.IRAM[170] [3], _08130_, clk);
  dff _55110_ (\uc8051golden_1.IRAM[170] [4], _08131_, clk);
  dff _55111_ (\uc8051golden_1.IRAM[170] [5], _08132_, clk);
  dff _55112_ (\uc8051golden_1.IRAM[170] [6], _08133_, clk);
  dff _55113_ (\uc8051golden_1.IRAM[170] [7], _08134_, clk);
  dff _55114_ (\uc8051golden_1.IRAM[171] [0], _08135_, clk);
  dff _55115_ (\uc8051golden_1.IRAM[171] [1], _08136_, clk);
  dff _55116_ (\uc8051golden_1.IRAM[171] [2], _08137_, clk);
  dff _55117_ (\uc8051golden_1.IRAM[171] [3], _08139_, clk);
  dff _55118_ (\uc8051golden_1.IRAM[171] [4], _08140_, clk);
  dff _55119_ (\uc8051golden_1.IRAM[171] [5], _08141_, clk);
  dff _55120_ (\uc8051golden_1.IRAM[171] [6], _08142_, clk);
  dff _55121_ (\uc8051golden_1.IRAM[171] [7], _08143_, clk);
  dff _55122_ (\uc8051golden_1.IRAM[172] [0], _08144_, clk);
  dff _55123_ (\uc8051golden_1.IRAM[172] [1], _08145_, clk);
  dff _55124_ (\uc8051golden_1.IRAM[172] [2], _08146_, clk);
  dff _55125_ (\uc8051golden_1.IRAM[172] [3], _08147_, clk);
  dff _55126_ (\uc8051golden_1.IRAM[172] [4], _08148_, clk);
  dff _55127_ (\uc8051golden_1.IRAM[172] [5], _08149_, clk);
  dff _55128_ (\uc8051golden_1.IRAM[172] [6], _08150_, clk);
  dff _55129_ (\uc8051golden_1.IRAM[172] [7], _08151_, clk);
  dff _55130_ (\uc8051golden_1.IRAM[173] [0], _08152_, clk);
  dff _55131_ (\uc8051golden_1.IRAM[173] [1], _08153_, clk);
  dff _55132_ (\uc8051golden_1.IRAM[173] [2], _08154_, clk);
  dff _55133_ (\uc8051golden_1.IRAM[173] [3], _08155_, clk);
  dff _55134_ (\uc8051golden_1.IRAM[173] [4], _08156_, clk);
  dff _55135_ (\uc8051golden_1.IRAM[173] [5], _08157_, clk);
  dff _55136_ (\uc8051golden_1.IRAM[173] [6], _08158_, clk);
  dff _55137_ (\uc8051golden_1.IRAM[173] [7], _08159_, clk);
  dff _55138_ (\uc8051golden_1.IRAM[174] [0], _08160_, clk);
  dff _55139_ (\uc8051golden_1.IRAM[174] [1], _08161_, clk);
  dff _55140_ (\uc8051golden_1.IRAM[174] [2], _08162_, clk);
  dff _55141_ (\uc8051golden_1.IRAM[174] [3], _08163_, clk);
  dff _55142_ (\uc8051golden_1.IRAM[174] [4], _08164_, clk);
  dff _55143_ (\uc8051golden_1.IRAM[174] [5], _08165_, clk);
  dff _55144_ (\uc8051golden_1.IRAM[174] [6], _08166_, clk);
  dff _55145_ (\uc8051golden_1.IRAM[174] [7], _08167_, clk);
  dff _55146_ (\uc8051golden_1.IRAM[175] [0], _08168_, clk);
  dff _55147_ (\uc8051golden_1.IRAM[175] [1], _08169_, clk);
  dff _55148_ (\uc8051golden_1.IRAM[175] [2], _08170_, clk);
  dff _55149_ (\uc8051golden_1.IRAM[175] [3], _08171_, clk);
  dff _55150_ (\uc8051golden_1.IRAM[175] [4], _08172_, clk);
  dff _55151_ (\uc8051golden_1.IRAM[175] [5], _08174_, clk);
  dff _55152_ (\uc8051golden_1.IRAM[175] [6], _08175_, clk);
  dff _55153_ (\uc8051golden_1.IRAM[175] [7], _08176_, clk);
  dff _55154_ (\uc8051golden_1.IRAM[176] [0], _08177_, clk);
  dff _55155_ (\uc8051golden_1.IRAM[176] [1], _08178_, clk);
  dff _55156_ (\uc8051golden_1.IRAM[176] [2], _08179_, clk);
  dff _55157_ (\uc8051golden_1.IRAM[176] [3], _08180_, clk);
  dff _55158_ (\uc8051golden_1.IRAM[176] [4], _08181_, clk);
  dff _55159_ (\uc8051golden_1.IRAM[176] [5], _08182_, clk);
  dff _55160_ (\uc8051golden_1.IRAM[176] [6], _08183_, clk);
  dff _55161_ (\uc8051golden_1.IRAM[176] [7], _08184_, clk);
  dff _55162_ (\uc8051golden_1.IRAM[177] [0], _08185_, clk);
  dff _55163_ (\uc8051golden_1.IRAM[177] [1], _08186_, clk);
  dff _55164_ (\uc8051golden_1.IRAM[177] [2], _08187_, clk);
  dff _55165_ (\uc8051golden_1.IRAM[177] [3], _08188_, clk);
  dff _55166_ (\uc8051golden_1.IRAM[177] [4], _08189_, clk);
  dff _55167_ (\uc8051golden_1.IRAM[177] [5], _08190_, clk);
  dff _55168_ (\uc8051golden_1.IRAM[177] [6], _08191_, clk);
  dff _55169_ (\uc8051golden_1.IRAM[177] [7], _08192_, clk);
  dff _55170_ (\uc8051golden_1.IRAM[178] [0], _08193_, clk);
  dff _55171_ (\uc8051golden_1.IRAM[178] [1], _08194_, clk);
  dff _55172_ (\uc8051golden_1.IRAM[178] [2], _08195_, clk);
  dff _55173_ (\uc8051golden_1.IRAM[178] [3], _08196_, clk);
  dff _55174_ (\uc8051golden_1.IRAM[178] [4], _08197_, clk);
  dff _55175_ (\uc8051golden_1.IRAM[178] [5], _08198_, clk);
  dff _55176_ (\uc8051golden_1.IRAM[178] [6], _08199_, clk);
  dff _55177_ (\uc8051golden_1.IRAM[178] [7], _08200_, clk);
  dff _55178_ (\uc8051golden_1.IRAM[179] [0], _08201_, clk);
  dff _55179_ (\uc8051golden_1.IRAM[179] [1], _08202_, clk);
  dff _55180_ (\uc8051golden_1.IRAM[179] [2], _08203_, clk);
  dff _55181_ (\uc8051golden_1.IRAM[179] [3], _08204_, clk);
  dff _55182_ (\uc8051golden_1.IRAM[179] [4], _08205_, clk);
  dff _55183_ (\uc8051golden_1.IRAM[179] [5], _08206_, clk);
  dff _55184_ (\uc8051golden_1.IRAM[179] [6], _08208_, clk);
  dff _55185_ (\uc8051golden_1.IRAM[179] [7], _08209_, clk);
  dff _55186_ (\uc8051golden_1.IRAM[180] [0], _08210_, clk);
  dff _55187_ (\uc8051golden_1.IRAM[180] [1], _08211_, clk);
  dff _55188_ (\uc8051golden_1.IRAM[180] [2], _08212_, clk);
  dff _55189_ (\uc8051golden_1.IRAM[180] [3], _08213_, clk);
  dff _55190_ (\uc8051golden_1.IRAM[180] [4], _08214_, clk);
  dff _55191_ (\uc8051golden_1.IRAM[180] [5], _08215_, clk);
  dff _55192_ (\uc8051golden_1.IRAM[180] [6], _08216_, clk);
  dff _55193_ (\uc8051golden_1.IRAM[180] [7], _08217_, clk);
  dff _55194_ (\uc8051golden_1.IRAM[181] [0], _08218_, clk);
  dff _55195_ (\uc8051golden_1.IRAM[181] [1], _08219_, clk);
  dff _55196_ (\uc8051golden_1.IRAM[181] [2], _08220_, clk);
  dff _55197_ (\uc8051golden_1.IRAM[181] [3], _08221_, clk);
  dff _55198_ (\uc8051golden_1.IRAM[181] [4], _08222_, clk);
  dff _55199_ (\uc8051golden_1.IRAM[181] [5], _08223_, clk);
  dff _55200_ (\uc8051golden_1.IRAM[181] [6], _08224_, clk);
  dff _55201_ (\uc8051golden_1.IRAM[181] [7], _08225_, clk);
  dff _55202_ (\uc8051golden_1.IRAM[182] [0], _08226_, clk);
  dff _55203_ (\uc8051golden_1.IRAM[182] [1], _08227_, clk);
  dff _55204_ (\uc8051golden_1.IRAM[182] [2], _08228_, clk);
  dff _55205_ (\uc8051golden_1.IRAM[182] [3], _08229_, clk);
  dff _55206_ (\uc8051golden_1.IRAM[182] [4], _08230_, clk);
  dff _55207_ (\uc8051golden_1.IRAM[182] [5], _08231_, clk);
  dff _55208_ (\uc8051golden_1.IRAM[182] [6], _08232_, clk);
  dff _55209_ (\uc8051golden_1.IRAM[182] [7], _08233_, clk);
  dff _55210_ (\uc8051golden_1.IRAM[183] [0], _08234_, clk);
  dff _55211_ (\uc8051golden_1.IRAM[183] [1], _08235_, clk);
  dff _55212_ (\uc8051golden_1.IRAM[183] [2], _08236_, clk);
  dff _55213_ (\uc8051golden_1.IRAM[183] [3], _08237_, clk);
  dff _55214_ (\uc8051golden_1.IRAM[183] [4], _08238_, clk);
  dff _55215_ (\uc8051golden_1.IRAM[183] [5], _08239_, clk);
  dff _55216_ (\uc8051golden_1.IRAM[183] [6], _08240_, clk);
  dff _55217_ (\uc8051golden_1.IRAM[183] [7], _08242_, clk);
  dff _55218_ (\uc8051golden_1.IRAM[184] [0], _08243_, clk);
  dff _55219_ (\uc8051golden_1.IRAM[184] [1], _08244_, clk);
  dff _55220_ (\uc8051golden_1.IRAM[184] [2], _08245_, clk);
  dff _55221_ (\uc8051golden_1.IRAM[184] [3], _08246_, clk);
  dff _55222_ (\uc8051golden_1.IRAM[184] [4], _08247_, clk);
  dff _55223_ (\uc8051golden_1.IRAM[184] [5], _08248_, clk);
  dff _55224_ (\uc8051golden_1.IRAM[184] [6], _08249_, clk);
  dff _55225_ (\uc8051golden_1.IRAM[184] [7], _08250_, clk);
  dff _55226_ (\uc8051golden_1.IRAM[185] [0], _08251_, clk);
  dff _55227_ (\uc8051golden_1.IRAM[185] [1], _08252_, clk);
  dff _55228_ (\uc8051golden_1.IRAM[185] [2], _08253_, clk);
  dff _55229_ (\uc8051golden_1.IRAM[185] [3], _08254_, clk);
  dff _55230_ (\uc8051golden_1.IRAM[185] [4], _08255_, clk);
  dff _55231_ (\uc8051golden_1.IRAM[185] [5], _08256_, clk);
  dff _55232_ (\uc8051golden_1.IRAM[185] [6], _08257_, clk);
  dff _55233_ (\uc8051golden_1.IRAM[185] [7], _08258_, clk);
  dff _55234_ (\uc8051golden_1.IRAM[186] [0], _08259_, clk);
  dff _55235_ (\uc8051golden_1.IRAM[186] [1], _08260_, clk);
  dff _55236_ (\uc8051golden_1.IRAM[186] [2], _08261_, clk);
  dff _55237_ (\uc8051golden_1.IRAM[186] [3], _08262_, clk);
  dff _55238_ (\uc8051golden_1.IRAM[186] [4], _08263_, clk);
  dff _55239_ (\uc8051golden_1.IRAM[186] [5], _08264_, clk);
  dff _55240_ (\uc8051golden_1.IRAM[186] [6], _08265_, clk);
  dff _55241_ (\uc8051golden_1.IRAM[186] [7], _08266_, clk);
  dff _55242_ (\uc8051golden_1.IRAM[187] [0], _08267_, clk);
  dff _55243_ (\uc8051golden_1.IRAM[187] [1], _08268_, clk);
  dff _55244_ (\uc8051golden_1.IRAM[187] [2], _08269_, clk);
  dff _55245_ (\uc8051golden_1.IRAM[187] [3], _08270_, clk);
  dff _55246_ (\uc8051golden_1.IRAM[187] [4], _08271_, clk);
  dff _55247_ (\uc8051golden_1.IRAM[187] [5], _08272_, clk);
  dff _55248_ (\uc8051golden_1.IRAM[187] [6], _08273_, clk);
  dff _55249_ (\uc8051golden_1.IRAM[187] [7], _08274_, clk);
  dff _55250_ (\uc8051golden_1.IRAM[188] [0], _08276_, clk);
  dff _55251_ (\uc8051golden_1.IRAM[188] [1], _08277_, clk);
  dff _55252_ (\uc8051golden_1.IRAM[188] [2], _08278_, clk);
  dff _55253_ (\uc8051golden_1.IRAM[188] [3], _08279_, clk);
  dff _55254_ (\uc8051golden_1.IRAM[188] [4], _08280_, clk);
  dff _55255_ (\uc8051golden_1.IRAM[188] [5], _08281_, clk);
  dff _55256_ (\uc8051golden_1.IRAM[188] [6], _08282_, clk);
  dff _55257_ (\uc8051golden_1.IRAM[188] [7], _08283_, clk);
  dff _55258_ (\uc8051golden_1.IRAM[189] [0], _08284_, clk);
  dff _55259_ (\uc8051golden_1.IRAM[189] [1], _08285_, clk);
  dff _55260_ (\uc8051golden_1.IRAM[189] [2], _08286_, clk);
  dff _55261_ (\uc8051golden_1.IRAM[189] [3], _08287_, clk);
  dff _55262_ (\uc8051golden_1.IRAM[189] [4], _08288_, clk);
  dff _55263_ (\uc8051golden_1.IRAM[189] [5], _08289_, clk);
  dff _55264_ (\uc8051golden_1.IRAM[189] [6], _08290_, clk);
  dff _55265_ (\uc8051golden_1.IRAM[189] [7], _08291_, clk);
  dff _55266_ (\uc8051golden_1.IRAM[190] [0], _08292_, clk);
  dff _55267_ (\uc8051golden_1.IRAM[190] [1], _08293_, clk);
  dff _55268_ (\uc8051golden_1.IRAM[190] [2], _08294_, clk);
  dff _55269_ (\uc8051golden_1.IRAM[190] [3], _08295_, clk);
  dff _55270_ (\uc8051golden_1.IRAM[190] [4], _08296_, clk);
  dff _55271_ (\uc8051golden_1.IRAM[190] [5], _08297_, clk);
  dff _55272_ (\uc8051golden_1.IRAM[190] [6], _08298_, clk);
  dff _55273_ (\uc8051golden_1.IRAM[190] [7], _08299_, clk);
  dff _55274_ (\uc8051golden_1.IRAM[191] [0], _08300_, clk);
  dff _55275_ (\uc8051golden_1.IRAM[191] [1], _08301_, clk);
  dff _55276_ (\uc8051golden_1.IRAM[191] [2], _08302_, clk);
  dff _55277_ (\uc8051golden_1.IRAM[191] [3], _08303_, clk);
  dff _55278_ (\uc8051golden_1.IRAM[191] [4], _08304_, clk);
  dff _55279_ (\uc8051golden_1.IRAM[191] [5], _08305_, clk);
  dff _55280_ (\uc8051golden_1.IRAM[191] [6], _08306_, clk);
  dff _55281_ (\uc8051golden_1.IRAM[191] [7], _08307_, clk);
  dff _55282_ (\uc8051golden_1.IRAM[192] [0], _08308_, clk);
  dff _55283_ (\uc8051golden_1.IRAM[192] [1], _08310_, clk);
  dff _55284_ (\uc8051golden_1.IRAM[192] [2], _08311_, clk);
  dff _55285_ (\uc8051golden_1.IRAM[192] [3], _08312_, clk);
  dff _55286_ (\uc8051golden_1.IRAM[192] [4], _08313_, clk);
  dff _55287_ (\uc8051golden_1.IRAM[192] [5], _08314_, clk);
  dff _55288_ (\uc8051golden_1.IRAM[192] [6], _08315_, clk);
  dff _55289_ (\uc8051golden_1.IRAM[192] [7], _08316_, clk);
  dff _55290_ (\uc8051golden_1.IRAM[193] [0], _08317_, clk);
  dff _55291_ (\uc8051golden_1.IRAM[193] [1], _08318_, clk);
  dff _55292_ (\uc8051golden_1.IRAM[193] [2], _08319_, clk);
  dff _55293_ (\uc8051golden_1.IRAM[193] [3], _08320_, clk);
  dff _55294_ (\uc8051golden_1.IRAM[193] [4], _08321_, clk);
  dff _55295_ (\uc8051golden_1.IRAM[193] [5], _08322_, clk);
  dff _55296_ (\uc8051golden_1.IRAM[193] [6], _08323_, clk);
  dff _55297_ (\uc8051golden_1.IRAM[193] [7], _08324_, clk);
  dff _55298_ (\uc8051golden_1.IRAM[194] [0], _08325_, clk);
  dff _55299_ (\uc8051golden_1.IRAM[194] [1], _08326_, clk);
  dff _55300_ (\uc8051golden_1.IRAM[194] [2], _08327_, clk);
  dff _55301_ (\uc8051golden_1.IRAM[194] [3], _08328_, clk);
  dff _55302_ (\uc8051golden_1.IRAM[194] [4], _08329_, clk);
  dff _55303_ (\uc8051golden_1.IRAM[194] [5], _08330_, clk);
  dff _55304_ (\uc8051golden_1.IRAM[194] [6], _08331_, clk);
  dff _55305_ (\uc8051golden_1.IRAM[194] [7], _08332_, clk);
  dff _55306_ (\uc8051golden_1.IRAM[195] [0], _08333_, clk);
  dff _55307_ (\uc8051golden_1.IRAM[195] [1], _08334_, clk);
  dff _55308_ (\uc8051golden_1.IRAM[195] [2], _08335_, clk);
  dff _55309_ (\uc8051golden_1.IRAM[195] [3], _08336_, clk);
  dff _55310_ (\uc8051golden_1.IRAM[195] [4], _08337_, clk);
  dff _55311_ (\uc8051golden_1.IRAM[195] [5], _08338_, clk);
  dff _55312_ (\uc8051golden_1.IRAM[195] [6], _08339_, clk);
  dff _55313_ (\uc8051golden_1.IRAM[195] [7], _08340_, clk);
  dff _55314_ (\uc8051golden_1.IRAM[196] [0], _08341_, clk);
  dff _55315_ (\uc8051golden_1.IRAM[196] [1], _08342_, clk);
  dff _55316_ (\uc8051golden_1.IRAM[196] [2], _08344_, clk);
  dff _55317_ (\uc8051golden_1.IRAM[196] [3], _08345_, clk);
  dff _55318_ (\uc8051golden_1.IRAM[196] [4], _08346_, clk);
  dff _55319_ (\uc8051golden_1.IRAM[196] [5], _08347_, clk);
  dff _55320_ (\uc8051golden_1.IRAM[196] [6], _08348_, clk);
  dff _55321_ (\uc8051golden_1.IRAM[196] [7], _08349_, clk);
  dff _55322_ (\uc8051golden_1.IRAM[197] [0], _08350_, clk);
  dff _55323_ (\uc8051golden_1.IRAM[197] [1], _08351_, clk);
  dff _55324_ (\uc8051golden_1.IRAM[197] [2], _08352_, clk);
  dff _55325_ (\uc8051golden_1.IRAM[197] [3], _08353_, clk);
  dff _55326_ (\uc8051golden_1.IRAM[197] [4], _08354_, clk);
  dff _55327_ (\uc8051golden_1.IRAM[197] [5], _08355_, clk);
  dff _55328_ (\uc8051golden_1.IRAM[197] [6], _08356_, clk);
  dff _55329_ (\uc8051golden_1.IRAM[197] [7], _08357_, clk);
  dff _55330_ (\uc8051golden_1.IRAM[198] [0], _08358_, clk);
  dff _55331_ (\uc8051golden_1.IRAM[198] [1], _08359_, clk);
  dff _55332_ (\uc8051golden_1.IRAM[198] [2], _08360_, clk);
  dff _55333_ (\uc8051golden_1.IRAM[198] [3], _08361_, clk);
  dff _55334_ (\uc8051golden_1.IRAM[198] [4], _08362_, clk);
  dff _55335_ (\uc8051golden_1.IRAM[198] [5], _08363_, clk);
  dff _55336_ (\uc8051golden_1.IRAM[198] [6], _08364_, clk);
  dff _55337_ (\uc8051golden_1.IRAM[198] [7], _08365_, clk);
  dff _55338_ (\uc8051golden_1.IRAM[199] [0], _08366_, clk);
  dff _55339_ (\uc8051golden_1.IRAM[199] [1], _08367_, clk);
  dff _55340_ (\uc8051golden_1.IRAM[199] [2], _08368_, clk);
  dff _55341_ (\uc8051golden_1.IRAM[199] [3], _08369_, clk);
  dff _55342_ (\uc8051golden_1.IRAM[199] [4], _08370_, clk);
  dff _55343_ (\uc8051golden_1.IRAM[199] [5], _08371_, clk);
  dff _55344_ (\uc8051golden_1.IRAM[199] [6], _08372_, clk);
  dff _55345_ (\uc8051golden_1.IRAM[199] [7], _08373_, clk);
  dff _55346_ (\uc8051golden_1.IRAM[200] [0], _08374_, clk);
  dff _55347_ (\uc8051golden_1.IRAM[200] [1], _08375_, clk);
  dff _55348_ (\uc8051golden_1.IRAM[200] [2], _08376_, clk);
  dff _55349_ (\uc8051golden_1.IRAM[200] [3], _08377_, clk);
  dff _55350_ (\uc8051golden_1.IRAM[200] [4], _08379_, clk);
  dff _55351_ (\uc8051golden_1.IRAM[200] [5], _08380_, clk);
  dff _55352_ (\uc8051golden_1.IRAM[200] [6], _08381_, clk);
  dff _55353_ (\uc8051golden_1.IRAM[200] [7], _08382_, clk);
  dff _55354_ (\uc8051golden_1.IRAM[201] [0], _08383_, clk);
  dff _55355_ (\uc8051golden_1.IRAM[201] [1], _08384_, clk);
  dff _55356_ (\uc8051golden_1.IRAM[201] [2], _08385_, clk);
  dff _55357_ (\uc8051golden_1.IRAM[201] [3], _08386_, clk);
  dff _55358_ (\uc8051golden_1.IRAM[201] [4], _08387_, clk);
  dff _55359_ (\uc8051golden_1.IRAM[201] [5], _08388_, clk);
  dff _55360_ (\uc8051golden_1.IRAM[201] [6], _08389_, clk);
  dff _55361_ (\uc8051golden_1.IRAM[201] [7], _08390_, clk);
  dff _55362_ (\uc8051golden_1.IRAM[202] [0], _08391_, clk);
  dff _55363_ (\uc8051golden_1.IRAM[202] [1], _08392_, clk);
  dff _55364_ (\uc8051golden_1.IRAM[202] [2], _08393_, clk);
  dff _55365_ (\uc8051golden_1.IRAM[202] [3], _08394_, clk);
  dff _55366_ (\uc8051golden_1.IRAM[202] [4], _08395_, clk);
  dff _55367_ (\uc8051golden_1.IRAM[202] [5], _08396_, clk);
  dff _55368_ (\uc8051golden_1.IRAM[202] [6], _08397_, clk);
  dff _55369_ (\uc8051golden_1.IRAM[202] [7], _08398_, clk);
  dff _55370_ (\uc8051golden_1.IRAM[203] [0], _08399_, clk);
  dff _55371_ (\uc8051golden_1.IRAM[203] [1], _08400_, clk);
  dff _55372_ (\uc8051golden_1.IRAM[203] [2], _08401_, clk);
  dff _55373_ (\uc8051golden_1.IRAM[203] [3], _08402_, clk);
  dff _55374_ (\uc8051golden_1.IRAM[203] [4], _08403_, clk);
  dff _55375_ (\uc8051golden_1.IRAM[203] [5], _08404_, clk);
  dff _55376_ (\uc8051golden_1.IRAM[203] [6], _08405_, clk);
  dff _55377_ (\uc8051golden_1.IRAM[203] [7], _08406_, clk);
  dff _55378_ (\uc8051golden_1.IRAM[204] [0], _08407_, clk);
  dff _55379_ (\uc8051golden_1.IRAM[204] [1], _08408_, clk);
  dff _55380_ (\uc8051golden_1.IRAM[204] [2], _08409_, clk);
  dff _55381_ (\uc8051golden_1.IRAM[204] [3], _08410_, clk);
  dff _55382_ (\uc8051golden_1.IRAM[204] [4], _08411_, clk);
  dff _55383_ (\uc8051golden_1.IRAM[204] [5], _08413_, clk);
  dff _55384_ (\uc8051golden_1.IRAM[204] [6], _08414_, clk);
  dff _55385_ (\uc8051golden_1.IRAM[204] [7], _08415_, clk);
  dff _55386_ (\uc8051golden_1.IRAM[205] [0], _08416_, clk);
  dff _55387_ (\uc8051golden_1.IRAM[205] [1], _08417_, clk);
  dff _55388_ (\uc8051golden_1.IRAM[205] [2], _08418_, clk);
  dff _55389_ (\uc8051golden_1.IRAM[205] [3], _08419_, clk);
  dff _55390_ (\uc8051golden_1.IRAM[205] [4], _08420_, clk);
  dff _55391_ (\uc8051golden_1.IRAM[205] [5], _08421_, clk);
  dff _55392_ (\uc8051golden_1.IRAM[205] [6], _08422_, clk);
  dff _55393_ (\uc8051golden_1.IRAM[205] [7], _08423_, clk);
  dff _55394_ (\uc8051golden_1.IRAM[206] [0], _08424_, clk);
  dff _55395_ (\uc8051golden_1.IRAM[206] [1], _08425_, clk);
  dff _55396_ (\uc8051golden_1.IRAM[206] [2], _08426_, clk);
  dff _55397_ (\uc8051golden_1.IRAM[206] [3], _08427_, clk);
  dff _55398_ (\uc8051golden_1.IRAM[206] [4], _08428_, clk);
  dff _55399_ (\uc8051golden_1.IRAM[206] [5], _08429_, clk);
  dff _55400_ (\uc8051golden_1.IRAM[206] [6], _08430_, clk);
  dff _55401_ (\uc8051golden_1.IRAM[206] [7], _08431_, clk);
  dff _55402_ (\uc8051golden_1.IRAM[207] [0], _08432_, clk);
  dff _55403_ (\uc8051golden_1.IRAM[207] [1], _08433_, clk);
  dff _55404_ (\uc8051golden_1.IRAM[207] [2], _08434_, clk);
  dff _55405_ (\uc8051golden_1.IRAM[207] [3], _08435_, clk);
  dff _55406_ (\uc8051golden_1.IRAM[207] [4], _08436_, clk);
  dff _55407_ (\uc8051golden_1.IRAM[207] [5], _08437_, clk);
  dff _55408_ (\uc8051golden_1.IRAM[207] [6], _08438_, clk);
  dff _55409_ (\uc8051golden_1.IRAM[207] [7], _08439_, clk);
  dff _55410_ (\uc8051golden_1.IRAM[208] [0], _08440_, clk);
  dff _55411_ (\uc8051golden_1.IRAM[208] [1], _08441_, clk);
  dff _55412_ (\uc8051golden_1.IRAM[208] [2], _08442_, clk);
  dff _55413_ (\uc8051golden_1.IRAM[208] [3], _08443_, clk);
  dff _55414_ (\uc8051golden_1.IRAM[208] [4], _08444_, clk);
  dff _55415_ (\uc8051golden_1.IRAM[208] [5], _08445_, clk);
  dff _55416_ (\uc8051golden_1.IRAM[208] [6], _08447_, clk);
  dff _55417_ (\uc8051golden_1.IRAM[208] [7], _08448_, clk);
  dff _55418_ (\uc8051golden_1.IRAM[209] [0], _08449_, clk);
  dff _55419_ (\uc8051golden_1.IRAM[209] [1], _08450_, clk);
  dff _55420_ (\uc8051golden_1.IRAM[209] [2], _08451_, clk);
  dff _55421_ (\uc8051golden_1.IRAM[209] [3], _08452_, clk);
  dff _55422_ (\uc8051golden_1.IRAM[209] [4], _08453_, clk);
  dff _55423_ (\uc8051golden_1.IRAM[209] [5], _08454_, clk);
  dff _55424_ (\uc8051golden_1.IRAM[209] [6], _08455_, clk);
  dff _55425_ (\uc8051golden_1.IRAM[209] [7], _08456_, clk);
  dff _55426_ (\uc8051golden_1.IRAM[210] [0], _08457_, clk);
  dff _55427_ (\uc8051golden_1.IRAM[210] [1], _08458_, clk);
  dff _55428_ (\uc8051golden_1.IRAM[210] [2], _08459_, clk);
  dff _55429_ (\uc8051golden_1.IRAM[210] [3], _08460_, clk);
  dff _55430_ (\uc8051golden_1.IRAM[210] [4], _08461_, clk);
  dff _55431_ (\uc8051golden_1.IRAM[210] [5], _08462_, clk);
  dff _55432_ (\uc8051golden_1.IRAM[210] [6], _08463_, clk);
  dff _55433_ (\uc8051golden_1.IRAM[210] [7], _08464_, clk);
  dff _55434_ (\uc8051golden_1.IRAM[211] [0], _08465_, clk);
  dff _55435_ (\uc8051golden_1.IRAM[211] [1], _08466_, clk);
  dff _55436_ (\uc8051golden_1.IRAM[211] [2], _08467_, clk);
  dff _55437_ (\uc8051golden_1.IRAM[211] [3], _08468_, clk);
  dff _55438_ (\uc8051golden_1.IRAM[211] [4], _08469_, clk);
  dff _55439_ (\uc8051golden_1.IRAM[211] [5], _08470_, clk);
  dff _55440_ (\uc8051golden_1.IRAM[211] [6], _08471_, clk);
  dff _55441_ (\uc8051golden_1.IRAM[211] [7], _08472_, clk);
  dff _55442_ (\uc8051golden_1.IRAM[212] [0], _08473_, clk);
  dff _55443_ (\uc8051golden_1.IRAM[212] [1], _08474_, clk);
  dff _55444_ (\uc8051golden_1.IRAM[212] [2], _08475_, clk);
  dff _55445_ (\uc8051golden_1.IRAM[212] [3], _08476_, clk);
  dff _55446_ (\uc8051golden_1.IRAM[212] [4], _08477_, clk);
  dff _55447_ (\uc8051golden_1.IRAM[212] [5], _08478_, clk);
  dff _55448_ (\uc8051golden_1.IRAM[212] [6], _08479_, clk);
  dff _55449_ (\uc8051golden_1.IRAM[212] [7], _08480_, clk);
  dff _55450_ (\uc8051golden_1.IRAM[213] [0], _08482_, clk);
  dff _55451_ (\uc8051golden_1.IRAM[213] [1], _08483_, clk);
  dff _55452_ (\uc8051golden_1.IRAM[213] [2], _08484_, clk);
  dff _55453_ (\uc8051golden_1.IRAM[213] [3], _08485_, clk);
  dff _55454_ (\uc8051golden_1.IRAM[213] [4], _08486_, clk);
  dff _55455_ (\uc8051golden_1.IRAM[213] [5], _08487_, clk);
  dff _55456_ (\uc8051golden_1.IRAM[213] [6], _08488_, clk);
  dff _55457_ (\uc8051golden_1.IRAM[213] [7], _08489_, clk);
  dff _55458_ (\uc8051golden_1.IRAM[214] [0], _08490_, clk);
  dff _55459_ (\uc8051golden_1.IRAM[214] [1], _08491_, clk);
  dff _55460_ (\uc8051golden_1.IRAM[214] [2], _08492_, clk);
  dff _55461_ (\uc8051golden_1.IRAM[214] [3], _08493_, clk);
  dff _55462_ (\uc8051golden_1.IRAM[214] [4], _08494_, clk);
  dff _55463_ (\uc8051golden_1.IRAM[214] [5], _08495_, clk);
  dff _55464_ (\uc8051golden_1.IRAM[214] [6], _08496_, clk);
  dff _55465_ (\uc8051golden_1.IRAM[214] [7], _08497_, clk);
  dff _55466_ (\uc8051golden_1.IRAM[215] [0], _08498_, clk);
  dff _55467_ (\uc8051golden_1.IRAM[215] [1], _08499_, clk);
  dff _55468_ (\uc8051golden_1.IRAM[215] [2], _08500_, clk);
  dff _55469_ (\uc8051golden_1.IRAM[215] [3], _08501_, clk);
  dff _55470_ (\uc8051golden_1.IRAM[215] [4], _08502_, clk);
  dff _55471_ (\uc8051golden_1.IRAM[215] [5], _08503_, clk);
  dff _55472_ (\uc8051golden_1.IRAM[215] [6], _08504_, clk);
  dff _55473_ (\uc8051golden_1.IRAM[215] [7], _08505_, clk);
  dff _55474_ (\uc8051golden_1.IRAM[216] [0], _08506_, clk);
  dff _55475_ (\uc8051golden_1.IRAM[216] [1], _08507_, clk);
  dff _55476_ (\uc8051golden_1.IRAM[216] [2], _08508_, clk);
  dff _55477_ (\uc8051golden_1.IRAM[216] [3], _08509_, clk);
  dff _55478_ (\uc8051golden_1.IRAM[216] [4], _08510_, clk);
  dff _55479_ (\uc8051golden_1.IRAM[216] [5], _08511_, clk);
  dff _55480_ (\uc8051golden_1.IRAM[216] [6], _08512_, clk);
  dff _55481_ (\uc8051golden_1.IRAM[216] [7], _08513_, clk);
  dff _55482_ (\uc8051golden_1.IRAM[217] [0], _08514_, clk);
  dff _55483_ (\uc8051golden_1.IRAM[217] [1], _08516_, clk);
  dff _55484_ (\uc8051golden_1.IRAM[217] [2], _08517_, clk);
  dff _55485_ (\uc8051golden_1.IRAM[217] [3], _08518_, clk);
  dff _55486_ (\uc8051golden_1.IRAM[217] [4], _08519_, clk);
  dff _55487_ (\uc8051golden_1.IRAM[217] [5], _08520_, clk);
  dff _55488_ (\uc8051golden_1.IRAM[217] [6], _08521_, clk);
  dff _55489_ (\uc8051golden_1.IRAM[217] [7], _08522_, clk);
  dff _55490_ (\uc8051golden_1.IRAM[218] [0], _08523_, clk);
  dff _55491_ (\uc8051golden_1.IRAM[218] [1], _08524_, clk);
  dff _55492_ (\uc8051golden_1.IRAM[218] [2], _08525_, clk);
  dff _55493_ (\uc8051golden_1.IRAM[218] [3], _08526_, clk);
  dff _55494_ (\uc8051golden_1.IRAM[218] [4], _08527_, clk);
  dff _55495_ (\uc8051golden_1.IRAM[218] [5], _08528_, clk);
  dff _55496_ (\uc8051golden_1.IRAM[218] [6], _08529_, clk);
  dff _55497_ (\uc8051golden_1.IRAM[218] [7], _08530_, clk);
  dff _55498_ (\uc8051golden_1.IRAM[219] [0], _08531_, clk);
  dff _55499_ (\uc8051golden_1.IRAM[219] [1], _08532_, clk);
  dff _55500_ (\uc8051golden_1.IRAM[219] [2], _08533_, clk);
  dff _55501_ (\uc8051golden_1.IRAM[219] [3], _08534_, clk);
  dff _55502_ (\uc8051golden_1.IRAM[219] [4], _08535_, clk);
  dff _55503_ (\uc8051golden_1.IRAM[219] [5], _08536_, clk);
  dff _55504_ (\uc8051golden_1.IRAM[219] [6], _08537_, clk);
  dff _55505_ (\uc8051golden_1.IRAM[219] [7], _08538_, clk);
  dff _55506_ (\uc8051golden_1.IRAM[220] [0], _08539_, clk);
  dff _55507_ (\uc8051golden_1.IRAM[220] [1], _08540_, clk);
  dff _55508_ (\uc8051golden_1.IRAM[220] [2], _08541_, clk);
  dff _55509_ (\uc8051golden_1.IRAM[220] [3], _08542_, clk);
  dff _55510_ (\uc8051golden_1.IRAM[220] [4], _08543_, clk);
  dff _55511_ (\uc8051golden_1.IRAM[220] [5], _08544_, clk);
  dff _55512_ (\uc8051golden_1.IRAM[220] [6], _08545_, clk);
  dff _55513_ (\uc8051golden_1.IRAM[220] [7], _08546_, clk);
  dff _55514_ (\uc8051golden_1.IRAM[221] [0], _08547_, clk);
  dff _55515_ (\uc8051golden_1.IRAM[221] [1], _08548_, clk);
  dff _55516_ (\uc8051golden_1.IRAM[221] [2], _08550_, clk);
  dff _55517_ (\uc8051golden_1.IRAM[221] [3], _08551_, clk);
  dff _55518_ (\uc8051golden_1.IRAM[221] [4], _08552_, clk);
  dff _55519_ (\uc8051golden_1.IRAM[221] [5], _08553_, clk);
  dff _55520_ (\uc8051golden_1.IRAM[221] [6], _08554_, clk);
  dff _55521_ (\uc8051golden_1.IRAM[221] [7], _08555_, clk);
  dff _55522_ (\uc8051golden_1.IRAM[222] [0], _08556_, clk);
  dff _55523_ (\uc8051golden_1.IRAM[222] [1], _08557_, clk);
  dff _55524_ (\uc8051golden_1.IRAM[222] [2], _08558_, clk);
  dff _55525_ (\uc8051golden_1.IRAM[222] [3], _08559_, clk);
  dff _55526_ (\uc8051golden_1.IRAM[222] [4], _08560_, clk);
  dff _55527_ (\uc8051golden_1.IRAM[222] [5], _08561_, clk);
  dff _55528_ (\uc8051golden_1.IRAM[222] [6], _08562_, clk);
  dff _55529_ (\uc8051golden_1.IRAM[222] [7], _08563_, clk);
  dff _55530_ (\uc8051golden_1.IRAM[223] [0], _08564_, clk);
  dff _55531_ (\uc8051golden_1.IRAM[223] [1], _08565_, clk);
  dff _55532_ (\uc8051golden_1.IRAM[223] [2], _08566_, clk);
  dff _55533_ (\uc8051golden_1.IRAM[223] [3], _08567_, clk);
  dff _55534_ (\uc8051golden_1.IRAM[223] [4], _08568_, clk);
  dff _55535_ (\uc8051golden_1.IRAM[223] [5], _08569_, clk);
  dff _55536_ (\uc8051golden_1.IRAM[223] [6], _08570_, clk);
  dff _55537_ (\uc8051golden_1.IRAM[223] [7], _08571_, clk);
  dff _55538_ (\uc8051golden_1.IRAM[224] [0], _08572_, clk);
  dff _55539_ (\uc8051golden_1.IRAM[224] [1], _08573_, clk);
  dff _55540_ (\uc8051golden_1.IRAM[224] [2], _08574_, clk);
  dff _55541_ (\uc8051golden_1.IRAM[224] [3], _08575_, clk);
  dff _55542_ (\uc8051golden_1.IRAM[224] [4], _08576_, clk);
  dff _55543_ (\uc8051golden_1.IRAM[224] [5], _08577_, clk);
  dff _55544_ (\uc8051golden_1.IRAM[224] [6], _08578_, clk);
  dff _55545_ (\uc8051golden_1.IRAM[224] [7], _08579_, clk);
  dff _55546_ (\uc8051golden_1.IRAM[225] [0], _08580_, clk);
  dff _55547_ (\uc8051golden_1.IRAM[225] [1], _08581_, clk);
  dff _55548_ (\uc8051golden_1.IRAM[225] [2], _08582_, clk);
  dff _55549_ (\uc8051golden_1.IRAM[225] [3], _08584_, clk);
  dff _55550_ (\uc8051golden_1.IRAM[225] [4], _08585_, clk);
  dff _55551_ (\uc8051golden_1.IRAM[225] [5], _08586_, clk);
  dff _55552_ (\uc8051golden_1.IRAM[225] [6], _08587_, clk);
  dff _55553_ (\uc8051golden_1.IRAM[225] [7], _08588_, clk);
  dff _55554_ (\uc8051golden_1.IRAM[226] [0], _08589_, clk);
  dff _55555_ (\uc8051golden_1.IRAM[226] [1], _08590_, clk);
  dff _55556_ (\uc8051golden_1.IRAM[226] [2], _08591_, clk);
  dff _55557_ (\uc8051golden_1.IRAM[226] [3], _08592_, clk);
  dff _55558_ (\uc8051golden_1.IRAM[226] [4], _08593_, clk);
  dff _55559_ (\uc8051golden_1.IRAM[226] [5], _08594_, clk);
  dff _55560_ (\uc8051golden_1.IRAM[226] [6], _08595_, clk);
  dff _55561_ (\uc8051golden_1.IRAM[226] [7], _08596_, clk);
  dff _55562_ (\uc8051golden_1.IRAM[227] [0], _08597_, clk);
  dff _55563_ (\uc8051golden_1.IRAM[227] [1], _08598_, clk);
  dff _55564_ (\uc8051golden_1.IRAM[227] [2], _08599_, clk);
  dff _55565_ (\uc8051golden_1.IRAM[227] [3], _08600_, clk);
  dff _55566_ (\uc8051golden_1.IRAM[227] [4], _08601_, clk);
  dff _55567_ (\uc8051golden_1.IRAM[227] [5], _08602_, clk);
  dff _55568_ (\uc8051golden_1.IRAM[227] [6], _08603_, clk);
  dff _55569_ (\uc8051golden_1.IRAM[227] [7], _08604_, clk);
  dff _55570_ (\uc8051golden_1.IRAM[228] [0], _08605_, clk);
  dff _55571_ (\uc8051golden_1.IRAM[228] [1], _08606_, clk);
  dff _55572_ (\uc8051golden_1.IRAM[228] [2], _08607_, clk);
  dff _55573_ (\uc8051golden_1.IRAM[228] [3], _08608_, clk);
  dff _55574_ (\uc8051golden_1.IRAM[228] [4], _08609_, clk);
  dff _55575_ (\uc8051golden_1.IRAM[228] [5], _08610_, clk);
  dff _55576_ (\uc8051golden_1.IRAM[228] [6], _08611_, clk);
  dff _55577_ (\uc8051golden_1.IRAM[228] [7], _08612_, clk);
  dff _55578_ (\uc8051golden_1.IRAM[229] [0], _08613_, clk);
  dff _55579_ (\uc8051golden_1.IRAM[229] [1], _08614_, clk);
  dff _55580_ (\uc8051golden_1.IRAM[229] [2], _08615_, clk);
  dff _55581_ (\uc8051golden_1.IRAM[229] [3], _08616_, clk);
  dff _55582_ (\uc8051golden_1.IRAM[229] [4], _08618_, clk);
  dff _55583_ (\uc8051golden_1.IRAM[229] [5], _08619_, clk);
  dff _55584_ (\uc8051golden_1.IRAM[229] [6], _08620_, clk);
  dff _55585_ (\uc8051golden_1.IRAM[229] [7], _08621_, clk);
  dff _55586_ (\uc8051golden_1.IRAM[230] [0], _08622_, clk);
  dff _55587_ (\uc8051golden_1.IRAM[230] [1], _08623_, clk);
  dff _55588_ (\uc8051golden_1.IRAM[230] [2], _08624_, clk);
  dff _55589_ (\uc8051golden_1.IRAM[230] [3], _08625_, clk);
  dff _55590_ (\uc8051golden_1.IRAM[230] [4], _08626_, clk);
  dff _55591_ (\uc8051golden_1.IRAM[230] [5], _08627_, clk);
  dff _55592_ (\uc8051golden_1.IRAM[230] [6], _08628_, clk);
  dff _55593_ (\uc8051golden_1.IRAM[230] [7], _08629_, clk);
  dff _55594_ (\uc8051golden_1.IRAM[231] [0], _08630_, clk);
  dff _55595_ (\uc8051golden_1.IRAM[231] [1], _08631_, clk);
  dff _55596_ (\uc8051golden_1.IRAM[231] [2], _08632_, clk);
  dff _55597_ (\uc8051golden_1.IRAM[231] [3], _08633_, clk);
  dff _55598_ (\uc8051golden_1.IRAM[231] [4], _08634_, clk);
  dff _55599_ (\uc8051golden_1.IRAM[231] [5], _08635_, clk);
  dff _55600_ (\uc8051golden_1.IRAM[231] [6], _08636_, clk);
  dff _55601_ (\uc8051golden_1.IRAM[231] [7], _08637_, clk);
  dff _55602_ (\uc8051golden_1.IRAM[232] [0], _08638_, clk);
  dff _55603_ (\uc8051golden_1.IRAM[232] [1], _08639_, clk);
  dff _55604_ (\uc8051golden_1.IRAM[232] [2], _08640_, clk);
  dff _55605_ (\uc8051golden_1.IRAM[232] [3], _08641_, clk);
  dff _55606_ (\uc8051golden_1.IRAM[232] [4], _08642_, clk);
  dff _55607_ (\uc8051golden_1.IRAM[232] [5], _08643_, clk);
  dff _55608_ (\uc8051golden_1.IRAM[232] [6], _08644_, clk);
  dff _55609_ (\uc8051golden_1.IRAM[232] [7], _08645_, clk);
  dff _55610_ (\uc8051golden_1.IRAM[233] [0], _08646_, clk);
  dff _55611_ (\uc8051golden_1.IRAM[233] [1], _08647_, clk);
  dff _55612_ (\uc8051golden_1.IRAM[233] [2], _08648_, clk);
  dff _55613_ (\uc8051golden_1.IRAM[233] [3], _08649_, clk);
  dff _55614_ (\uc8051golden_1.IRAM[233] [4], _08650_, clk);
  dff _55615_ (\uc8051golden_1.IRAM[233] [5], _08651_, clk);
  dff _55616_ (\uc8051golden_1.IRAM[233] [6], _08653_, clk);
  dff _55617_ (\uc8051golden_1.IRAM[233] [7], _08654_, clk);
  dff _55618_ (\uc8051golden_1.IRAM[234] [0], _08655_, clk);
  dff _55619_ (\uc8051golden_1.IRAM[234] [1], _08656_, clk);
  dff _55620_ (\uc8051golden_1.IRAM[234] [2], _08657_, clk);
  dff _55621_ (\uc8051golden_1.IRAM[234] [3], _08658_, clk);
  dff _55622_ (\uc8051golden_1.IRAM[234] [4], _08659_, clk);
  dff _55623_ (\uc8051golden_1.IRAM[234] [5], _08660_, clk);
  dff _55624_ (\uc8051golden_1.IRAM[234] [6], _08661_, clk);
  dff _55625_ (\uc8051golden_1.IRAM[234] [7], _08662_, clk);
  dff _55626_ (\uc8051golden_1.IRAM[235] [0], _08663_, clk);
  dff _55627_ (\uc8051golden_1.IRAM[235] [1], _08664_, clk);
  dff _55628_ (\uc8051golden_1.IRAM[235] [2], _08665_, clk);
  dff _55629_ (\uc8051golden_1.IRAM[235] [3], _08666_, clk);
  dff _55630_ (\uc8051golden_1.IRAM[235] [4], _08667_, clk);
  dff _55631_ (\uc8051golden_1.IRAM[235] [5], _08668_, clk);
  dff _55632_ (\uc8051golden_1.IRAM[235] [6], _08669_, clk);
  dff _55633_ (\uc8051golden_1.IRAM[235] [7], _08670_, clk);
  dff _55634_ (\uc8051golden_1.IRAM[236] [0], _08671_, clk);
  dff _55635_ (\uc8051golden_1.IRAM[236] [1], _08672_, clk);
  dff _55636_ (\uc8051golden_1.IRAM[236] [2], _08673_, clk);
  dff _55637_ (\uc8051golden_1.IRAM[236] [3], _08674_, clk);
  dff _55638_ (\uc8051golden_1.IRAM[236] [4], _08675_, clk);
  dff _55639_ (\uc8051golden_1.IRAM[236] [5], _08676_, clk);
  dff _55640_ (\uc8051golden_1.IRAM[236] [6], _08677_, clk);
  dff _55641_ (\uc8051golden_1.IRAM[236] [7], _08678_, clk);
  dff _55642_ (\uc8051golden_1.IRAM[237] [0], _08679_, clk);
  dff _55643_ (\uc8051golden_1.IRAM[237] [1], _08680_, clk);
  dff _55644_ (\uc8051golden_1.IRAM[237] [2], _08681_, clk);
  dff _55645_ (\uc8051golden_1.IRAM[237] [3], _08682_, clk);
  dff _55646_ (\uc8051golden_1.IRAM[237] [4], _08683_, clk);
  dff _55647_ (\uc8051golden_1.IRAM[237] [5], _08684_, clk);
  dff _55648_ (\uc8051golden_1.IRAM[237] [6], _08685_, clk);
  dff _55649_ (\uc8051golden_1.IRAM[237] [7], _08687_, clk);
  dff _55650_ (\uc8051golden_1.IRAM[238] [0], _08688_, clk);
  dff _55651_ (\uc8051golden_1.IRAM[238] [1], _08689_, clk);
  dff _55652_ (\uc8051golden_1.IRAM[238] [2], _08690_, clk);
  dff _55653_ (\uc8051golden_1.IRAM[238] [3], _08691_, clk);
  dff _55654_ (\uc8051golden_1.IRAM[238] [4], _08692_, clk);
  dff _55655_ (\uc8051golden_1.IRAM[238] [5], _08693_, clk);
  dff _55656_ (\uc8051golden_1.IRAM[238] [6], _08694_, clk);
  dff _55657_ (\uc8051golden_1.IRAM[238] [7], _08695_, clk);
  dff _55658_ (\uc8051golden_1.IRAM[239] [0], _08696_, clk);
  dff _55659_ (\uc8051golden_1.IRAM[239] [1], _08697_, clk);
  dff _55660_ (\uc8051golden_1.IRAM[239] [2], _08698_, clk);
  dff _55661_ (\uc8051golden_1.IRAM[239] [3], _08699_, clk);
  dff _55662_ (\uc8051golden_1.IRAM[239] [4], _08700_, clk);
  dff _55663_ (\uc8051golden_1.IRAM[239] [5], _08701_, clk);
  dff _55664_ (\uc8051golden_1.IRAM[239] [6], _08702_, clk);
  dff _55665_ (\uc8051golden_1.IRAM[239] [7], _08703_, clk);
  dff _55666_ (\uc8051golden_1.IRAM[240] [0], _08704_, clk);
  dff _55667_ (\uc8051golden_1.IRAM[240] [1], _08705_, clk);
  dff _55668_ (\uc8051golden_1.IRAM[240] [2], _08706_, clk);
  dff _55669_ (\uc8051golden_1.IRAM[240] [3], _08707_, clk);
  dff _55670_ (\uc8051golden_1.IRAM[240] [4], _08708_, clk);
  dff _55671_ (\uc8051golden_1.IRAM[240] [5], _08709_, clk);
  dff _55672_ (\uc8051golden_1.IRAM[240] [6], _08710_, clk);
  dff _55673_ (\uc8051golden_1.IRAM[240] [7], _08711_, clk);
  dff _55674_ (\uc8051golden_1.IRAM[241] [0], _08712_, clk);
  dff _55675_ (\uc8051golden_1.IRAM[241] [1], _08713_, clk);
  dff _55676_ (\uc8051golden_1.IRAM[241] [2], _08714_, clk);
  dff _55677_ (\uc8051golden_1.IRAM[241] [3], _08715_, clk);
  dff _55678_ (\uc8051golden_1.IRAM[241] [4], _08716_, clk);
  dff _55679_ (\uc8051golden_1.IRAM[241] [5], _08717_, clk);
  dff _55680_ (\uc8051golden_1.IRAM[241] [6], _08718_, clk);
  dff _55681_ (\uc8051golden_1.IRAM[241] [7], _08719_, clk);
  dff _55682_ (\uc8051golden_1.IRAM[242] [0], _08721_, clk);
  dff _55683_ (\uc8051golden_1.IRAM[242] [1], _08722_, clk);
  dff _55684_ (\uc8051golden_1.IRAM[242] [2], _08723_, clk);
  dff _55685_ (\uc8051golden_1.IRAM[242] [3], _08724_, clk);
  dff _55686_ (\uc8051golden_1.IRAM[242] [4], _08725_, clk);
  dff _55687_ (\uc8051golden_1.IRAM[242] [5], _08726_, clk);
  dff _55688_ (\uc8051golden_1.IRAM[242] [6], _08727_, clk);
  dff _55689_ (\uc8051golden_1.IRAM[242] [7], _08728_, clk);
  dff _55690_ (\uc8051golden_1.IRAM[243] [0], _08729_, clk);
  dff _55691_ (\uc8051golden_1.IRAM[243] [1], _08730_, clk);
  dff _55692_ (\uc8051golden_1.IRAM[243] [2], _08731_, clk);
  dff _55693_ (\uc8051golden_1.IRAM[243] [3], _08732_, clk);
  dff _55694_ (\uc8051golden_1.IRAM[243] [4], _08733_, clk);
  dff _55695_ (\uc8051golden_1.IRAM[243] [5], _08734_, clk);
  dff _55696_ (\uc8051golden_1.IRAM[243] [6], _08735_, clk);
  dff _55697_ (\uc8051golden_1.IRAM[243] [7], _08736_, clk);
  dff _55698_ (\uc8051golden_1.IRAM[244] [0], _08737_, clk);
  dff _55699_ (\uc8051golden_1.IRAM[244] [1], _08738_, clk);
  dff _55700_ (\uc8051golden_1.IRAM[244] [2], _08739_, clk);
  dff _55701_ (\uc8051golden_1.IRAM[244] [3], _08740_, clk);
  dff _55702_ (\uc8051golden_1.IRAM[244] [4], _08741_, clk);
  dff _55703_ (\uc8051golden_1.IRAM[244] [5], _08742_, clk);
  dff _55704_ (\uc8051golden_1.IRAM[244] [6], _08743_, clk);
  dff _55705_ (\uc8051golden_1.IRAM[244] [7], _08744_, clk);
  dff _55706_ (\uc8051golden_1.IRAM[245] [0], _08745_, clk);
  dff _55707_ (\uc8051golden_1.IRAM[245] [1], _08746_, clk);
  dff _55708_ (\uc8051golden_1.IRAM[245] [2], _08747_, clk);
  dff _55709_ (\uc8051golden_1.IRAM[245] [3], _08748_, clk);
  dff _55710_ (\uc8051golden_1.IRAM[245] [4], _08749_, clk);
  dff _55711_ (\uc8051golden_1.IRAM[245] [5], _08750_, clk);
  dff _55712_ (\uc8051golden_1.IRAM[245] [6], _08751_, clk);
  dff _55713_ (\uc8051golden_1.IRAM[245] [7], _08752_, clk);
  dff _55714_ (\uc8051golden_1.IRAM[246] [0], _08753_, clk);
  dff _55715_ (\uc8051golden_1.IRAM[246] [1], _08755_, clk);
  dff _55716_ (\uc8051golden_1.IRAM[246] [2], _08756_, clk);
  dff _55717_ (\uc8051golden_1.IRAM[246] [3], _08757_, clk);
  dff _55718_ (\uc8051golden_1.IRAM[246] [4], _08758_, clk);
  dff _55719_ (\uc8051golden_1.IRAM[246] [5], _08759_, clk);
  dff _55720_ (\uc8051golden_1.IRAM[246] [6], _08760_, clk);
  dff _55721_ (\uc8051golden_1.IRAM[246] [7], _08761_, clk);
  dff _55722_ (\uc8051golden_1.IRAM[247] [0], _08762_, clk);
  dff _55723_ (\uc8051golden_1.IRAM[247] [1], _08763_, clk);
  dff _55724_ (\uc8051golden_1.IRAM[247] [2], _08764_, clk);
  dff _55725_ (\uc8051golden_1.IRAM[247] [3], _08765_, clk);
  dff _55726_ (\uc8051golden_1.IRAM[247] [4], _08766_, clk);
  dff _55727_ (\uc8051golden_1.IRAM[247] [5], _08767_, clk);
  dff _55728_ (\uc8051golden_1.IRAM[247] [6], _08768_, clk);
  dff _55729_ (\uc8051golden_1.IRAM[247] [7], _08769_, clk);
  dff _55730_ (\uc8051golden_1.IRAM[248] [0], _08770_, clk);
  dff _55731_ (\uc8051golden_1.IRAM[248] [1], _08771_, clk);
  dff _55732_ (\uc8051golden_1.IRAM[248] [2], _08772_, clk);
  dff _55733_ (\uc8051golden_1.IRAM[248] [3], _08773_, clk);
  dff _55734_ (\uc8051golden_1.IRAM[248] [4], _08774_, clk);
  dff _55735_ (\uc8051golden_1.IRAM[248] [5], _08775_, clk);
  dff _55736_ (\uc8051golden_1.IRAM[248] [6], _08776_, clk);
  dff _55737_ (\uc8051golden_1.IRAM[248] [7], _08777_, clk);
  dff _55738_ (\uc8051golden_1.IRAM[249] [0], _08778_, clk);
  dff _55739_ (\uc8051golden_1.IRAM[249] [1], _08779_, clk);
  dff _55740_ (\uc8051golden_1.IRAM[249] [2], _08780_, clk);
  dff _55741_ (\uc8051golden_1.IRAM[249] [3], _08781_, clk);
  dff _55742_ (\uc8051golden_1.IRAM[249] [4], _08782_, clk);
  dff _55743_ (\uc8051golden_1.IRAM[249] [5], _08783_, clk);
  dff _55744_ (\uc8051golden_1.IRAM[249] [6], _08784_, clk);
  dff _55745_ (\uc8051golden_1.IRAM[249] [7], _08785_, clk);
  dff _55746_ (\uc8051golden_1.IRAM[250] [0], _08786_, clk);
  dff _55747_ (\uc8051golden_1.IRAM[250] [1], _08787_, clk);
  dff _55748_ (\uc8051golden_1.IRAM[250] [2], _08788_, clk);
  dff _55749_ (\uc8051golden_1.IRAM[250] [3], _08790_, clk);
  dff _55750_ (\uc8051golden_1.IRAM[250] [4], _08791_, clk);
  dff _55751_ (\uc8051golden_1.IRAM[250] [5], _08792_, clk);
  dff _55752_ (\uc8051golden_1.IRAM[250] [6], _08793_, clk);
  dff _55753_ (\uc8051golden_1.IRAM[250] [7], _08794_, clk);
  dff _55754_ (\uc8051golden_1.IRAM[251] [0], _08795_, clk);
  dff _55755_ (\uc8051golden_1.IRAM[251] [1], _08796_, clk);
  dff _55756_ (\uc8051golden_1.IRAM[251] [2], _08797_, clk);
  dff _55757_ (\uc8051golden_1.IRAM[251] [3], _08798_, clk);
  dff _55758_ (\uc8051golden_1.IRAM[251] [4], _08799_, clk);
  dff _55759_ (\uc8051golden_1.IRAM[251] [5], _08800_, clk);
  dff _55760_ (\uc8051golden_1.IRAM[251] [6], _08801_, clk);
  dff _55761_ (\uc8051golden_1.IRAM[251] [7], _08802_, clk);
  dff _55762_ (\uc8051golden_1.IRAM[252] [0], _08803_, clk);
  dff _55763_ (\uc8051golden_1.IRAM[252] [1], _08804_, clk);
  dff _55764_ (\uc8051golden_1.IRAM[252] [2], _08805_, clk);
  dff _55765_ (\uc8051golden_1.IRAM[252] [3], _08806_, clk);
  dff _55766_ (\uc8051golden_1.IRAM[252] [4], _08807_, clk);
  dff _55767_ (\uc8051golden_1.IRAM[252] [5], _08808_, clk);
  dff _55768_ (\uc8051golden_1.IRAM[252] [6], _08809_, clk);
  dff _55769_ (\uc8051golden_1.IRAM[252] [7], _08810_, clk);
  dff _55770_ (\uc8051golden_1.IRAM[253] [0], _08811_, clk);
  dff _55771_ (\uc8051golden_1.IRAM[253] [1], _08812_, clk);
  dff _55772_ (\uc8051golden_1.IRAM[253] [2], _08813_, clk);
  dff _55773_ (\uc8051golden_1.IRAM[253] [3], _08814_, clk);
  dff _55774_ (\uc8051golden_1.IRAM[253] [4], _08815_, clk);
  dff _55775_ (\uc8051golden_1.IRAM[253] [5], _08816_, clk);
  dff _55776_ (\uc8051golden_1.IRAM[253] [6], _08817_, clk);
  dff _55777_ (\uc8051golden_1.IRAM[253] [7], _08818_, clk);
  dff _55778_ (\uc8051golden_1.IRAM[254] [0], _08819_, clk);
  dff _55779_ (\uc8051golden_1.IRAM[254] [1], _08820_, clk);
  dff _55780_ (\uc8051golden_1.IRAM[254] [2], _08821_, clk);
  dff _55781_ (\uc8051golden_1.IRAM[254] [3], _08822_, clk);
  dff _55782_ (\uc8051golden_1.IRAM[254] [4], _08824_, clk);
  dff _55783_ (\uc8051golden_1.IRAM[254] [5], _08825_, clk);
  dff _55784_ (\uc8051golden_1.IRAM[254] [6], _08826_, clk);
  dff _55785_ (\uc8051golden_1.IRAM[254] [7], _08827_, clk);
  dff _55786_ (\uc8051golden_1.IRAM[255] [0], _08828_, clk);
  dff _55787_ (\uc8051golden_1.IRAM[255] [1], _08829_, clk);
  dff _55788_ (\uc8051golden_1.IRAM[255] [2], _08830_, clk);
  dff _55789_ (\uc8051golden_1.IRAM[255] [3], _08831_, clk);
  dff _55790_ (\uc8051golden_1.IRAM[255] [4], _08832_, clk);
  dff _55791_ (\uc8051golden_1.IRAM[255] [5], _08833_, clk);
  dff _55792_ (\uc8051golden_1.IRAM[255] [6], _08834_, clk);
  dff _55793_ (\uc8051golden_1.IRAM[255] [7], _06583_, clk);
  dff _55794_ (_06719_, _09422_, clk);
  dff _55795_ (_06717_, _09423_, clk);
  dff _55796_ (_06715_, _09424_, clk);
  dff _55797_ (_06714_, _09425_, clk);
  dff _55798_ (_06713_, _09426_, clk);
  dff _55799_ (_06712_, _09427_, clk);
  dff _55800_ (_06711_, _09428_, clk);
  dff _55801_ (_06710_, _06604_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\uc8051golden_1.clk , clk);
  buf(\uc8051golden_1.rst , rst);
  buf(\uc8051golden_1.ACC_03 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_03 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_03 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_03 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_03 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_03 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_03 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_03 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_13 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_13 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_13 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_13 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_13 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_13 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_13 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_13 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.ACC_23 [0], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_23 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_23 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_23 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_23 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_23 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_23 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_23 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_33 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.ACC_33 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_33 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_33 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_33 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_33 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_33 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_33 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_c4 [0], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_c4 [1], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_c4 [2], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_c4 [3], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_c4 [4], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.ACC_c4 [5], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.ACC_c4 [6], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.ACC_c4 [7], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.ACC_d6 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.ACC_d6 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.ACC_d6 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.ACC_d6 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.ACC_d6 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_d6 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_d6 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_d6 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_d7 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.ACC_d7 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.ACC_d7 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.ACC_d7 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.ACC_d7 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.ACC_d7 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.ACC_d7 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.ACC_d7 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.ACC_e6 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.ACC_e6 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.ACC_e6 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.ACC_e6 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.ACC_e6 [4], \uc8051golden_1.ACC_c6 [4]);
  buf(\uc8051golden_1.ACC_e6 [5], \uc8051golden_1.ACC_c6 [5]);
  buf(\uc8051golden_1.ACC_e6 [6], \uc8051golden_1.ACC_c6 [6]);
  buf(\uc8051golden_1.ACC_e6 [7], \uc8051golden_1.ACC_c6 [7]);
  buf(\uc8051golden_1.ACC_e7 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.ACC_e7 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.ACC_e7 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.ACC_e7 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.ACC_e7 [4], \uc8051golden_1.ACC_c7 [4]);
  buf(\uc8051golden_1.ACC_e7 [5], \uc8051golden_1.ACC_c7 [5]);
  buf(\uc8051golden_1.ACC_e7 [6], \uc8051golden_1.ACC_c7 [6]);
  buf(\uc8051golden_1.ACC_e7 [7], \uc8051golden_1.ACC_c7 [7]);
  buf(\uc8051golden_1.PSW_0d [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_0d [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_0d [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_0d [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_0d [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_0d [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_0d [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_0d [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.PSW_13 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_13 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_13 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_13 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_13 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_13 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_13 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_13 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.PSW_24 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_24 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_24 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_24 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_24 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_25 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_25 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_25 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_25 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_25 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_26 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_26 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_26 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_26 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_26 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_27 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_27 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_27 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_27 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_27 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_28 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_28 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_28 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_28 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_28 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_29 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_29 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_29 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_29 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_29 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2a [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2a [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2a [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2a [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2a [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2b [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2b [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2b [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2b [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2b [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2c [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2c [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2c [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2c [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2c [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2d [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2d [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2d [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2d [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2d [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2e [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2e [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2e [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2e [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2e [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_2f [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_2f [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_2f [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_2f [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_2f [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_33 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_33 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_33 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_33 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_33 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_33 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_33 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_33 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.PSW_34 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_34 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_34 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_34 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_34 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_35 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_35 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_35 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_35 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_35 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_36 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_36 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_36 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_36 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_36 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_37 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_37 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_37 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_37 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_37 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_38 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_38 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_38 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_38 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_38 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_39 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_39 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_39 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_39 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_39 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3a [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3a [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3a [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3a [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3a [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3b [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3b [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3b [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3b [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3b [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3c [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3c [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3c [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3c [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3c [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3d [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3d [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3d [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3d [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3d [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3e [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3e [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3e [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3e [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3e [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_3f [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_3f [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_3f [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_3f [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_3f [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_46 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_46 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_46 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_46 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_46 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_46 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_46 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_46 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.PSW_65 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_65 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_65 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_65 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_65 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_65 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_65 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_65 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.PSW_72 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_72 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_72 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_72 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_72 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_72 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_72 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_82 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_82 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_82 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_82 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_82 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_82 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_82 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_84 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_84 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_84 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_84 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_84 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_84 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_84 [7], 1'b0);
  buf(\uc8051golden_1.PSW_94 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_94 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_94 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_94 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_94 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_95 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_95 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_95 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_95 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_95 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_96 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_96 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_96 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_96 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_96 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_97 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_97 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_97 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_97 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_97 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_98 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_98 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_98 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_98 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_98 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_99 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_99 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_99 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_99 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_99 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9a [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9a [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9a [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9a [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9a [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9b [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9b [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9b [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9b [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9b [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9c [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9c [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9c [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9c [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9c [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9d [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9d [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9d [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9d [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9d [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9e [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9e [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9e [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9e [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9e [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_9f [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_9f [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_9f [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_9f [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_9f [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_a0 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_a0 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_a0 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_a0 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_a0 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_a0 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_a0 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_a2 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_a2 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_a2 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_a2 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_a2 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_a2 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_a2 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_a4 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_a4 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_a4 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_a4 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_a4 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_a4 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_a4 [7], 1'b0);
  buf(\uc8051golden_1.PSW_b0 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b0 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b0 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b0 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b0 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b0 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b0 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b3 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b3 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b3 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b3 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b3 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b3 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b3 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b4 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b4 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b4 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b4 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b4 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b4 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b4 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b5 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b5 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b5 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b5 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b5 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b5 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b5 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b6 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b6 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b6 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b6 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b6 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b6 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b6 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b7 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b7 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b7 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b7 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b7 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b7 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b7 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b8 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b8 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b8 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b8 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b8 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b8 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b8 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_b9 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_b9 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_b9 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_b9 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_b9 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_b9 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_b9 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_ba [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_ba [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_ba [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_ba [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_ba [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_ba [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_ba [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bb [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bb [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bb [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bb [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bb [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bb [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bb [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bc [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bc [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bc [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bc [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bc [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bc [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bc [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bd [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bd [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bd [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bd [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bd [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bd [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bd [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_be [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_be [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_be [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_be [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_be [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_be [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_be [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_bf [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_bf [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_bf [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_bf [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_bf [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_bf [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_bf [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_c0 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_c0 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_c0 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_c0 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_c0 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_c0 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_c0 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_c0 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.PSW_c3 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_c3 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_c3 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_c3 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_c3 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_c3 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_c3 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_c3 [7], 1'b0);
  buf(\uc8051golden_1.PSW_ce [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_ce [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_ce [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_ce [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_ce [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_ce [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_ce [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_ce [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.PSW_d3 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_d3 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_d3 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_d3 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_d3 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_d3 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_d3 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.PSW_d3 [7], 1'b1);
  buf(\uc8051golden_1.PSW_d4 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.PSW_d4 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.PSW_d4 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.PSW_d4 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.PSW_d4 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.PSW_d4 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.PSW_d4 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0014 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0014 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0014 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0014 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0014 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0014 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0014 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0014 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0109 [0], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0109 [1], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0110 [0], 1'b0);
  buf(\uc8051golden_1.n0110 [1], 1'b0);
  buf(\uc8051golden_1.n0110 [2], 1'b0);
  buf(\uc8051golden_1.n0110 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0110 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0110 [5], 1'b0);
  buf(\uc8051golden_1.n0110 [6], 1'b0);
  buf(\uc8051golden_1.n0110 [7], 1'b0);
  buf(\uc8051golden_1.n0112 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.n0112 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.n0112 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.n0112 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.n0112 [4], \uc8051golden_1.ACC_c6 [4]);
  buf(\uc8051golden_1.n0112 [5], \uc8051golden_1.ACC_c6 [5]);
  buf(\uc8051golden_1.n0112 [6], \uc8051golden_1.ACC_c6 [6]);
  buf(\uc8051golden_1.n0112 [7], \uc8051golden_1.ACC_c6 [7]);
  buf(\uc8051golden_1.n0115 [0], 1'b1);
  buf(\uc8051golden_1.n0115 [1], 1'b0);
  buf(\uc8051golden_1.n0115 [2], 1'b0);
  buf(\uc8051golden_1.n0115 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0115 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0115 [5], 1'b0);
  buf(\uc8051golden_1.n0115 [6], 1'b0);
  buf(\uc8051golden_1.n0115 [7], 1'b0);
  buf(\uc8051golden_1.n0117 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.n0117 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.n0117 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.n0117 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.n0117 [4], \uc8051golden_1.ACC_c7 [4]);
  buf(\uc8051golden_1.n0117 [5], \uc8051golden_1.ACC_c7 [5]);
  buf(\uc8051golden_1.n0117 [6], \uc8051golden_1.ACC_c7 [6]);
  buf(\uc8051golden_1.n0117 [7], \uc8051golden_1.ACC_c7 [7]);
  buf(\uc8051golden_1.n0124 [0], 1'b0);
  buf(\uc8051golden_1.n0124 [1], 1'b1);
  buf(\uc8051golden_1.n0124 [2], 1'b0);
  buf(\uc8051golden_1.n0124 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0124 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0124 [5], 1'b0);
  buf(\uc8051golden_1.n0124 [6], 1'b0);
  buf(\uc8051golden_1.n0124 [7], 1'b0);
  buf(\uc8051golden_1.n0128 [0], 1'b1);
  buf(\uc8051golden_1.n0128 [1], 1'b1);
  buf(\uc8051golden_1.n0128 [2], 1'b0);
  buf(\uc8051golden_1.n0128 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0128 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0128 [5], 1'b0);
  buf(\uc8051golden_1.n0128 [6], 1'b0);
  buf(\uc8051golden_1.n0128 [7], 1'b0);
  buf(\uc8051golden_1.n0132 [0], 1'b0);
  buf(\uc8051golden_1.n0132 [1], 1'b0);
  buf(\uc8051golden_1.n0132 [2], 1'b1);
  buf(\uc8051golden_1.n0132 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0132 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0132 [5], 1'b0);
  buf(\uc8051golden_1.n0132 [6], 1'b0);
  buf(\uc8051golden_1.n0132 [7], 1'b0);
  buf(\uc8051golden_1.n0136 [0], 1'b1);
  buf(\uc8051golden_1.n0136 [1], 1'b0);
  buf(\uc8051golden_1.n0136 [2], 1'b1);
  buf(\uc8051golden_1.n0136 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0136 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0136 [5], 1'b0);
  buf(\uc8051golden_1.n0136 [6], 1'b0);
  buf(\uc8051golden_1.n0136 [7], 1'b0);
  buf(\uc8051golden_1.n0139 , \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0140 , \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0141 [0], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0141 [1], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0141 [2], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0142 , \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n0143 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0143 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0144 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0144 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0144 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n0144 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0144 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0144 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0144 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0144 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0146 [0], 1'b0);
  buf(\uc8051golden_1.n0146 [1], 1'b1);
  buf(\uc8051golden_1.n0146 [2], 1'b1);
  buf(\uc8051golden_1.n0146 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0146 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0146 [5], 1'b0);
  buf(\uc8051golden_1.n0146 [6], 1'b0);
  buf(\uc8051golden_1.n0146 [7], 1'b0);
  buf(\uc8051golden_1.n0150 [0], 1'b1);
  buf(\uc8051golden_1.n0150 [1], 1'b1);
  buf(\uc8051golden_1.n0150 [2], 1'b1);
  buf(\uc8051golden_1.n0150 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0150 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0150 [5], 1'b0);
  buf(\uc8051golden_1.n0150 [6], 1'b0);
  buf(\uc8051golden_1.n0150 [7], 1'b0);
  buf(\uc8051golden_1.n0223 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0223 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0223 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0223 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0223 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0223 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0223 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0223 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0223 [8], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0224 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0224 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0224 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0224 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0224 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0224 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0224 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0224 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0224 [8], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0225 [0], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0225 [1], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0225 [2], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0225 [3], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0225 [4], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0225 [5], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0225 [6], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0225 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0226 , \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0227 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0227 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0227 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n0227 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0227 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0227 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0227 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0227 [7], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0266 [0], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0266 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0266 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0266 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0266 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0266 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0266 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0266 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0268 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0268 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0268 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0268 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0268 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0268 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0268 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0268 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0268 [8], 1'b0);
  buf(\uc8051golden_1.n0274 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0274 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0274 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0274 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0275 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0275 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0275 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0275 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0275 [4], 1'b0);
  buf(\uc8051golden_1.n0282 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0282 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0282 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0282 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0282 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0282 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0282 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0282 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0282 [8], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0291 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0291 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0291 [2], \uc8051golden_1.PSW_24 [2]);
  buf(\uc8051golden_1.n0291 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0291 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0291 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0291 [6], \uc8051golden_1.PSW_24 [6]);
  buf(\uc8051golden_1.n0291 [7], \uc8051golden_1.PSW_24 [7]);
  buf(\uc8051golden_1.n0359 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0359 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0359 [2], \uc8051golden_1.PSW_25 [2]);
  buf(\uc8051golden_1.n0359 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0359 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0359 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0359 [6], \uc8051golden_1.PSW_25 [6]);
  buf(\uc8051golden_1.n0359 [7], \uc8051golden_1.PSW_25 [7]);
  buf(\uc8051golden_1.n0361 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.n0361 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.n0361 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.n0361 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.n0361 [4], \uc8051golden_1.ACC_c6 [4]);
  buf(\uc8051golden_1.n0361 [5], \uc8051golden_1.ACC_c6 [5]);
  buf(\uc8051golden_1.n0361 [6], \uc8051golden_1.ACC_c6 [6]);
  buf(\uc8051golden_1.n0361 [7], \uc8051golden_1.ACC_c6 [7]);
  buf(\uc8051golden_1.n0361 [8], 1'b0);
  buf(\uc8051golden_1.n0365 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.n0365 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.n0365 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.n0365 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.n0366 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.n0366 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.n0366 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.n0366 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.n0366 [4], 1'b0);
  buf(\uc8051golden_1.n0370 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.n0370 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.n0370 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.n0370 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.n0370 [4], \uc8051golden_1.ACC_c6 [4]);
  buf(\uc8051golden_1.n0370 [5], \uc8051golden_1.ACC_c6 [5]);
  buf(\uc8051golden_1.n0370 [6], \uc8051golden_1.ACC_c6 [6]);
  buf(\uc8051golden_1.n0370 [7], \uc8051golden_1.ACC_c6 [7]);
  buf(\uc8051golden_1.n0370 [8], \uc8051golden_1.ACC_c6 [7]);
  buf(\uc8051golden_1.n0378 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0378 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0378 [2], \uc8051golden_1.PSW_26 [2]);
  buf(\uc8051golden_1.n0378 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0378 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0378 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0378 [6], \uc8051golden_1.PSW_26 [6]);
  buf(\uc8051golden_1.n0378 [7], \uc8051golden_1.PSW_26 [7]);
  buf(\uc8051golden_1.n0380 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.n0380 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.n0380 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.n0380 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.n0380 [4], \uc8051golden_1.ACC_c7 [4]);
  buf(\uc8051golden_1.n0380 [5], \uc8051golden_1.ACC_c7 [5]);
  buf(\uc8051golden_1.n0380 [6], \uc8051golden_1.ACC_c7 [6]);
  buf(\uc8051golden_1.n0380 [7], \uc8051golden_1.ACC_c7 [7]);
  buf(\uc8051golden_1.n0380 [8], 1'b0);
  buf(\uc8051golden_1.n0385 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.n0385 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.n0385 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.n0385 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.n0386 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.n0386 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.n0386 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.n0386 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.n0386 [4], 1'b0);
  buf(\uc8051golden_1.n0390 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.n0390 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.n0390 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.n0390 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.n0390 [4], \uc8051golden_1.ACC_c7 [4]);
  buf(\uc8051golden_1.n0390 [5], \uc8051golden_1.ACC_c7 [5]);
  buf(\uc8051golden_1.n0390 [6], \uc8051golden_1.ACC_c7 [6]);
  buf(\uc8051golden_1.n0390 [7], \uc8051golden_1.ACC_c7 [7]);
  buf(\uc8051golden_1.n0390 [8], \uc8051golden_1.ACC_c7 [7]);
  buf(\uc8051golden_1.n0398 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0398 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0398 [2], \uc8051golden_1.PSW_27 [2]);
  buf(\uc8051golden_1.n0398 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0398 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0398 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0398 [6], \uc8051golden_1.PSW_27 [6]);
  buf(\uc8051golden_1.n0398 [7], \uc8051golden_1.PSW_27 [7]);
  buf(\uc8051golden_1.n0417 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0417 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0417 [2], \uc8051golden_1.PSW_28 [2]);
  buf(\uc8051golden_1.n0417 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0417 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0417 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0417 [6], \uc8051golden_1.PSW_28 [6]);
  buf(\uc8051golden_1.n0417 [7], \uc8051golden_1.PSW_28 [7]);
  buf(\uc8051golden_1.n0436 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0436 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0436 [2], \uc8051golden_1.PSW_29 [2]);
  buf(\uc8051golden_1.n0436 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0436 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0436 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0436 [6], \uc8051golden_1.PSW_29 [6]);
  buf(\uc8051golden_1.n0436 [7], \uc8051golden_1.PSW_29 [7]);
  buf(\uc8051golden_1.n0455 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0455 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0455 [2], \uc8051golden_1.PSW_2a [2]);
  buf(\uc8051golden_1.n0455 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0455 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0455 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0455 [6], \uc8051golden_1.PSW_2a [6]);
  buf(\uc8051golden_1.n0455 [7], \uc8051golden_1.PSW_2a [7]);
  buf(\uc8051golden_1.n0474 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0474 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0474 [2], \uc8051golden_1.PSW_2b [2]);
  buf(\uc8051golden_1.n0474 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0474 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0474 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0474 [6], \uc8051golden_1.PSW_2b [6]);
  buf(\uc8051golden_1.n0474 [7], \uc8051golden_1.PSW_2b [7]);
  buf(\uc8051golden_1.n0493 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0493 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0493 [2], \uc8051golden_1.PSW_2c [2]);
  buf(\uc8051golden_1.n0493 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0493 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0493 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0493 [6], \uc8051golden_1.PSW_2c [6]);
  buf(\uc8051golden_1.n0493 [7], \uc8051golden_1.PSW_2c [7]);
  buf(\uc8051golden_1.n0513 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0513 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0513 [2], \uc8051golden_1.PSW_2d [2]);
  buf(\uc8051golden_1.n0513 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0513 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0513 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0513 [6], \uc8051golden_1.PSW_2d [6]);
  buf(\uc8051golden_1.n0513 [7], \uc8051golden_1.PSW_2d [7]);
  buf(\uc8051golden_1.n0532 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0532 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0532 [2], \uc8051golden_1.PSW_2e [2]);
  buf(\uc8051golden_1.n0532 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0532 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0532 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0532 [6], \uc8051golden_1.PSW_2e [6]);
  buf(\uc8051golden_1.n0532 [7], \uc8051golden_1.PSW_2e [7]);
  buf(\uc8051golden_1.n0551 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0551 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0551 [2], \uc8051golden_1.PSW_2f [2]);
  buf(\uc8051golden_1.n0551 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0551 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0551 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0551 [6], \uc8051golden_1.PSW_2f [6]);
  buf(\uc8051golden_1.n0551 [7], \uc8051golden_1.PSW_2f [7]);
  buf(\uc8051golden_1.n0555 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0555 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0555 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0555 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0555 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0555 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0555 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0555 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0555 [8], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0556 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0556 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0556 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0556 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0556 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0556 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0556 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0556 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0556 [8], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0557 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0557 [1], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0557 [2], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0557 [3], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0557 [4], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0557 [5], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0557 [6], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0557 [7], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0558 , \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0559 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0559 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0559 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n0559 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0559 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0559 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0559 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0559 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0560 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0560 [1], 1'b0);
  buf(\uc8051golden_1.n0560 [2], 1'b0);
  buf(\uc8051golden_1.n0560 [3], 1'b0);
  buf(\uc8051golden_1.n0560 [4], 1'b0);
  buf(\uc8051golden_1.n0560 [5], 1'b0);
  buf(\uc8051golden_1.n0560 [6], 1'b0);
  buf(\uc8051golden_1.n0560 [7], 1'b0);
  buf(\uc8051golden_1.n0563 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0563 [1], 1'b0);
  buf(\uc8051golden_1.n0563 [2], 1'b0);
  buf(\uc8051golden_1.n0563 [3], 1'b0);
  buf(\uc8051golden_1.n0563 [4], 1'b0);
  buf(\uc8051golden_1.n0563 [5], 1'b0);
  buf(\uc8051golden_1.n0563 [6], 1'b0);
  buf(\uc8051golden_1.n0563 [7], 1'b0);
  buf(\uc8051golden_1.n0563 [8], 1'b0);
  buf(\uc8051golden_1.n0567 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n0567 [1], 1'b0);
  buf(\uc8051golden_1.n0567 [2], 1'b0);
  buf(\uc8051golden_1.n0567 [3], 1'b0);
  buf(\uc8051golden_1.n0567 [4], 1'b0);
  buf(\uc8051golden_1.n0578 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0578 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0578 [2], \uc8051golden_1.PSW_34 [2]);
  buf(\uc8051golden_1.n0578 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0578 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0578 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0578 [6], \uc8051golden_1.PSW_34 [6]);
  buf(\uc8051golden_1.n0578 [7], \uc8051golden_1.PSW_34 [7]);
  buf(\uc8051golden_1.n0594 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0594 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0594 [2], \uc8051golden_1.PSW_35 [2]);
  buf(\uc8051golden_1.n0594 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0594 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0594 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0594 [6], \uc8051golden_1.PSW_35 [6]);
  buf(\uc8051golden_1.n0594 [7], \uc8051golden_1.PSW_35 [7]);
  buf(\uc8051golden_1.n0610 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0610 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0610 [2], \uc8051golden_1.PSW_36 [2]);
  buf(\uc8051golden_1.n0610 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0610 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0610 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0610 [6], \uc8051golden_1.PSW_36 [6]);
  buf(\uc8051golden_1.n0610 [7], \uc8051golden_1.PSW_36 [7]);
  buf(\uc8051golden_1.n0626 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0626 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0626 [2], \uc8051golden_1.PSW_37 [2]);
  buf(\uc8051golden_1.n0626 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0626 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0626 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0626 [6], \uc8051golden_1.PSW_37 [6]);
  buf(\uc8051golden_1.n0626 [7], \uc8051golden_1.PSW_37 [7]);
  buf(\uc8051golden_1.n0642 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0642 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0642 [2], \uc8051golden_1.PSW_38 [2]);
  buf(\uc8051golden_1.n0642 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0642 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0642 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0642 [6], \uc8051golden_1.PSW_38 [6]);
  buf(\uc8051golden_1.n0642 [7], \uc8051golden_1.PSW_38 [7]);
  buf(\uc8051golden_1.n0658 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0658 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0658 [2], \uc8051golden_1.PSW_39 [2]);
  buf(\uc8051golden_1.n0658 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0658 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0658 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0658 [6], \uc8051golden_1.PSW_39 [6]);
  buf(\uc8051golden_1.n0658 [7], \uc8051golden_1.PSW_39 [7]);
  buf(\uc8051golden_1.n0674 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0674 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0674 [2], \uc8051golden_1.PSW_3a [2]);
  buf(\uc8051golden_1.n0674 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0674 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0674 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0674 [6], \uc8051golden_1.PSW_3a [6]);
  buf(\uc8051golden_1.n0674 [7], \uc8051golden_1.PSW_3a [7]);
  buf(\uc8051golden_1.n0690 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0690 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0690 [2], \uc8051golden_1.PSW_3b [2]);
  buf(\uc8051golden_1.n0690 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0690 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0690 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0690 [6], \uc8051golden_1.PSW_3b [6]);
  buf(\uc8051golden_1.n0690 [7], \uc8051golden_1.PSW_3b [7]);
  buf(\uc8051golden_1.n0706 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0706 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0706 [2], \uc8051golden_1.PSW_3c [2]);
  buf(\uc8051golden_1.n0706 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0706 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0706 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0706 [6], \uc8051golden_1.PSW_3c [6]);
  buf(\uc8051golden_1.n0706 [7], \uc8051golden_1.PSW_3c [7]);
  buf(\uc8051golden_1.n0722 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0722 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0722 [2], \uc8051golden_1.PSW_3d [2]);
  buf(\uc8051golden_1.n0722 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0722 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0722 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0722 [6], \uc8051golden_1.PSW_3d [6]);
  buf(\uc8051golden_1.n0722 [7], \uc8051golden_1.PSW_3d [7]);
  buf(\uc8051golden_1.n0738 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0738 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0738 [2], \uc8051golden_1.PSW_3e [2]);
  buf(\uc8051golden_1.n0738 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0738 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0738 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0738 [6], \uc8051golden_1.PSW_3e [6]);
  buf(\uc8051golden_1.n0738 [7], \uc8051golden_1.PSW_3e [7]);
  buf(\uc8051golden_1.n0754 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0754 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0754 [2], \uc8051golden_1.PSW_3f [2]);
  buf(\uc8051golden_1.n0754 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0754 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0754 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0754 [6], \uc8051golden_1.PSW_3f [6]);
  buf(\uc8051golden_1.n0754 [7], \uc8051golden_1.PSW_3f [7]);
  buf(\uc8051golden_1.n0934 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0934 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0934 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n0934 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0934 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0934 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0934 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0935 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0935 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0935 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n0935 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0935 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0935 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0935 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0935 [7], \uc8051golden_1.PSW_72 [7]);
  buf(\uc8051golden_1.n0936 [0], \uc8051golden_1.DPL [0]);
  buf(\uc8051golden_1.n0936 [1], \uc8051golden_1.DPL [1]);
  buf(\uc8051golden_1.n0936 [2], \uc8051golden_1.DPL [2]);
  buf(\uc8051golden_1.n0936 [3], \uc8051golden_1.DPL [3]);
  buf(\uc8051golden_1.n0936 [4], \uc8051golden_1.DPL [4]);
  buf(\uc8051golden_1.n0936 [5], \uc8051golden_1.DPL [5]);
  buf(\uc8051golden_1.n0936 [6], \uc8051golden_1.DPL [6]);
  buf(\uc8051golden_1.n0936 [7], \uc8051golden_1.DPL [7]);
  buf(\uc8051golden_1.n0936 [8], \uc8051golden_1.DPH [0]);
  buf(\uc8051golden_1.n0936 [9], \uc8051golden_1.DPH [1]);
  buf(\uc8051golden_1.n0936 [10], \uc8051golden_1.DPH [2]);
  buf(\uc8051golden_1.n0936 [11], \uc8051golden_1.DPH [3]);
  buf(\uc8051golden_1.n0936 [12], \uc8051golden_1.DPH [4]);
  buf(\uc8051golden_1.n0936 [13], \uc8051golden_1.DPH [5]);
  buf(\uc8051golden_1.n0936 [14], \uc8051golden_1.DPH [6]);
  buf(\uc8051golden_1.n0936 [15], \uc8051golden_1.DPH [7]);
  buf(\uc8051golden_1.n0937 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n0937 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n0937 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n0937 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n0937 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n0937 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n0937 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n0937 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n0937 [8], 1'b0);
  buf(\uc8051golden_1.n0937 [9], 1'b0);
  buf(\uc8051golden_1.n0937 [10], 1'b0);
  buf(\uc8051golden_1.n0937 [11], 1'b0);
  buf(\uc8051golden_1.n0937 [12], 1'b0);
  buf(\uc8051golden_1.n0937 [13], 1'b0);
  buf(\uc8051golden_1.n0937 [14], 1'b0);
  buf(\uc8051golden_1.n0937 [15], 1'b0);
  buf(\uc8051golden_1.n0962 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0962 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0962 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n0962 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0962 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0962 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0962 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0962 [7], \uc8051golden_1.PSW_82 [7]);
  buf(\uc8051golden_1.n0971 [0], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0971 [1], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0971 [2], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0971 [3], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0973 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n0973 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n0973 [2], \uc8051golden_1.PSW_84 [2]);
  buf(\uc8051golden_1.n0973 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n0973 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n0973 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n0973 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n0973 [7], 1'b0);
  buf(\uc8051golden_1.n1207 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1207 [1], 1'b0);
  buf(\uc8051golden_1.n1207 [2], 1'b0);
  buf(\uc8051golden_1.n1207 [3], 1'b0);
  buf(\uc8051golden_1.n1207 [4], 1'b0);
  buf(\uc8051golden_1.n1207 [5], 1'b0);
  buf(\uc8051golden_1.n1207 [6], 1'b0);
  buf(\uc8051golden_1.n1207 [7], 1'b0);
  buf(\uc8051golden_1.n1223 [0], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1223 [1], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1223 [2], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1223 [3], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1223 [4], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1223 [5], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1223 [6], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1223 [7], \uc8051golden_1.PSW [7]);
  buf(\uc8051golden_1.n1235 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1235 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1235 [2], \uc8051golden_1.PSW_94 [2]);
  buf(\uc8051golden_1.n1235 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1235 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1235 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1235 [6], \uc8051golden_1.PSW_94 [6]);
  buf(\uc8051golden_1.n1235 [7], \uc8051golden_1.PSW_94 [7]);
  buf(\uc8051golden_1.n1248 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1248 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1248 [2], \uc8051golden_1.PSW_95 [2]);
  buf(\uc8051golden_1.n1248 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1248 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1248 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1248 [6], \uc8051golden_1.PSW_95 [6]);
  buf(\uc8051golden_1.n1248 [7], \uc8051golden_1.PSW_95 [7]);
  buf(\uc8051golden_1.n1261 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1261 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1261 [2], \uc8051golden_1.PSW_96 [2]);
  buf(\uc8051golden_1.n1261 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1261 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1261 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1261 [6], \uc8051golden_1.PSW_96 [6]);
  buf(\uc8051golden_1.n1261 [7], \uc8051golden_1.PSW_96 [7]);
  buf(\uc8051golden_1.n1274 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1274 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1274 [2], \uc8051golden_1.PSW_97 [2]);
  buf(\uc8051golden_1.n1274 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1274 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1274 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1274 [6], \uc8051golden_1.PSW_97 [6]);
  buf(\uc8051golden_1.n1274 [7], \uc8051golden_1.PSW_97 [7]);
  buf(\uc8051golden_1.n1287 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1287 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1287 [2], \uc8051golden_1.PSW_98 [2]);
  buf(\uc8051golden_1.n1287 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1287 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1287 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1287 [6], \uc8051golden_1.PSW_98 [6]);
  buf(\uc8051golden_1.n1287 [7], \uc8051golden_1.PSW_98 [7]);
  buf(\uc8051golden_1.n1300 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1300 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1300 [2], \uc8051golden_1.PSW_99 [2]);
  buf(\uc8051golden_1.n1300 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1300 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1300 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1300 [6], \uc8051golden_1.PSW_99 [6]);
  buf(\uc8051golden_1.n1300 [7], \uc8051golden_1.PSW_99 [7]);
  buf(\uc8051golden_1.n1313 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1313 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1313 [2], \uc8051golden_1.PSW_9a [2]);
  buf(\uc8051golden_1.n1313 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1313 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1313 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1313 [6], \uc8051golden_1.PSW_9a [6]);
  buf(\uc8051golden_1.n1313 [7], \uc8051golden_1.PSW_9a [7]);
  buf(\uc8051golden_1.n1326 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1326 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1326 [2], \uc8051golden_1.PSW_9b [2]);
  buf(\uc8051golden_1.n1326 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1326 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1326 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1326 [6], \uc8051golden_1.PSW_9b [6]);
  buf(\uc8051golden_1.n1326 [7], \uc8051golden_1.PSW_9b [7]);
  buf(\uc8051golden_1.n1339 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1339 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1339 [2], \uc8051golden_1.PSW_9c [2]);
  buf(\uc8051golden_1.n1339 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1339 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1339 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1339 [6], \uc8051golden_1.PSW_9c [6]);
  buf(\uc8051golden_1.n1339 [7], \uc8051golden_1.PSW_9c [7]);
  buf(\uc8051golden_1.n1352 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1352 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1352 [2], \uc8051golden_1.PSW_9d [2]);
  buf(\uc8051golden_1.n1352 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1352 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1352 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1352 [6], \uc8051golden_1.PSW_9d [6]);
  buf(\uc8051golden_1.n1352 [7], \uc8051golden_1.PSW_9d [7]);
  buf(\uc8051golden_1.n1365 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1365 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1365 [2], \uc8051golden_1.PSW_9e [2]);
  buf(\uc8051golden_1.n1365 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1365 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1365 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1365 [6], \uc8051golden_1.PSW_9e [6]);
  buf(\uc8051golden_1.n1365 [7], \uc8051golden_1.PSW_9e [7]);
  buf(\uc8051golden_1.n1378 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1378 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1378 [2], \uc8051golden_1.PSW_9f [2]);
  buf(\uc8051golden_1.n1378 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1378 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1378 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1378 [6], \uc8051golden_1.PSW_9f [6]);
  buf(\uc8051golden_1.n1378 [7], \uc8051golden_1.PSW_9f [7]);
  buf(\uc8051golden_1.n1381 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1381 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1381 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1381 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1381 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1381 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1381 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1381 [7], \uc8051golden_1.PSW_a0 [7]);
  buf(\uc8051golden_1.n1382 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1382 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1382 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1382 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1382 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1382 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1382 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1382 [7], \uc8051golden_1.PSW_a2 [7]);
  buf(\uc8051golden_1.n1386 [0], \uc8051golden_1.B [0]);
  buf(\uc8051golden_1.n1386 [1], \uc8051golden_1.B [1]);
  buf(\uc8051golden_1.n1386 [2], \uc8051golden_1.B [2]);
  buf(\uc8051golden_1.n1386 [3], \uc8051golden_1.B [3]);
  buf(\uc8051golden_1.n1386 [4], \uc8051golden_1.B [4]);
  buf(\uc8051golden_1.n1386 [5], \uc8051golden_1.B [5]);
  buf(\uc8051golden_1.n1386 [6], \uc8051golden_1.B [6]);
  buf(\uc8051golden_1.n1386 [7], \uc8051golden_1.B [7]);
  buf(\uc8051golden_1.n1386 [8], 1'b0);
  buf(\uc8051golden_1.n1386 [9], 1'b0);
  buf(\uc8051golden_1.n1386 [10], 1'b0);
  buf(\uc8051golden_1.n1386 [11], 1'b0);
  buf(\uc8051golden_1.n1386 [12], 1'b0);
  buf(\uc8051golden_1.n1386 [13], 1'b0);
  buf(\uc8051golden_1.n1386 [14], 1'b0);
  buf(\uc8051golden_1.n1386 [15], 1'b0);
  buf(\uc8051golden_1.n1393 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1393 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1393 [2], \uc8051golden_1.PSW_a4 [2]);
  buf(\uc8051golden_1.n1393 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1393 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1393 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1393 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1393 [7], 1'b0);
  buf(\uc8051golden_1.n1395 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1395 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1395 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1395 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1395 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1395 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1395 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1395 [7], \uc8051golden_1.PSW_b0 [7]);
  buf(\uc8051golden_1.n1411 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1411 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1411 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1411 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1411 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1411 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1411 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1411 [7], \uc8051golden_1.PSW_b3 [7]);
  buf(\uc8051golden_1.n1417 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1417 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1417 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1417 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1417 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1417 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1417 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1417 [7], \uc8051golden_1.PSW_b4 [7]);
  buf(\uc8051golden_1.n1423 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1423 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1423 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1423 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1423 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1423 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1423 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1423 [7], \uc8051golden_1.PSW_b5 [7]);
  buf(\uc8051golden_1.n1429 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1429 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1429 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1429 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1429 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1429 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1429 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1429 [7], \uc8051golden_1.PSW_b6 [7]);
  buf(\uc8051golden_1.n1436 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1436 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1436 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1436 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1436 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1436 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1436 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1436 [7], \uc8051golden_1.PSW_b7 [7]);
  buf(\uc8051golden_1.n1442 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1442 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1442 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1442 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1442 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1442 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1442 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1442 [7], \uc8051golden_1.PSW_b8 [7]);
  buf(\uc8051golden_1.n1448 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1448 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1448 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1448 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1448 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1448 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1448 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1448 [7], \uc8051golden_1.PSW_b9 [7]);
  buf(\uc8051golden_1.n1454 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1454 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1454 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1454 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1454 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1454 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1454 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1454 [7], \uc8051golden_1.PSW_ba [7]);
  buf(\uc8051golden_1.n1460 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1460 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1460 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1460 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1460 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1460 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1460 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1460 [7], \uc8051golden_1.PSW_bb [7]);
  buf(\uc8051golden_1.n1466 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1466 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1466 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1466 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1466 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1466 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1466 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1466 [7], \uc8051golden_1.PSW_bc [7]);
  buf(\uc8051golden_1.n1473 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1473 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1473 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1473 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1473 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1473 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1473 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1473 [7], \uc8051golden_1.PSW_bd [7]);
  buf(\uc8051golden_1.n1479 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1479 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1479 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1479 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1479 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1479 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1479 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1479 [7], \uc8051golden_1.PSW_be [7]);
  buf(\uc8051golden_1.n1485 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1485 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1485 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1485 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1485 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1485 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1485 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1485 [7], \uc8051golden_1.PSW_bf [7]);
  buf(\uc8051golden_1.n1486 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1486 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1486 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1486 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1486 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1486 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1486 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1486 [7], 1'b0);
  buf(\uc8051golden_1.n1487 [0], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1487 [1], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1487 [2], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1487 [3], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1488 [0], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1488 [1], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1488 [2], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1488 [3], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1488 [4], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1488 [5], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1488 [6], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1488 [7], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1544 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1544 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1544 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1544 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1544 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1544 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1544 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1544 [7], 1'b1);
  buf(\uc8051golden_1.n1564 [0], \uc8051golden_1.PSW [0]);
  buf(\uc8051golden_1.n1564 [1], \uc8051golden_1.PSW [1]);
  buf(\uc8051golden_1.n1564 [2], \uc8051golden_1.PSW [2]);
  buf(\uc8051golden_1.n1564 [3], \uc8051golden_1.PSW [3]);
  buf(\uc8051golden_1.n1564 [4], \uc8051golden_1.PSW [4]);
  buf(\uc8051golden_1.n1564 [5], \uc8051golden_1.PSW [5]);
  buf(\uc8051golden_1.n1564 [6], \uc8051golden_1.PSW [6]);
  buf(\uc8051golden_1.n1564 [7], \uc8051golden_1.PSW_d4 [7]);
  buf(\uc8051golden_1.n1568 [0], \uc8051golden_1.ACC_c6 [0]);
  buf(\uc8051golden_1.n1568 [1], \uc8051golden_1.ACC_c6 [1]);
  buf(\uc8051golden_1.n1568 [2], \uc8051golden_1.ACC_c6 [2]);
  buf(\uc8051golden_1.n1568 [3], \uc8051golden_1.ACC_c6 [3]);
  buf(\uc8051golden_1.n1568 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1568 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1568 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1568 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1569 [0], \uc8051golden_1.ACC_c6 [4]);
  buf(\uc8051golden_1.n1569 [1], \uc8051golden_1.ACC_c6 [5]);
  buf(\uc8051golden_1.n1569 [2], \uc8051golden_1.ACC_c6 [6]);
  buf(\uc8051golden_1.n1569 [3], \uc8051golden_1.ACC_c6 [7]);
  buf(\uc8051golden_1.n1570 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1570 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1570 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1570 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1570 [4], \uc8051golden_1.ACC_c6 [4]);
  buf(\uc8051golden_1.n1570 [5], \uc8051golden_1.ACC_c6 [5]);
  buf(\uc8051golden_1.n1570 [6], \uc8051golden_1.ACC_c6 [6]);
  buf(\uc8051golden_1.n1570 [7], \uc8051golden_1.ACC_c6 [7]);
  buf(\uc8051golden_1.n1571 [0], \uc8051golden_1.ACC_c7 [0]);
  buf(\uc8051golden_1.n1571 [1], \uc8051golden_1.ACC_c7 [1]);
  buf(\uc8051golden_1.n1571 [2], \uc8051golden_1.ACC_c7 [2]);
  buf(\uc8051golden_1.n1571 [3], \uc8051golden_1.ACC_c7 [3]);
  buf(\uc8051golden_1.n1571 [4], \uc8051golden_1.ACC [4]);
  buf(\uc8051golden_1.n1571 [5], \uc8051golden_1.ACC [5]);
  buf(\uc8051golden_1.n1571 [6], \uc8051golden_1.ACC [6]);
  buf(\uc8051golden_1.n1571 [7], \uc8051golden_1.ACC [7]);
  buf(\uc8051golden_1.n1572 [0], \uc8051golden_1.ACC_c7 [4]);
  buf(\uc8051golden_1.n1572 [1], \uc8051golden_1.ACC_c7 [5]);
  buf(\uc8051golden_1.n1572 [2], \uc8051golden_1.ACC_c7 [6]);
  buf(\uc8051golden_1.n1572 [3], \uc8051golden_1.ACC_c7 [7]);
  buf(\uc8051golden_1.n1573 [0], \uc8051golden_1.ACC [0]);
  buf(\uc8051golden_1.n1573 [1], \uc8051golden_1.ACC [1]);
  buf(\uc8051golden_1.n1573 [2], \uc8051golden_1.ACC [2]);
  buf(\uc8051golden_1.n1573 [3], \uc8051golden_1.ACC [3]);
  buf(\uc8051golden_1.n1573 [4], \uc8051golden_1.ACC_c7 [4]);
  buf(\uc8051golden_1.n1573 [5], \uc8051golden_1.ACC_c7 [5]);
  buf(\uc8051golden_1.n1573 [6], \uc8051golden_1.ACC_c7 [6]);
  buf(\uc8051golden_1.n1573 [7], \uc8051golden_1.ACC_c7 [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
