
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire [15:0] _31420_;
  wire [15:0] _31421_;
  wire [15:0] _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire [7:0] _33298_;
  wire [3:0] _33299_;
  wire [1:0] _33300_;
  wire [7:0] _33301_;
  wire [3:0] _33302_;
  wire [1:0] _33303_;
  wire [7:0] _33304_;
  wire [3:0] _33305_;
  wire [1:0] _33306_;
  wire [15:0] _33307_;
  wire [15:0] _33308_;
  wire [15:0] _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire [15:0] _33476_;
  wire [15:0] _33477_;
  wire [15:0] _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire [3:0] _33493_;
  wire [7:0] _33494_;
  wire [7:0] _33495_;
  wire [3:0] _33496_;
  wire [7:0] _33497_;
  wire [7:0] _33498_;
  wire [3:0] _33499_;
  wire [7:0] _33500_;
  wire [7:0] _33501_;
  wire [3:0] _33502_;
  wire [7:0] _33503_;
  wire [7:0] _33504_;
  wire [15:0] _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire [1:0] _33638_;
  wire [1:0] _33639_;
  wire [1:0] _33640_;
  wire [1:0] _33641_;
  wire [1:0] _33642_;
  wire [1:0] _33643_;
  wire [1:0] _33644_;
  wire [1:0] _33645_;
  wire [1:0] _33646_;
  wire [1:0] _33647_;
  wire [1:0] _33648_;
  wire [1:0] _33649_;
  wire [1:0] _33650_;
  wire [1:0] _33651_;
  wire [1:0] _33652_;
  wire [1:0] _33653_;
  wire [1:0] _33654_;
  wire [1:0] _33655_;
  wire [1:0] _33656_;
  wire [1:0] _33657_;
  wire [1:0] _33658_;
  wire [1:0] _33659_;
  wire [6:0] _33660_;
  wire [3:0] _33661_;
  wire [1:0] _33662_;
  wire [6:0] _33663_;
  wire [3:0] _33664_;
  wire [1:0] _33665_;
  wire [6:0] _33666_;
  wire [3:0] _33667_;
  wire [1:0] _33668_;
  wire [6:0] _33669_;
  wire [3:0] _33670_;
  wire [1:0] _33671_;
  wire [3:0] _33672_;
  wire [3:0] _33673_;
  wire [3:0] _33674_;
  wire [3:0] _33675_;
  wire [3:0] _33676_;
  wire [3:0] _33677_;
  wire [3:0] _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire [7:0] _33759_;
  wire [7:0] _33760_;
  wire [7:0] _33761_;
  wire [7:0] _33762_;
  wire [7:0] _33763_;
  wire [7:0] _33764_;
  wire [7:0] _33765_;
  wire [7:0] _33766_;
  wire [7:0] _33767_;
  wire [7:0] _33768_;
  wire [7:0] _33769_;
  wire [7:0] _33770_;
  wire [7:0] _33771_;
  wire [7:0] _33772_;
  wire [7:0] _33773_;
  wire [7:0] _33774_;
  wire [7:0] _33775_;
  wire [7:0] _33776_;
  wire [7:0] _33777_;
  wire [7:0] _33778_;
  wire [7:0] _33779_;
  wire [7:0] _33780_;
  wire [7:0] _33781_;
  wire [7:0] _33782_;
  wire [7:0] _33783_;
  wire [7:0] _33784_;
  wire [7:0] _33785_;
  wire [7:0] _33786_;
  wire [7:0] _33787_;
  wire [7:0] _33788_;
  wire [7:0] _33789_;
  wire [7:0] _33790_;
  wire [7:0] _33791_;
  wire [7:0] _33792_;
  wire [7:0] _33793_;
  wire [7:0] _33794_;
  wire [7:0] _33795_;
  wire [7:0] _33796_;
  wire [7:0] _33797_;
  wire [7:0] _33798_;
  wire [7:0] _33799_;
  wire [7:0] _33800_;
  wire [7:0] _33801_;
  wire [7:0] _33802_;
  wire [7:0] _33803_;
  wire [7:0] _33804_;
  wire [7:0] _33805_;
  wire [7:0] _33806_;
  wire [7:0] _33807_;
  wire [7:0] _33808_;
  wire [7:0] _33809_;
  wire [7:0] _33810_;
  wire [7:0] _33811_;
  wire [7:0] _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire [7:0] _33877_;
  wire [7:0] _33878_;
  wire [7:0] _33879_;
  wire [7:0] _33880_;
  wire [7:0] _33881_;
  wire [7:0] _33882_;
  wire [7:0] _33883_;
  wire [7:0] _33884_;
  wire [7:0] _33885_;
  wire [7:0] _33886_;
  wire [7:0] _33887_;
  wire [7:0] _33888_;
  wire [7:0] _33889_;
  wire [7:0] _33890_;
  wire [7:0] _33891_;
  wire [7:0] _33892_;
  wire [7:0] _33893_;
  wire [7:0] _33894_;
  wire [7:0] _33895_;
  wire [7:0] _33896_;
  wire [7:0] _33897_;
  wire [7:0] _33898_;
  wire [7:0] _33899_;
  wire [7:0] _33900_;
  wire [7:0] _33901_;
  wire [7:0] _33902_;
  wire [7:0] _33903_;
  wire [7:0] _33904_;
  wire [7:0] _33905_;
  wire [7:0] _33906_;
  wire [7:0] _33907_;
  wire [7:0] _33908_;
  wire [7:0] _33909_;
  wire [7:0] _33910_;
  wire [7:0] _33911_;
  wire [7:0] _33912_;
  wire [7:0] _33913_;
  wire [7:0] _33914_;
  wire [7:0] _33915_;
  wire [7:0] _33916_;
  wire [7:0] _33917_;
  wire [7:0] _33918_;
  wire [7:0] _33919_;
  wire [7:0] _33920_;
  wire [7:0] _33921_;
  wire [7:0] _33922_;
  wire [7:0] _33923_;
  wire [7:0] _33924_;
  wire [7:0] _33925_;
  wire [7:0] _33926_;
  wire [7:0] _33927_;
  wire [7:0] _33928_;
  wire [7:0] _33929_;
  wire [7:0] _33930_;
  wire [7:0] _33931_;
  wire [7:0] _33932_;
  wire [7:0] _33933_;
  wire [7:0] _33934_;
  wire [7:0] _33935_;
  wire [7:0] _33936_;
  wire [7:0] _33937_;
  wire [7:0] _33938_;
  wire [7:0] _33939_;
  wire [7:0] _33940_;
  wire [7:0] _33941_;
  wire [7:0] _33942_;
  wire [7:0] _33943_;
  wire [7:0] _33944_;
  wire [7:0] _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire [3:0] _34135_;
  wire [7:0] _34136_;
  wire [7:0] _34137_;
  wire [3:0] _34138_;
  wire [7:0] _34139_;
  wire [7:0] _34140_;
  wire [3:0] _34141_;
  wire [7:0] _34142_;
  wire [7:0] _34143_;
  wire [3:0] _34144_;
  wire [7:0] _34145_;
  wire [7:0] _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire [15:0] _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire [15:0] _34155_;
  wire [15:0] _34156_;
  wire [15:0] _34157_;
  wire [15:0] _34158_;
  wire [31:0] _34159_;
  wire [31:0] _34160_;
  wire [31:0] _34161_;
  wire [31:0] _34162_;
  wire [31:0] _34163_;
  wire [31:0] _34164_;
  wire [15:0] _34165_;
  wire [15:0] _34166_;
  wire [15:0] _34167_;
  wire [15:0] _34168_;
  wire [15:0] _34169_;
  wire [15:0] _34170_;
  wire [15:0] _34171_;
  wire [15:0] _34172_;
  wire [15:0] _34173_;
  wire [15:0] _34174_;
  wire [15:0] _34175_;
  wire [15:0] _34176_;
  wire [15:0] _34177_;
  wire [15:0] _34178_;
  wire [15:0] _34179_;
  wire [15:0] _34180_;
  wire [15:0] _34181_;
  wire [15:0] _34182_;
  wire [15:0] _34183_;
  wire [15:0] _34184_;
  wire [15:0] _34185_;
  wire [15:0] _34186_;
  wire [15:0] _34187_;
  wire [15:0] _34188_;
  wire [15:0] _34189_;
  wire [15:0] _34190_;
  wire [15:0] _34191_;
  wire [15:0] _34192_;
  wire [15:0] _34193_;
  wire [15:0] _34194_;
  wire [15:0] _34195_;
  wire [15:0] _34196_;
  wire [15:0] _34197_;
  wire [15:0] _34198_;
  wire [15:0] _34199_;
  wire [15:0] _34200_;
  wire [15:0] _34201_;
  wire [15:0] _34202_;
  wire [15:0] _34203_;
  wire [15:0] _34204_;
  wire [15:0] _34205_;
  wire [15:0] _34206_;
  wire [15:0] _34207_;
  wire [15:0] _34208_;
  wire [15:0] _34209_;
  wire [15:0] _34210_;
  wire [15:0] _34211_;
  wire [15:0] _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire [7:0] _34220_;
  wire [3:0] _34221_;
  wire [7:0] _34222_;
  wire [7:0] _34223_;
  wire [3:0] _34224_;
  wire [7:0] _34225_;
  wire [4:0] _34226_;
  wire [3:0] _34227_;
  wire [1:0] _34228_;
  wire [7:0] _34229_;
  wire [4:0] _34230_;
  wire [4:0] _34231_;
  wire [4:0] _34232_;
  wire [4:0] _34233_;
  wire [7:0] _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire [3:0] _34242_;
  wire [1:0] _34243_;
  wire _34244_;
  wire [5:0] _34245_;
  wire [2:0] _34246_;
  wire [1:0] _34247_;
  wire [1:0] _34248_;
  wire [1:0] _34249_;
  wire [1:0] _34250_;
  wire [1:0] _34251_;
  wire [1:0] _34252_;
  wire [1:0] _34253_;
  wire [6:0] _34254_;
  wire [2:0] _34255_;
  wire [1:0] _34256_;
  wire [6:0] _34257_;
  wire [2:0] _34258_;
  wire [1:0] _34259_;
  wire [6:0] _34260_;
  wire [2:0] _34261_;
  wire [1:0] _34262_;
  wire [6:0] _34263_;
  wire [2:0] _34264_;
  wire [1:0] _34265_;
  wire [6:0] _34266_;
  wire [2:0] _34267_;
  wire [1:0] _34268_;
  wire [6:0] _34269_;
  wire [2:0] _34270_;
  wire [1:0] _34271_;
  wire [6:0] _34272_;
  wire [2:0] _34273_;
  wire [1:0] _34274_;
  wire [6:0] _34275_;
  wire [2:0] _34276_;
  wire [1:0] _34277_;
  wire [6:0] _34278_;
  wire [2:0] _34279_;
  wire [1:0] _34280_;
  wire [6:0] _34281_;
  wire [2:0] _34282_;
  wire [1:0] _34283_;
  wire [2:0] _34284_;
  wire [1:0] _34285_;
  wire [2:0] _34286_;
  wire [1:0] _34287_;
  wire [2:0] _34288_;
  wire [1:0] _34289_;
  wire [2:0] _34290_;
  wire [1:0] _34291_;
  wire [2:0] _34292_;
  wire [1:0] _34293_;
  wire [2:0] _34294_;
  wire [1:0] _34295_;
  wire [2:0] _34296_;
  wire [1:0] _34297_;
  wire [2:0] _34298_;
  wire [1:0] _34299_;
  wire [1:0] _34300_;
  wire [2:0] _34301_;
  wire [1:0] _34302_;
  wire [2:0] _34303_;
  wire [1:0] _34304_;
  wire [2:0] _34305_;
  wire [1:0] _34306_;
  wire [2:0] _34307_;
  wire [1:0] _34308_;
  wire [2:0] _34309_;
  wire [1:0] _34310_;
  wire [2:0] _34311_;
  wire [1:0] _34312_;
  wire [2:0] _34313_;
  wire [1:0] _34314_;
  wire [2:0] _34315_;
  wire [1:0] _34316_;
  wire [2:0] _34317_;
  wire [1:0] _34318_;
  wire [5:0] _34319_;
  wire [2:0] _34320_;
  wire _34321_;
  wire [5:0] _34322_;
  wire [2:0] _34323_;
  wire _34324_;
  wire _34325_;
  wire [1:0] _34326_;
  wire [3:0] _34327_;
  wire [3:0] _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire [7:0] _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire [7:0] _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire [4:0] _34370_;
  wire [4:0] _34371_;
  wire [4:0] _34372_;
  wire [3:0] _34373_;
  wire [1:0] _34374_;
  wire [4:0] _34375_;
  wire [4:0] _34376_;
  wire [3:0] _34377_;
  wire [3:0] _34378_;
  wire [1:0] _34379_;
  wire [15:0] _34380_;
  wire [7:0] _34381_;
  wire [4:0] _34382_;
  wire [4:0] _34383_;
  wire [4:0] _34384_;
  wire [4:0] _34385_;
  wire [3:0] _34386_;
  wire [3:0] _34387_;
  wire [3:0] _34388_;
  wire [3:0] _34389_;
  wire [3:0] _34390_;
  wire [3:0] _34391_;
  wire [3:0] _34392_;
  wire [3:0] _34393_;
  wire [3:0] _34394_;
  wire [3:0] _34395_;
  wire [3:0] _34396_;
  wire [3:0] _34397_;
  wire [3:0] _34398_;
  wire [3:0] _34399_;
  wire [3:0] _34400_;
  wire [3:0] _34401_;
  wire [3:0] _34402_;
  wire [3:0] _34403_;
  wire [3:0] _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire [3:0] _34410_;
  wire [3:0] _34411_;
  wire [3:0] _34412_;
  wire [3:0] _34413_;
  wire [3:0] _34414_;
  wire [3:0] _34415_;
  wire [3:0] _34416_;
  wire [3:0] _34417_;
  wire [3:0] _34418_;
  wire [3:0] _34419_;
  wire [3:0] _34420_;
  wire [3:0] _34421_;
  wire [3:0] _34422_;
  wire [3:0] _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire [7:0] _34438_;
  wire [7:0] _34439_;
  wire [7:0] _34440_;
  wire [7:0] _34441_;
  wire [7:0] _34442_;
  wire [7:0] _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire [4:0] _34475_;
  wire [4:0] _34476_;
  wire [4:0] _34477_;
  wire [4:0] _34478_;
  wire [4:0] _34479_;
  wire [4:0] _34480_;
  wire [3:0] _34481_;
  wire [3:0] _34482_;
  wire [3:0] _34483_;
  wire [3:0] _34484_;
  wire [3:0] _34485_;
  wire [3:0] _34486_;
  wire [1:0] _34487_;
  wire [1:0] _34488_;
  wire [15:0] _34489_;
  wire [15:0] _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire [4:0] _34524_;
  wire [4:0] _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire [4:0] _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire [3:0] _34539_;
  wire [3:0] _34540_;
  wire _34541_;
  wire _34542_;
  wire [3:0] _34543_;
  wire _34544_;
  wire _34545_;
  wire [1:0] _34546_;
  wire [1:0] _34547_;
  wire _34548_;
  wire [1:0] _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire [7:0] _34591_;
  wire _34592_;
  wire [1:0] _34593_;
  wire [1:0] _34594_;
  wire [3:0] _34595_;
  wire [1:0] _34596_;
  wire [3:0] _34597_;
  wire [1:0] _34598_;
  wire [3:0] _34599_;
  wire [1:0] _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire [1:0] _34607_;
  wire [15:0] _34608_;
  wire [1:0] _34609_;
  wire [1:0] _34610_;
  wire [1:0] _34611_;
  wire [8:0] _34612_;
  wire [8:0] _34613_;
  wire [8:0] _34614_;
  wire [8:0] _34615_;
  wire [8:0] _34616_;
  wire [1:0] _34617_;
  wire [8:0] _34618_;
  wire [8:0] _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire [8:0] _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire [1:0] _34661_;
  wire [1:0] _34662_;
  wire [15:0] _34663_;
  wire [15:0] _34664_;
  wire [15:0] _34665_;
  wire [15:0] _34666_;
  wire [15:0] _34667_;
  wire [15:0] _34668_;
  wire [15:0] _34669_;
  wire [15:0] _34670_;
  wire [15:0] _34671_;
  wire [15:0] _34672_;
  wire [15:0] _34673_;
  wire [15:0] _34674_;
  wire [15:0] _34675_;
  wire [15:0] _34676_;
  wire [15:0] _34677_;
  wire [15:0] _34678_;
  wire [15:0] _34679_;
  wire [15:0] _34680_;
  wire [15:0] _34681_;
  wire [15:0] _34682_;
  wire [15:0] _34683_;
  wire [15:0] _34684_;
  wire [3:0] _34685_;
  wire [1:0] _34686_;
  wire [1:0] _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire [15:0] _34691_;
  wire [15:0] _34692_;
  wire [15:0] _34693_;
  wire [15:0] _34694_;
  wire [15:0] _34695_;
  wire [15:0] _34696_;
  wire [15:0] _34697_;
  wire [15:0] _34698_;
  wire [15:0] _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire [15:0] _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire [1:0] _34737_;
  wire [15:0] _34738_;
  wire [15:0] _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire [2:0] _34744_;
  wire [1:0] _34745_;
  wire [2:0] _34746_;
  wire [1:0] _34747_;
  wire [2:0] _34748_;
  wire [1:0] _34749_;
  wire [2:0] _34750_;
  wire [1:0] _34751_;
  wire [2:0] _34752_;
  wire [1:0] _34753_;
  wire [2:0] _34754_;
  wire [1:0] _34755_;
  wire [2:0] _34756_;
  wire [1:0] _34757_;
  wire [2:0] _34758_;
  wire [1:0] _34759_;
  wire [2:0] _34760_;
  wire [1:0] _34761_;
  wire _34762_;
  wire [1:0] _34763_;
  wire [1:0] _34764_;
  wire [2:0] _34765_;
  wire [2:0] _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire [23:0] _34777_;
  wire [7:0] _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire [6:0] _34782_;
  wire [6:0] _34783_;
  wire [6:0] _34784_;
  wire [6:0] _34785_;
  wire [6:0] _34786_;
  wire [6:0] _34787_;
  wire [6:0] _34788_;
  wire [6:0] _34789_;
  wire [7:0] _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire [3:0] _34800_;
  wire [1:0] _34801_;
  wire [3:0] _34802_;
  wire [1:0] _34803_;
  wire _34804_;
  wire _34805_;
  wire [1:0] _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire [1:0] _34823_;
  wire [1:0] _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire [3:0] _34835_;
  wire [1:0] _34836_;
  wire [2:0] _34837_;
  wire [7:0] _34838_;
  wire [1:0] _34839_;
  wire [2:0] _34840_;
  wire [2:0] _34841_;
  wire [1:0] _34842_;
  wire _34843_;
  wire [1:0] _34844_;
  wire _34845_;
  wire [1:0] _34846_;
  wire _34847_;
  wire [1:0] _34848_;
  wire [2:0] _34849_;
  wire _34850_;
  wire [2:0] _34851_;
  wire _34852_;
  wire _34853_;
  wire [1:0] _34854_;
  wire _34855_;
  wire [2:0] _34856_;
  wire [2:0] _34857_;
  wire _34858_;
  wire [2:0] _34859_;
  wire [2:0] _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire [8:0] _34917_;
  wire [4:0] _34918_;
  wire [1:0] _34919_;
  wire _34920_;
  wire [2:0] _34921_;
  wire [1:0] _34922_;
  wire [2:0] _34923_;
  wire _34924_;
  wire [1:0] _34925_;
  wire [3:0] _34926_;
  wire [1:0] _34927_;
  wire _34928_;
  wire [2:0] _34929_;
  wire [1:0] _34930_;
  wire [5:0] _34931_;
  wire [2:0] _34932_;
  wire _34933_;
  wire [4:0] _34934_;
  wire [1:0] _34935_;
  wire _34936_;
  wire _34937_;
  wire [2:0] _34938_;
  wire [1:0] _34939_;
  wire [14:0] _34940_;
  wire [7:0] _34941_;
  wire [3:0] _34942_;
  wire [1:0] _34943_;
  wire [17:0] _34944_;
  wire [8:0] _34945_;
  wire [4:0] _34946_;
  wire [1:0] _34947_;
  wire _34948_;
  wire [1:0] _34949_;
  wire _34950_;
  wire [11:0] _34951_;
  wire [3:0] _34952_;
  wire [1:0] _34953_;
  wire [2:0] _34954_;
  wire _34955_;
  wire [5:0] _34956_;
  wire [2:0] _34957_;
  wire _34958_;
  wire [6:0] _34959_;
  wire [3:0] _34960_;
  wire [1:0] _34961_;
  wire [1:0] _34962_;
  wire _34963_;
  wire [3:0] _34964_;
  wire [1:0] _34965_;
  wire [15:0] _34966_;
  wire [7:0] _34967_;
  wire [3:0] _34968_;
  wire [1:0] _34969_;
  wire _34970_;
  wire [5:0] _34971_;
  wire [2:0] _34972_;
  wire _34973_;
  wire [3:0] _34974_;
  wire [1:0] _34975_;
  wire _34976_;
  wire [1:0] _34977_;
  wire [1:0] _34978_;
  wire [16:0] _34979_;
  wire [7:0] _34980_;
  wire [3:0] _34981_;
  wire [1:0] _34982_;
  wire _34983_;
  wire _34984_;
  wire [5:0] _34985_;
  wire [2:0] _34986_;
  wire [1:0] _34987_;
  wire [8:0] _34988_;
  wire [4:0] _34989_;
  wire [1:0] _34990_;
  wire _34991_;
  wire [1:0] _34992_;
  wire _34993_;
  wire [2:0] _34994_;
  wire [17:0] _34995_;
  wire [8:0] _34996_;
  wire [4:0] _34997_;
  wire [1:0] _34998_;
  wire _34999_;
  wire [5:0] _35000_;
  wire [2:0] _35001_;
  wire _35002_;
  wire [7:0] _35003_;
  wire [3:0] _35004_;
  wire [1:0] _35005_;
  wire _35006_;
  wire [6:0] _35007_;
  wire [2:0] _35008_;
  wire [1:0] _35009_;
  wire [2:0] _35010_;
  wire _35011_;
  wire [10:0] _35012_;
  wire [5:0] _35013_;
  wire [2:0] _35014_;
  wire _35015_;
  wire [3:0] _35016_;
  wire [1:0] _35017_;
  wire [3:0] _35018_;
  wire [1:0] _35019_;
  wire [3:0] _35020_;
  wire [1:0] _35021_;
  wire [3:0] _35022_;
  wire [1:0] _35023_;
  wire [3:0] _35024_;
  wire [1:0] _35025_;
  wire [3:0] _35026_;
  wire [1:0] _35027_;
  wire [3:0] _35028_;
  wire [1:0] _35029_;
  wire [1:0] _35030_;
  wire [1:0] _35031_;
  wire [1:0] _35032_;
  wire [3:0] _35033_;
  wire [1:0] _35034_;
  wire [3:0] _35035_;
  wire [1:0] _35036_;
  wire [1:0] _35037_;
  wire [2:0] _35038_;
  wire [1:0] _35039_;
  wire [2:0] _35040_;
  wire [1:0] _35041_;
  wire [1:0] _35042_;
  wire [3:0] _35043_;
  wire [1:0] _35044_;
  wire [1:0] _35045_;
  wire _35046_;
  wire [1:0] _35047_;
  wire [1:0] _35048_;
  wire [2:0] _35049_;
  wire [1:0] _35050_;
  wire _35051_;
  wire _35052_;
  wire [3:0] _35053_;
  wire [1:0] _35054_;
  wire [3:0] _35055_;
  wire [1:0] _35056_;
  wire [3:0] _35057_;
  wire [1:0] _35058_;
  wire [3:0] _35059_;
  wire [1:0] _35060_;
  wire [3:0] _35061_;
  wire [1:0] _35062_;
  wire [1:0] _35063_;
  wire [3:0] _35064_;
  wire [1:0] _35065_;
  wire [1:0] _35066_;
  wire [1:0] _35067_;
  wire [1:0] _35068_;
  wire [3:0] _35069_;
  wire [1:0] _35070_;
  wire [1:0] _35071_;
  wire [1:0] _35072_;
  wire [1:0] _35073_;
  wire [2:0] _35074_;
  wire [1:0] _35075_;
  wire [1:0] _35076_;
  wire [1:0] _35077_;
  wire _35078_;
  wire [1:0] _35079_;
  wire [1:0] _35080_;
  wire [3:0] _35081_;
  wire [1:0] _35082_;
  wire [1:0] _35083_;
  wire [2:0] _35084_;
  wire [1:0] _35085_;
  wire [2:0] _35086_;
  wire [1:0] _35087_;
  wire [2:0] _35088_;
  wire [1:0] _35089_;
  wire [1:0] _35090_;
  wire [2:0] _35091_;
  wire [1:0] _35092_;
  wire [1:0] _35093_;
  wire [2:0] _35094_;
  wire [1:0] _35095_;
  wire [1:0] _35096_;
  wire [1:0] _35097_;
  wire [1:0] _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire [1:0] _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire [1:0] _35112_;
  wire [1:0] _35113_;
  wire [1:0] _35114_;
  wire [1:0] _35115_;
  wire _35116_;
  wire [6:0] _35117_;
  wire [3:0] _35118_;
  wire [1:0] _35119_;
  wire [6:0] _35120_;
  wire [3:0] _35121_;
  wire [1:0] _35122_;
  wire [6:0] _35123_;
  wire [3:0] _35124_;
  wire [1:0] _35125_;
  wire [6:0] _35126_;
  wire [3:0] _35127_;
  wire [1:0] _35128_;
  wire [3:0] _35129_;
  wire [1:0] _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire [7:0] _35139_;
  wire [7:0] _35140_;
  wire [4:0] _35141_;
  wire [1:0] _35142_;
  wire [7:0] _35143_;
  wire [7:0] _35144_;
  wire [7:0] _35145_;
  wire [7:0] _35146_;
  wire [4:0] _35147_;
  wire [1:0] _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire [2:0] _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire [1:0] _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire [1:0] _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire [1:0] _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire [1:0] _35452_;
  wire [1:0] _35453_;
  wire [1:0] _35454_;
  wire _35455_;
  wire [1:0] _35456_;
  wire [2:0] _35457_;
  wire _35458_;
  wire [2:0] _35459_;
  wire [2:0] _35460_;
  wire [2:0] _35461_;
  wire [2:0] _35462_;
  wire [2:0] _35463_;
  wire [2:0] _35464_;
  wire [1:0] _35465_;
  wire [1:0] _35466_;
  wire [3:0] _35467_;
  wire [3:0] _35468_;
  wire [3:0] _35469_;
  wire [1:0] _35470_;
  wire [1:0] _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire [1:0] _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire [2:0] _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire [2:0] _35501_;
  wire [2:0] _35502_;
  wire [2:0] _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire [2:0] _35520_;
  wire [2:0] _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire [2:0] _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire [1:0] _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire [7:0] _35553_;
  wire [7:0] _35554_;
  wire [7:0] _35555_;
  wire [7:0] _35556_;
  wire [7:0] _35557_;
  wire [7:0] _35558_;
  wire [7:0] _35559_;
  wire [7:0] _35560_;
  wire [7:0] _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire [3:0] _35565_;
  wire [1:0] _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire [1:0] _35571_;
  wire [1:0] _35572_;
  wire [2:0] _35573_;
  wire [1:0] _35574_;
  wire [2:0] _35575_;
  wire [1:0] _35576_;
  wire [2:0] _35577_;
  wire [1:0] _35578_;
  wire [2:0] _35579_;
  wire [1:0] _35580_;
  wire [2:0] _35581_;
  wire [1:0] _35582_;
  wire [2:0] _35583_;
  wire [1:0] _35584_;
  wire [2:0] _35585_;
  wire [1:0] _35586_;
  wire [2:0] _35587_;
  wire [1:0] _35588_;
  wire [2:0] _35589_;
  wire [1:0] _35590_;
  wire [7:0] _35591_;
  wire [2:0] _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire [7:0] _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire [7:0] _35618_;
  wire [7:0] _35619_;
  wire [7:0] _35620_;
  wire [7:0] _35621_;
  wire [7:0] _35622_;
  wire [7:0] _35623_;
  wire [7:0] _35624_;
  wire [7:0] _35625_;
  wire [7:0] _35626_;
  wire [7:0] _35627_;
  wire [7:0] _35628_;
  wire [7:0] _35629_;
  wire [7:0] _35630_;
  wire [7:0] _35631_;
  wire [7:0] _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire [7:0] _35642_;
  wire _35643_;
  wire [15:0] _35644_;
  wire [31:0] _35645_;
  wire [31:0] _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire [7:0] _35650_;
  wire _35651_;
  wire [2:0] _35652_;
  wire _35653_;
  wire [3:0] _35654_;
  wire [15:0] _35655_;
  wire [15:0] _35656_;
  wire [15:0] _35657_;
  wire [15:0] _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire [7:0] _35662_;
  wire [31:0] _35663_;
  wire [1:0] _35664_;
  wire [2:0] _35665_;
  wire [8:0] _35666_;
  wire [15:0] _35667_;
  wire [15:0] _35668_;
  wire [15:0] _35669_;
  wire [15:0] _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire [1:0] _35687_;
  wire [3:0] _35688_;
  wire [1:0] _35689_;
  wire _35690_;
  wire [7:0] _35691_;
  wire [3:0] _35692_;
  wire [1:0] _35693_;
  wire [22:0] _35694_;
  wire [10:0] _35695_;
  wire [5:0] _35696_;
  wire [2:0] _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire [1:0] _35702_;
  wire [1:0] _35703_;
  wire [1:0] _35704_;
  wire [2:0] _35705_;
  wire [1:0] _35706_;
  wire [1:0] _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire [1:0] _35724_;
  wire [1:0] _35725_;
  wire [1:0] _35726_;
  wire [1:0] _35727_;
  wire [1:0] _35728_;
  wire [1:0] _35729_;
  wire [1:0] _35730_;
  wire [1:0] _35731_;
  wire [1:0] _35732_;
  wire [1:0] _35733_;
  wire [1:0] _35734_;
  wire _35735_;
  wire [1:0] _35736_;
  wire _35737_;
  wire [1:0] _35738_;
  wire _35739_;
  wire [1:0] _35740_;
  wire _35741_;
  wire [1:0] _35742_;
  wire [1:0] _35743_;
  wire [1:0] _35744_;
  wire [1:0] _35745_;
  wire [1:0] _35746_;
  wire [1:0] _35747_;
  wire [1:0] _35748_;
  wire _35749_;
  wire [1:0] _35750_;
  wire _35751_;
  wire [1:0] _35752_;
  wire _35753_;
  wire [1:0] _35754_;
  wire _35755_;
  wire [1:0] _35756_;
  wire _35757_;
  wire [1:0] _35758_;
  wire _35759_;
  wire [1:0] _35760_;
  wire _35761_;
  wire [1:0] _35762_;
  wire _35763_;
  wire [1:0] _35764_;
  wire _35765_;
  wire [1:0] _35766_;
  wire _35767_;
  wire [1:0] _35768_;
  wire _35769_;
  wire [1:0] _35770_;
  wire _35771_;
  wire [1:0] _35772_;
  wire _35773_;
  wire [1:0] _35774_;
  wire _35775_;
  wire [1:0] _35776_;
  wire _35777_;
  wire [1:0] _35778_;
  wire _35779_;
  wire [1:0] _35780_;
  wire _35781_;
  wire [1:0] _35782_;
  wire _35783_;
  wire [1:0] _35784_;
  wire _35785_;
  wire [1:0] _35786_;
  wire _35787_;
  wire [1:0] _35788_;
  wire _35789_;
  wire [1:0] _35790_;
  wire _35791_;
  wire [1:0] _35792_;
  wire _35793_;
  wire [1:0] _35794_;
  wire _35795_;
  wire [1:0] _35796_;
  wire _35797_;
  wire [2:0] _35798_;
  wire _35799_;
  wire [2:0] _35800_;
  wire _35801_;
  wire [2:0] _35802_;
  wire _35803_;
  wire [2:0] _35804_;
  wire _35805_;
  wire [2:0] _35806_;
  wire _35807_;
  wire [2:0] _35808_;
  wire _35809_;
  wire [2:0] _35810_;
  wire _35811_;
  wire [2:0] _35812_;
  wire _35813_;
  wire [2:0] _35814_;
  wire _35815_;
  wire [2:0] _35816_;
  wire [1:0] _35817_;
  wire [2:0] _35818_;
  wire [1:0] _35819_;
  wire [2:0] _35820_;
  wire [1:0] _35821_;
  wire [2:0] _35822_;
  wire [1:0] _35823_;
  wire [2:0] _35824_;
  wire [1:0] _35825_;
  wire [2:0] _35826_;
  wire [2:0] _35827_;
  wire [1:0] _35828_;
  wire [2:0] _35829_;
  wire [1:0] _35830_;
  wire [2:0] _35831_;
  wire [1:0] _35832_;
  wire [2:0] _35833_;
  wire [3:0] _35834_;
  wire [7:0] _35835_;
  wire [2:0] _35836_;
  wire [2:0] _35837_;
  wire [2:0] _35838_;
  wire [7:0] _35839_;
  wire [2:0] _35840_;
  wire [2:0] _35841_;
  wire [2:0] _35842_;
  wire [2:0] _35843_;
  wire [2:0] _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire [15:0] _35939_;
  wire [15:0] _35940_;
  wire [7:0] _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire [2:0] _35949_;
  wire [4:0] _35950_;
  wire [15:0] _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire [1:0] _35955_;
  wire [1:0] _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire [7:0] _36026_;
  wire [15:0] _36027_;
  wire [31:0] _36028_;
  wire [1:0] _36029_;
  wire [1:0] _36030_;
  wire [8:0] _36031_;
  wire [15:0] _36032_;
  wire [15:0] _36033_;
  wire [15:0] _36034_;
  wire [15:0] _36035_;
  wire [15:0] _36036_;
  wire [15:0] _36037_;
  wire [3:0] _36038_;
  wire [3:0] _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire [7:0] _36043_;
  wire [7:0] _36044_;
  wire [7:0] _36045_;
  wire [7:0] _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire [2:0] _36056_;
  wire [2:0] _36057_;
  wire [2:0] _36058_;
  wire [2:0] _36059_;
  wire [2:0] _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire [4:0] _36065_;
  wire [4:0] _36066_;
  wire [4:0] _36067_;
  wire [4:0] _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire [7:0] _36076_;
  wire [7:0] _36077_;
  wire [7:0] _36078_;
  wire [7:0] _36079_;
  wire [7:0] _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire [7:0] _36090_;
  wire [7:0] _36091_;
  wire [7:0] _36092_;
  wire [7:0] _36093_;
  wire [7:0] _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire [7:0] _36103_;
  wire [7:0] _36104_;
  wire [7:0] _36105_;
  wire [7:0] _36106_;
  wire [7:0] _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire [7:0] _36116_;
  wire [7:0] _36117_;
  wire [7:0] _36118_;
  wire [7:0] _36119_;
  wire [7:0] _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire [7:0] _36130_;
  wire [7:0] _36131_;
  wire [7:0] _36132_;
  wire [7:0] _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire [7:0] _36143_;
  wire [7:0] _36144_;
  wire [15:0] _36145_;
  wire [15:0] _36146_;
  wire [15:0] _36147_;
  wire [1:0] _36148_;
  wire _36149_;
  wire [8:0] _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire [15:0] _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire [15:0] _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire [3:0] _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire [31:0] _36256_;
  wire [1:0] _36257_;
  wire [1:0] _36258_;
  wire [1:0] _36259_;
  wire [1:0] _36260_;
  wire [1:0] _36261_;
  wire [3:0] _36262_;
  wire [1:0] _36263_;
  wire [3:0] _36264_;
  wire [1:0] _36265_;
  wire [3:0] _36266_;
  wire [1:0] _36267_;
  wire [3:0] _36268_;
  wire [1:0] _36269_;
  wire [3:0] _36270_;
  wire [1:0] _36271_;
  wire [3:0] _36272_;
  wire [1:0] _36273_;
  wire [3:0] _36274_;
  wire [1:0] _36275_;
  wire [3:0] _36276_;
  wire [1:0] _36277_;
  wire [3:0] _36278_;
  wire [1:0] _36279_;
  wire [3:0] _36280_;
  wire [3:0] _36281_;
  wire [3:0] _36282_;
  wire [1:0] _36283_;
  wire [1:0] _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire [63:0] _36294_;
  wire [7:0] _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire [15:0] _36303_;
  wire [7:0] _36304_;
  wire _36305_;
  wire [15:0] _36306_;
  wire [7:0] _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire [7:0] _36313_;
  wire [7:0] _36314_;
  wire [7:0] _36315_;
  wire [7:0] _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire [3:0] _36640_;
  wire [1:0] _36641_;
  wire [7:0] _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire [7:0] _36653_;
  wire [7:0] _36654_;
  wire [7:0] _36655_;
  wire [7:0] _36656_;
  wire [7:0] _36657_;
  wire [7:0] _36658_;
  wire [7:0] _36659_;
  wire [7:0] _36660_;
  wire [7:0] _36661_;
  wire [7:0] _36662_;
  wire [7:0] _36663_;
  wire [7:0] _36664_;
  wire [7:0] _36665_;
  wire [7:0] _36666_;
  wire [7:0] _36667_;
  wire [7:0] _36668_;
  wire [7:0] _36669_;
  wire [7:0] _36670_;
  wire [7:0] _36671_;
  wire [7:0] _36672_;
  wire [7:0] _36673_;
  wire [7:0] _36674_;
  wire [7:0] _36675_;
  wire [7:0] _36676_;
  wire [7:0] _36677_;
  wire [7:0] _36678_;
  wire [7:0] _36679_;
  wire [7:0] _36680_;
  wire [7:0] _36681_;
  wire [7:0] _36682_;
  wire [7:0] _36683_;
  wire [7:0] _36684_;
  wire [7:0] _36685_;
  wire [7:0] _36686_;
  wire [7:0] _36687_;
  wire [7:0] _36688_;
  wire [7:0] _36689_;
  wire [7:0] _36690_;
  wire [7:0] _36691_;
  wire [7:0] _36692_;
  wire [7:0] _36693_;
  wire [7:0] _36694_;
  wire [7:0] _36695_;
  wire [7:0] _36696_;
  wire [7:0] _36697_;
  wire [7:0] _36698_;
  wire [7:0] _36699_;
  wire [7:0] _36700_;
  wire [7:0] _36701_;
  wire [7:0] _36702_;
  wire [7:0] _36703_;
  wire [7:0] _36704_;
  wire [7:0] _36705_;
  wire [7:0] _36706_;
  wire [7:0] _36707_;
  wire [7:0] _36708_;
  wire [7:0] _36709_;
  wire [7:0] _36710_;
  wire [7:0] _36711_;
  wire [7:0] _36712_;
  wire [7:0] _36713_;
  wire [7:0] _36714_;
  wire [7:0] _36715_;
  wire [7:0] _36716_;
  wire [7:0] _36717_;
  wire [7:0] _36718_;
  wire [7:0] _36719_;
  wire [7:0] _36720_;
  wire [7:0] _36721_;
  wire [7:0] _36722_;
  wire [7:0] _36723_;
  wire [7:0] _36724_;
  wire [7:0] _36725_;
  wire [7:0] _36726_;
  wire [7:0] _36727_;
  wire [7:0] _36728_;
  wire [7:0] _36729_;
  wire [7:0] _36730_;
  wire [7:0] _36731_;
  wire [7:0] _36732_;
  wire [7:0] _36733_;
  wire [7:0] _36734_;
  wire [7:0] _36735_;
  wire [7:0] _36736_;
  wire [7:0] _36737_;
  wire [7:0] _36738_;
  wire [7:0] _36739_;
  wire [7:0] _36740_;
  wire [7:0] _36741_;
  wire [7:0] _36742_;
  wire [7:0] _36743_;
  wire [7:0] _36744_;
  wire [7:0] _36745_;
  wire [7:0] _36746_;
  wire [7:0] _36747_;
  wire [7:0] _36748_;
  wire [7:0] _36749_;
  wire [7:0] _36750_;
  wire [7:0] _36751_;
  wire [7:0] _36752_;
  wire [7:0] _36753_;
  wire [7:0] _36754_;
  wire [7:0] _36755_;
  wire [7:0] _36756_;
  wire [7:0] _36757_;
  wire [7:0] _36758_;
  wire [7:0] _36759_;
  wire [7:0] _36760_;
  wire [7:0] _36761_;
  wire [7:0] _36762_;
  wire [7:0] _36763_;
  wire [7:0] _36764_;
  wire [7:0] _36765_;
  wire [7:0] _36766_;
  wire [7:0] _36767_;
  wire [7:0] _36768_;
  wire [7:0] _36769_;
  wire [7:0] _36770_;
  wire [7:0] _36771_;
  wire [7:0] _36772_;
  wire [7:0] _36773_;
  wire [7:0] _36774_;
  wire [7:0] _36775_;
  wire [7:0] _36776_;
  wire [7:0] _36777_;
  wire [7:0] _36778_;
  wire [7:0] _36779_;
  wire [7:0] _36780_;
  wire [7:0] _36781_;
  wire [7:0] _36782_;
  wire [7:0] _36783_;
  wire [7:0] _36784_;
  wire [7:0] _36785_;
  wire [7:0] _36786_;
  wire [7:0] _36787_;
  wire [7:0] _36788_;
  wire [7:0] _36789_;
  wire [7:0] _36790_;
  wire [7:0] _36791_;
  wire [7:0] _36792_;
  wire [7:0] _36793_;
  wire [7:0] _36794_;
  wire [7:0] _36795_;
  wire [7:0] _36796_;
  wire [7:0] _36797_;
  wire [7:0] _36798_;
  wire [7:0] _36799_;
  wire [7:0] _36800_;
  wire [7:0] _36801_;
  wire [7:0] _36802_;
  wire [7:0] _36803_;
  wire [7:0] _36804_;
  wire [7:0] _36805_;
  wire [7:0] _36806_;
  wire [7:0] _36807_;
  wire [7:0] _36808_;
  wire [7:0] _36809_;
  wire [7:0] _36810_;
  wire [7:0] _36811_;
  wire [7:0] _36812_;
  wire [7:0] _36813_;
  wire [7:0] _36814_;
  wire [7:0] _36815_;
  wire [7:0] _36816_;
  wire [7:0] _36817_;
  wire [7:0] _36818_;
  wire [7:0] _36819_;
  wire [7:0] _36820_;
  wire [7:0] _36821_;
  wire [7:0] _36822_;
  wire [7:0] _36823_;
  wire [7:0] _36824_;
  wire [7:0] _36825_;
  wire [7:0] _36826_;
  wire [7:0] _36827_;
  wire [7:0] _36828_;
  wire [7:0] _36829_;
  wire [7:0] _36830_;
  wire [7:0] _36831_;
  wire [7:0] _36832_;
  wire [7:0] _36833_;
  wire [7:0] _36834_;
  wire [7:0] _36835_;
  wire [7:0] _36836_;
  wire [7:0] _36837_;
  wire [7:0] _36838_;
  wire [7:0] _36839_;
  wire [7:0] _36840_;
  wire [7:0] _36841_;
  wire [7:0] _36842_;
  wire [7:0] _36843_;
  wire [7:0] _36844_;
  wire [7:0] _36845_;
  wire [7:0] _36846_;
  wire [7:0] _36847_;
  wire [7:0] _36848_;
  wire [7:0] _36849_;
  wire [7:0] _36850_;
  wire [7:0] _36851_;
  wire [7:0] _36852_;
  wire [7:0] _36853_;
  wire [7:0] _36854_;
  wire [7:0] _36855_;
  wire [7:0] _36856_;
  wire [7:0] _36857_;
  wire [7:0] _36858_;
  wire [7:0] _36859_;
  wire [7:0] _36860_;
  wire [7:0] _36861_;
  wire [7:0] _36862_;
  wire [7:0] _36863_;
  wire [7:0] _36864_;
  wire [7:0] _36865_;
  wire [7:0] _36866_;
  wire [7:0] _36867_;
  wire [7:0] _36868_;
  wire [7:0] _36869_;
  wire [7:0] _36870_;
  wire [7:0] _36871_;
  wire [7:0] _36872_;
  wire [7:0] _36873_;
  wire [7:0] _36874_;
  wire [7:0] _36875_;
  wire [7:0] _36876_;
  wire [7:0] _36877_;
  wire [7:0] _36878_;
  wire [7:0] _36879_;
  wire [7:0] _36880_;
  wire [7:0] _36881_;
  wire [7:0] _36882_;
  wire [7:0] _36883_;
  wire [7:0] _36884_;
  wire [7:0] _36885_;
  wire [7:0] _36886_;
  wire [7:0] _36887_;
  wire [7:0] _36888_;
  wire [7:0] _36889_;
  wire [7:0] _36890_;
  wire [7:0] _36891_;
  wire [7:0] _36892_;
  wire [7:0] _36893_;
  wire [7:0] _36894_;
  wire [7:0] _36895_;
  wire [7:0] _36896_;
  wire [7:0] _36897_;
  wire [7:0] _36898_;
  wire [7:0] _36899_;
  wire [7:0] _36900_;
  wire [7:0] _36901_;
  wire [7:0] _36902_;
  wire [7:0] _36903_;
  wire [7:0] _36904_;
  wire [7:0] _36905_;
  wire [7:0] _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire [7:0] _37163_;
  wire [7:0] _37164_;
  wire [7:0] _37165_;
  wire [7:0] _37166_;
  wire [7:0] _37167_;
  wire [7:0] _37168_;
  wire [7:0] _37169_;
  wire [7:0] _37170_;
  wire [7:0] _37171_;
  wire [7:0] _37172_;
  wire [7:0] _37173_;
  wire [7:0] _37174_;
  wire [7:0] _37175_;
  wire [7:0] _37176_;
  wire [7:0] _37177_;
  wire [7:0] _37178_;
  wire [7:0] _37179_;
  wire [7:0] _37180_;
  wire [7:0] _37181_;
  wire [7:0] _37182_;
  wire [7:0] _37183_;
  wire [7:0] _37184_;
  wire [7:0] _37185_;
  wire [7:0] _37186_;
  wire [7:0] _37187_;
  wire [7:0] _37188_;
  wire [7:0] _37189_;
  wire [7:0] _37190_;
  wire [7:0] _37191_;
  wire [7:0] _37192_;
  wire [7:0] _37193_;
  wire [7:0] _37194_;
  wire [7:0] _37195_;
  wire [7:0] _37196_;
  wire [7:0] _37197_;
  wire [7:0] _37198_;
  wire [7:0] _37199_;
  wire [7:0] _37200_;
  wire [7:0] _37201_;
  wire [7:0] _37202_;
  wire [7:0] _37203_;
  wire [7:0] _37204_;
  wire [7:0] _37205_;
  wire [7:0] _37206_;
  wire [7:0] _37207_;
  wire [7:0] _37208_;
  wire [7:0] _37209_;
  wire [7:0] _37210_;
  wire [7:0] _37211_;
  wire [7:0] _37212_;
  wire [7:0] _37213_;
  wire [7:0] _37214_;
  wire [7:0] _37215_;
  wire [7:0] _37216_;
  wire [7:0] _37217_;
  wire [7:0] _37218_;
  wire [7:0] _37219_;
  wire [7:0] _37220_;
  wire [7:0] _37221_;
  wire [7:0] _37222_;
  wire [7:0] _37223_;
  wire [7:0] _37224_;
  wire [7:0] _37225_;
  wire [7:0] _37226_;
  wire [7:0] _37227_;
  wire [7:0] _37228_;
  wire [7:0] _37229_;
  wire [7:0] _37230_;
  wire [7:0] _37231_;
  wire [7:0] _37232_;
  wire [7:0] _37233_;
  wire [7:0] _37234_;
  wire [7:0] _37235_;
  wire [7:0] _37236_;
  wire [7:0] _37237_;
  wire [7:0] _37238_;
  wire [7:0] _37239_;
  wire [7:0] _37240_;
  wire [7:0] _37241_;
  wire [7:0] _37242_;
  wire [7:0] _37243_;
  wire [7:0] _37244_;
  wire [7:0] _37245_;
  wire [7:0] _37246_;
  wire [7:0] _37247_;
  wire [7:0] _37248_;
  wire [7:0] _37249_;
  wire [7:0] _37250_;
  wire [7:0] _37251_;
  wire [7:0] _37252_;
  wire [7:0] _37253_;
  wire [7:0] _37254_;
  wire [7:0] _37255_;
  wire [7:0] _37256_;
  wire [7:0] _37257_;
  wire [7:0] _37258_;
  wire [7:0] _37259_;
  wire [7:0] _37260_;
  wire [7:0] _37261_;
  wire [7:0] _37262_;
  wire [7:0] _37263_;
  wire [7:0] _37264_;
  wire [7:0] _37265_;
  wire [7:0] _37266_;
  wire [7:0] _37267_;
  wire [7:0] _37268_;
  wire [7:0] _37269_;
  wire [7:0] _37270_;
  wire [7:0] _37271_;
  wire [7:0] _37272_;
  wire [7:0] _37273_;
  wire [7:0] _37274_;
  wire [7:0] _37275_;
  wire [7:0] _37276_;
  wire [7:0] _37277_;
  wire [7:0] _37278_;
  wire [7:0] _37279_;
  wire [7:0] _37280_;
  wire [7:0] _37281_;
  wire [7:0] _37282_;
  wire [7:0] _37283_;
  wire [7:0] _37284_;
  wire [7:0] _37285_;
  wire [7:0] _37286_;
  wire [7:0] _37287_;
  wire [7:0] _37288_;
  wire [7:0] _37289_;
  wire [7:0] _37290_;
  wire [7:0] _37291_;
  wire [7:0] _37292_;
  wire [7:0] _37293_;
  wire [7:0] _37294_;
  wire [7:0] _37295_;
  wire [7:0] _37296_;
  wire [7:0] _37297_;
  wire [7:0] _37298_;
  wire [7:0] _37299_;
  wire [7:0] _37300_;
  wire [7:0] _37301_;
  wire [7:0] _37302_;
  wire [7:0] _37303_;
  wire [7:0] _37304_;
  wire [7:0] _37305_;
  wire [7:0] _37306_;
  wire [7:0] _37307_;
  wire [7:0] _37308_;
  wire [7:0] _37309_;
  wire [7:0] _37310_;
  wire [7:0] _37311_;
  wire [7:0] _37312_;
  wire [7:0] _37313_;
  wire [7:0] _37314_;
  wire [7:0] _37315_;
  wire [7:0] _37316_;
  wire [7:0] _37317_;
  wire [7:0] _37318_;
  wire [7:0] _37319_;
  wire [7:0] _37320_;
  wire [7:0] _37321_;
  wire [7:0] _37322_;
  wire [7:0] _37323_;
  wire [7:0] _37324_;
  wire [7:0] _37325_;
  wire [7:0] _37326_;
  wire [7:0] _37327_;
  wire [7:0] _37328_;
  wire [7:0] _37329_;
  wire [7:0] _37330_;
  wire [7:0] _37331_;
  wire [7:0] _37332_;
  wire [7:0] _37333_;
  wire [7:0] _37334_;
  wire [7:0] _37335_;
  wire [7:0] _37336_;
  wire [7:0] _37337_;
  wire [7:0] _37338_;
  wire [7:0] _37339_;
  wire [7:0] _37340_;
  wire [7:0] _37341_;
  wire [7:0] _37342_;
  wire [7:0] _37343_;
  wire [7:0] _37344_;
  wire [7:0] _37345_;
  wire [7:0] _37346_;
  wire [7:0] _37347_;
  wire [7:0] _37348_;
  wire [7:0] _37349_;
  wire [7:0] _37350_;
  wire [7:0] _37351_;
  wire [7:0] _37352_;
  wire [7:0] _37353_;
  wire [7:0] _37354_;
  wire [7:0] _37355_;
  wire [7:0] _37356_;
  wire [7:0] _37357_;
  wire [7:0] _37358_;
  wire [7:0] _37359_;
  wire [7:0] _37360_;
  wire [7:0] _37361_;
  wire [7:0] _37362_;
  wire [7:0] _37363_;
  wire [7:0] _37364_;
  wire [7:0] _37365_;
  wire [7:0] _37366_;
  wire [7:0] _37367_;
  wire [7:0] _37368_;
  wire [7:0] _37369_;
  wire [7:0] _37370_;
  wire [7:0] _37371_;
  wire [7:0] _37372_;
  wire [7:0] _37373_;
  wire [7:0] _37374_;
  wire [7:0] _37375_;
  wire [7:0] _37376_;
  wire [7:0] _37377_;
  wire [7:0] _37378_;
  wire [7:0] _37379_;
  wire [7:0] _37380_;
  wire [7:0] _37381_;
  wire [7:0] _37382_;
  wire [7:0] _37383_;
  wire [7:0] _37384_;
  wire [7:0] _37385_;
  wire [7:0] _37386_;
  wire [7:0] _37387_;
  wire [7:0] _37388_;
  wire [7:0] _37389_;
  wire [7:0] _37390_;
  wire [7:0] _37391_;
  wire [7:0] _37392_;
  wire [7:0] _37393_;
  wire [7:0] _37394_;
  wire [7:0] _37395_;
  wire [7:0] _37396_;
  wire [7:0] _37397_;
  wire [7:0] _37398_;
  wire [7:0] _37399_;
  wire [7:0] _37400_;
  wire [7:0] _37401_;
  wire [7:0] _37402_;
  wire [7:0] _37403_;
  wire [7:0] _37404_;
  wire [7:0] _37405_;
  wire [7:0] _37406_;
  wire [7:0] _37407_;
  wire [7:0] _37408_;
  wire [7:0] _37409_;
  wire [7:0] _37410_;
  wire [7:0] _37411_;
  wire [7:0] _37412_;
  wire [7:0] _37413_;
  wire [7:0] _37414_;
  wire [7:0] _37415_;
  wire [7:0] _37416_;
  wire [7:0] _37417_;
  wire [7:0] _37418_;
  wire [7:0] _37419_;
  wire [7:0] _37420_;
  wire [7:0] _37421_;
  wire _37422_;
  wire [8:0] _37423_;
  wire [7:0] _37424_;
  wire _37425_;
  wire [3:0] _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire [3:0] _37452_;
  wire [1:0] _37453_;
  wire [3:0] _37454_;
  wire [1:0] _37455_;
  wire [3:0] _37456_;
  wire [1:0] _37457_;
  wire [1:0] _37458_;
  wire [1:0] _37459_;
  wire [3:0] _37460_;
  wire [1:0] _37461_;
  wire [3:0] _37462_;
  wire [1:0] _37463_;
  wire [1:0] _37464_;
  wire [3:0] _37465_;
  wire [1:0] _37466_;
  wire [3:0] _37467_;
  wire [1:0] _37468_;
  wire [3:0] _37469_;
  wire [1:0] _37470_;
  wire [1:0] _37471_;
  wire [3:0] _37472_;
  wire [1:0] _37473_;
  wire [3:0] _37474_;
  wire [1:0] _37475_;
  wire [1:0] _37476_;
  wire [1:0] _37477_;
  wire [1:0] _37478_;
  wire [1:0] _37479_;
  wire [1:0] _37480_;
  wire _37481_;
  wire [1:0] _37482_;
  wire _37483_;
  wire [1:0] _37484_;
  wire _37485_;
  wire _37486_;
  wire [1:0] _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire [1:0] _37491_;
  wire _37492_;
  wire [1:0] _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire [1:0] _37499_;
  wire _37500_;
  wire _37501_;
  wire [3:0] _37502_;
  wire [1:0] _37503_;
  wire [1:0] _37504_;
  wire [12:0] _37505_;
  wire [5:0] _37506_;
  wire [2:0] _37507_;
  wire [1:0] _37508_;
  wire [12:0] _37509_;
  wire [5:0] _37510_;
  wire [2:0] _37511_;
  wire [1:0] _37512_;
  wire [12:0] _37513_;
  wire [5:0] _37514_;
  wire [2:0] _37515_;
  wire [1:0] _37516_;
  wire [12:0] _37517_;
  wire [5:0] _37518_;
  wire [2:0] _37519_;
  wire [1:0] _37520_;
  wire [12:0] _37521_;
  wire [5:0] _37522_;
  wire [2:0] _37523_;
  wire [1:0] _37524_;
  wire [12:0] _37525_;
  wire [5:0] _37526_;
  wire [2:0] _37527_;
  wire [1:0] _37528_;
  wire [12:0] _37529_;
  wire [5:0] _37530_;
  wire [2:0] _37531_;
  wire [1:0] _37532_;
  wire [12:0] _37533_;
  wire [5:0] _37534_;
  wire [2:0] _37535_;
  wire [1:0] _37536_;
  wire [12:0] _37537_;
  wire [5:0] _37538_;
  wire [2:0] _37539_;
  wire [1:0] _37540_;
  wire [5:0] _37541_;
  wire [2:0] _37542_;
  wire _37543_;
  wire [5:0] _37544_;
  wire [2:0] _37545_;
  wire _37546_;
  wire [7:0] _37547_;
  wire [7:0] _37548_;
  wire [7:0] _37549_;
  wire [7:0] _37550_;
  wire [7:0] _37551_;
  wire [7:0] _37552_;
  wire [1:0] _37553_;
  wire [1:0] _37554_;
  wire [1:0] _37555_;
  wire [4:0] _37556_;
  wire [7:0] _37557_;
  wire [3:0] _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire [3:0] _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire [7:0] _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire [7:0] _37670_;
  wire _37671_;
  wire [7:0] _37672_;
  wire _37673_;
  wire [7:0] _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire [3:0] _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire [7:0] _37707_;
  wire [7:0] _37708_;
  wire [7:0] _37709_;
  wire [7:0] _37710_;
  wire [7:0] _37711_;
  wire [7:0] _37712_;
  wire [7:0] _37713_;
  wire [7:0] _37714_;
  wire [7:0] _37715_;
  wire [7:0] _37716_;
  wire [7:0] _37717_;
  wire [7:0] _37718_;
  wire [7:0] _37719_;
  wire [7:0] _37720_;
  wire [7:0] _37721_;
  wire [7:0] _37722_;
  wire [7:0] _37723_;
  wire [7:0] _37724_;
  wire [7:0] _37725_;
  wire [7:0] _37726_;
  wire [7:0] _37727_;
  wire [7:0] _37728_;
  wire [7:0] _37729_;
  wire [7:0] _37730_;
  wire [7:0] _37731_;
  wire [7:0] _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire [7:0] _37742_;
  wire [7:0] _37743_;
  wire [7:0] _37744_;
  wire [7:0] _37745_;
  wire [7:0] _37746_;
  wire [7:0] _37747_;
  wire [7:0] _37748_;
  wire [7:0] _37749_;
  wire [7:0] _37750_;
  wire [7:0] _37751_;
  wire [7:0] _37752_;
  wire [7:0] _37753_;
  wire [7:0] _37754_;
  wire [7:0] _37755_;
  wire [7:0] _37756_;
  wire [7:0] _37757_;
  wire [7:0] _37758_;
  wire [7:0] _37759_;
  wire [7:0] _37760_;
  wire [7:0] _37761_;
  wire [7:0] _37762_;
  wire [7:0] _37763_;
  wire [7:0] _37764_;
  wire [7:0] _37765_;
  wire [7:0] _37766_;
  wire [7:0] _37767_;
  wire [7:0] _37768_;
  wire [7:0] _37769_;
  wire [7:0] _37770_;
  wire [7:0] _37771_;
  wire [7:0] _37772_;
  wire [7:0] _37773_;
  wire [7:0] _37774_;
  wire [7:0] _37775_;
  wire [7:0] _37776_;
  wire [7:0] _37777_;
  wire [7:0] _37778_;
  wire [7:0] _37779_;
  wire [7:0] _37780_;
  wire [7:0] _37781_;
  wire [7:0] _37782_;
  wire [7:0] _37783_;
  wire [7:0] _37784_;
  wire [7:0] _37785_;
  wire [7:0] _37786_;
  wire [7:0] _37787_;
  wire [7:0] _37788_;
  wire [7:0] _37789_;
  wire [7:0] _37790_;
  wire [7:0] _37791_;
  wire [7:0] _37792_;
  wire [7:0] _37793_;
  wire [7:0] _37794_;
  wire [7:0] _37795_;
  wire [7:0] _37796_;
  wire _37797_;
  wire [3:0] _37798_;
  wire [1:0] _37799_;
  wire [3:0] _37800_;
  wire [1:0] _37801_;
  wire _37802_;
  wire [2:0] _37803_;
  wire [1:0] _37804_;
  wire [2:0] _37805_;
  wire [1:0] _37806_;
  wire [2:0] _37807_;
  wire [1:0] _37808_;
  wire [2:0] _37809_;
  wire [1:0] _37810_;
  wire [2:0] _37811_;
  wire [1:0] _37812_;
  wire [2:0] _37813_;
  wire [1:0] _37814_;
  wire [2:0] _37815_;
  wire [1:0] _37816_;
  wire [2:0] _37817_;
  wire [1:0] _37818_;
  wire [2:0] _37819_;
  wire [1:0] _37820_;
  wire [7:0] _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire [7:0] _37829_;
  wire [7:0] _37830_;
  wire [7:0] _37831_;
  wire [7:0] _37832_;
  wire [7:0] _37833_;
  wire [7:0] _37834_;
  wire [7:0] _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire [7:0] _37845_;
  wire [1:0] _37846_;
  wire [1:0] _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire [7:0] _37885_;
  wire [7:0] _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire [1:0] _37891_;
  wire [1:0] _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire [7:0] _37897_;
  wire [7:0] _37898_;
  wire [7:0] _37899_;
  wire [7:0] _37900_;
  wire [1:0] _37901_;
  wire [1:0] _37902_;
  wire [1:0] _37903_;
  wire _37904_;
  wire [7:0] _37905_;
  wire [7:0] _37906_;
  wire [2:0] _37907_;
  wire [2:0] _37908_;
  wire _37909_;
  wire _37910_;
  wire [3:0] _37911_;
  wire _37912_;
  wire _37913_;
  wire [1:0] _37914_;
  wire [5:0] _37915_;
  wire [5:0] _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire [2:0] _37943_;
  wire _37944_;
  wire [2:0] _37945_;
  wire _37946_;
  wire [3:0] _37947_;
  wire [1:0] _37948_;
  wire [3:0] _37949_;
  wire [1:0] _37950_;
  wire [1:0] _37951_;
  wire _37952_;
  wire [3:0] _37953_;
  wire [1:0] _37954_;
  wire [1:0] _37955_;
  wire _37956_;
  wire _37957_;
  wire [1:0] _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire [2:0] _37963_;
  wire [1:0] _37964_;
  wire [7:0] _37965_;
  wire [2:0] _37966_;
  wire [2:0] _37967_;
  wire [2:0] _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire [2:0] _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire [7:0] _38059_;
  wire [7:0] _38060_;
  wire [7:0] _38061_;
  wire [7:0] _38062_;
  wire [7:0] _38063_;
  wire [7:0] _38064_;
  wire [7:0] _38065_;
  wire [7:0] _38066_;
  wire [7:0] _38067_;
  wire [7:0] _38068_;
  wire [7:0] _38069_;
  wire [7:0] _38070_;
  wire [7:0] _38071_;
  wire [7:0] _38072_;
  wire [1:0] _38073_;
  wire [1:0] _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire [2:0] _38078_;
  wire [2:0] _38079_;
  wire [2:0] _38080_;
  wire [2:0] _38081_;
  wire [2:0] _38082_;
  wire [2:0] _38083_;
  wire [2:0] _38084_;
  wire [2:0] _38085_;
  wire [2:0] _38086_;
  wire [2:0] _38087_;
  wire [2:0] _38088_;
  wire [2:0] _38089_;
  wire [2:0] _38090_;
  wire [2:0] _38091_;
  wire [2:0] _38092_;
  wire [2:0] _38093_;
  wire [2:0] _38094_;
  wire [2:0] _38095_;
  wire [2:0] _38096_;
  wire [2:0] _38097_;
  wire [2:0] _38098_;
  wire [2:0] _38099_;
  wire [2:0] _38100_;
  wire [2:0] _38101_;
  wire [2:0] _38102_;
  wire [2:0] _38103_;
  wire [2:0] _38104_;
  wire [2:0] _38105_;
  wire [2:0] _38106_;
  wire [2:0] _38107_;
  wire [2:0] _38108_;
  wire [2:0] _38109_;
  wire [2:0] _38110_;
  wire [2:0] _38111_;
  wire [1:0] _38112_;
  wire [1:0] _38113_;
  wire [1:0] _38114_;
  wire [1:0] _38115_;
  wire [1:0] _38116_;
  wire [1:0] _38117_;
  wire [1:0] _38118_;
  wire [1:0] _38119_;
  wire [1:0] _38120_;
  wire [7:0] _38121_;
  wire [7:0] _38122_;
  wire [7:0] _38123_;
  wire [7:0] _38124_;
  wire [1:0] _38125_;
  wire _38126_;
  wire [1:0] _38127_;
  wire _38128_;
  wire [1:0] _38129_;
  wire _38130_;
  wire _38131_;
  wire [1:0] _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire [6:0] _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire [3:0] _38275_;
  wire [1:0] _38276_;
  wire _38277_;
  wire _38278_;
  wire [1:0] _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire [7:0] _38308_;
  wire [7:0] _38309_;
  wire [7:0] _38310_;
  wire [7:0] _38311_;
  wire _38312_;
  wire [1:0] _38313_;
  wire _38314_;
  wire _38315_;
  wire [2:0] _38316_;
  wire [2:0] _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire [7:0] _38322_;
  wire [7:0] _38323_;
  wire [7:0] _38324_;
  wire [7:0] _38325_;
  wire [7:0] _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire [7:0] _38331_;
  wire [7:0] _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire [7:0] _38348_;
  wire [7:0] _38349_;
  wire [7:0] _38350_;
  wire [7:0] _38351_;
  wire [7:0] _38352_;
  wire [13:0] _38353_;
  wire [16:0] _38354_;
  wire [8:0] _38355_;
  wire [13:0] _38356_;
  wire [16:0] _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire [3:0] _38373_;
  wire [1:0] _38374_;
  wire [3:0] _38375_;
  wire [1:0] _38376_;
  wire [3:0] _38377_;
  wire [1:0] _38378_;
  wire [3:0] _38379_;
  wire [1:0] _38380_;
  wire [3:0] _38381_;
  wire [1:0] _38382_;
  wire [1:0] _38383_;
  wire [3:0] _38384_;
  wire [1:0] _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire [7:0] _38411_;
  wire [7:0] _38412_;
  wire [7:0] _38413_;
  wire [7:0] _38414_;
  wire [7:0] _38415_;
  wire [1:0] _38416_;
  wire [1:0] _38417_;
  wire [1:0] _38418_;
  wire [1:0] _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire [4:0] _38447_;
  wire [4:0] _38448_;
  wire [4:0] _38449_;
  wire _38450_;
  wire [4:0] _38451_;
  wire _38452_;
  wire _38453_;
  wire [4:0] _38454_;
  wire [2:0] _38455_;
  wire [2:0] _38456_;
  wire [2:0] _38457_;
  wire [2:0] _38458_;
  wire [2:0] _38459_;
  wire [7:0] _38460_;
  wire [7:0] _38461_;
  wire [7:0] _38462_;
  wire [7:0] _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire [4:0] _38478_;
  wire [4:0] _38479_;
  wire [4:0] _38480_;
  wire [4:0] _38481_;
  wire [4:0] _38482_;
  wire [2:0] _38483_;
  wire [2:0] _38484_;
  wire [2:0] _38485_;
  wire [2:0] _38486_;
  wire [2:0] _38487_;
  wire [7:0] _38488_;
  wire [7:0] _38489_;
  wire [7:0] _38490_;
  wire [7:0] _38491_;
  wire [7:0] _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire [13:0] _38496_;
  wire [16:0] _38497_;
  wire [7:0] _38498_;
  wire [7:0] _38499_;
  wire [8:0] _38500_;
  wire [13:0] _38501_;
  wire [16:0] _38502_;
  wire [4:0] _38503_;
  wire [4:0] _38504_;
  wire [4:0] _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire [2:0] _38512_;
  wire [2:0] _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire [7:0] _38518_;
  wire [7:0] _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire [4:0] _38538_;
  wire [4:0] _38539_;
  wire [4:0] _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire [2:0] _38546_;
  wire [2:0] _38547_;
  wire [2:0] _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire [7:0] _38552_;
  wire [7:0] _38553_;
  wire [7:0] _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire [7:0] _38611_;
  wire [7:0] _38612_;
  wire _38613_;
  wire [7:0] _38614_;
  wire _38615_;
  wire _38616_;
  wire [7:0] _38617_;
  wire [7:0] _38618_;
  wire [16:0] _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire [1:0] _38636_;
  wire _38637_;
  wire [1:0] _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire [7:0] _38658_;
  wire [7:0] _38659_;
  wire [7:0] _38660_;
  wire [7:0] _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire [7:0] _38667_;
  wire [7:0] _38668_;
  wire [7:0] _38669_;
  wire [7:0] _38670_;
  wire [7:0] _38671_;
  wire [7:0] _38672_;
  wire [7:0] _38673_;
  wire [7:0] _38674_;
  wire [7:0] _38675_;
  wire [7:0] _38676_;
  wire [7:0] _38677_;
  wire [7:0] _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire [16:0] _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire [7:0] _38718_;
  wire [3:0] _38719_;
  wire _38720_;
  wire _38721_;
  wire [1:0] _38722_;
  wire _38723_;
  wire [7:0] _38724_;
  wire [11:0] _38725_;
  wire [10:0] _38726_;
  wire [7:0] _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire [3:0] _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire [3:0] _38737_;
  wire [3:0] _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire [4:0] _38756_;
  wire [1:0] _38757_;
  wire _38758_;
  wire [1:0] _38759_;
  wire [2:0] _38760_;
  wire [1:0] _38761_;
  wire [1:0] _38762_;
  wire [1:0] _38763_;
  wire [1:0] _38764_;
  wire [3:0] _38765_;
  wire [3:0] _38766_;
  wire [1:0] _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire [3:0] _38816_;
  wire [3:0] _38817_;
  wire [3:0] _38818_;
  wire [3:0] _38819_;
  wire [11:0] _38820_;
  wire [11:0] _38821_;
  wire [11:0] _38822_;
  wire [11:0] _38823_;
  wire [11:0] _38824_;
  wire [11:0] _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire [3:0] _38839_;
  wire [3:0] _38840_;
  wire [10:0] _38841_;
  wire [10:0] _38842_;
  wire [10:0] _38843_;
  wire [10:0] _38844_;
  wire [10:0] _38845_;
  wire [10:0] _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire [3:0] _38876_;
  wire [3:0] _38877_;
  wire [10:0] _38878_;
  wire [10:0] _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  input clk;
  wire [15:0] cxrom_addr;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [3:0] \oc8051_symbolic_cxrom1.addr0 ;
  wire [3:0] \oc8051_symbolic_cxrom1.addr1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.addr2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.addr3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [15:0] \oc8051_symbolic_cxrom1.cxrom_addr ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [7:0] \oc8051_symbolic_cxrom1.op_out ;
  wire \oc8051_symbolic_cxrom1.op_valid ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc11 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc13 ;
  wire \oc8051_symbolic_cxrom1.pc1_valid ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc21 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc23 ;
  wire \oc8051_symbolic_cxrom1.pc2_valid ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.alu_cy ;
  wire [3:0] \oc8051_top_1.alu_op ;
  wire [1:0] \oc8051_top_1.bank_sel ;
  wire \oc8051_top_1.bit_addr ;
  wire \oc8051_top_1.bit_addr_o ;
  wire \oc8051_top_1.bit_data ;
  wire \oc8051_top_1.bit_out ;
  wire [1:0] \oc8051_top_1.comp_sel ;
  wire \oc8051_top_1.comp_wait ;
  wire [15:0] \oc8051_top_1.cxrom_addr ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.des1 ;
  wire [7:0] \oc8051_top_1.des2 ;
  wire \oc8051_top_1.desAc ;
  wire \oc8051_top_1.desCy ;
  wire \oc8051_top_1.desOv ;
  wire [7:0] \oc8051_top_1.des_acc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire \oc8051_top_1.eq ;
  wire \oc8051_top_1.iack_i ;
  wire [15:0] \oc8051_top_1.iadr_o ;
  wire [31:0] \oc8051_top_1.idat_i ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.intr ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.mem_wait ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.add1 ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.add2 ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.add3 ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.add4 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.add5 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.add6 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.add7 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.add8 ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.add9 ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.adda ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.addb ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.addc ;
  wire \oc8051_top_1.oc8051_alu1.bit_in ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.dec ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.desAc ;
  wire \oc8051_top_1.oc8051_alu1.desCy ;
  wire \oc8051_top_1.oc8051_alu1.desOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.des_acc ;
  wire \oc8051_top_1.oc8051_alu1.divOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.enable_div ;
  wire \oc8051_top_1.oc8051_alu1.enable_mul ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.inc ;
  wire \oc8051_top_1.oc8051_alu1.mulOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.desOv ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.enable ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.rem1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.rem2 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 ;
  wire [8:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.sub0 ;
  wire [8:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.sub1 ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.desOv ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.enable ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.shifted ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.op_code ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.src1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.src2 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.src3 ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire \oc8051_top_1.oc8051_alu1.srcCy ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.sub1 ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.sub2 ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.sub3 ;
  wire [4:0] \oc8051_top_1.oc8051_alu1.sub4 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.sub5 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.sub6 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.sub7 ;
  wire [3:0] \oc8051_top_1.oc8051_alu1.sub8 ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.sub9 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.sub_result ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.suba ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.subb ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.subc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2 ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3 ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.ram ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rd ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.src1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.src2 ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.src3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.b_in ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.des ;
  wire \oc8051_top_1.oc8051_comp1.eq ;
  wire \oc8051_top_1.oc8051_comp1.eq_r ;
  wire [1:0] \oc8051_top_1.oc8051_comp1.sel ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire \oc8051_top_1.oc8051_cy_select1.data_in ;
  wire \oc8051_top_1.oc8051_cy_select1.data_out ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op_o ;
  wire \oc8051_top_1.oc8051_decoder1.bit_addr ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.comp_sel ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.eq ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.mem_wait ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.op1_c ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op_cur ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op_in ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.pc_sel ;
  wire \oc8051_top_1.oc8051_decoder1.pc_wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o ;
  wire \oc8051_top_1.oc8051_decoder1.rd ;
  wire \oc8051_top_1.oc8051_decoder1.rmw ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state_dec ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire \oc8051_top_1.oc8051_decoder1.wr_o ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr_o ;
  wire [1:0] \oc8051_top_1.oc8051_indi_addr1.bank ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.ri_out ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.sel ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.wr_addr ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.alu ;
  wire [1:0] \oc8051_top_1.oc8051_memory_interface1.bank ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_out ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des_acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_rom_sel ;
  wire \oc8051_top_1.oc8051_memory_interface1.iack_i ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_i ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.inc_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.iram_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire \oc8051_top_1.oc8051_memory_interface1.mem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op1 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op1_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op1_out ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_out ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_out ;
  wire [1:0] \oc8051_top_1.oc8051_memory_interface1.op_length ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.pc_wr_sel ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pcs_result ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.pcs_source ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.rd_addr ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.rd_sel ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sp ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sp_w ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.wr_addr ;
  wire \oc8051_top_1.oc8051_memory_interface1.wr_bit_i ;
  wire \oc8051_top_1.oc8051_memory_interface1.wr_bit_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.wr_dat ;
  wire \oc8051_top_1.oc8051_memory_interface1.wr_i ;
  wire \oc8051_top_1.oc8051_memory_interface1.wr_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.wr_o ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.wr_sel ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_data_in ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_data_out ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_en ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_addr ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_addr_m ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire \oc8051_top_1.oc8051_ram_top1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_addr ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_addr_m ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_m ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.adr0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.adr1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.bank_sel ;
  wire \oc8051_top_1.oc8051_sfr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.comp_sel ;
  wire \oc8051_top_1.oc8051_sfr1.comp_wait ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat2 ;
  wire \oc8051_top_1.oc8051_sfr1.desAc ;
  wire \oc8051_top_1.oc8051_sfr1.desOv ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.des_acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire \oc8051_top_1.oc8051_sfr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.acc ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit_acc ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_sfr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_sfr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.cur_lev ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.il0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.il1 ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept_1 ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_l0 ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_l1 ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l0 ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc_cur ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rmw ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.bank_sel ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_psw ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_rd_sel ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_t ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.write ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tc0_add ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tc1_add ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.run ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sc_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sc_clk_tr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_sbuf ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.ram_rd_sel ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.ram_wr_sel ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rmw ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sp ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sp_w ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.tf1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.we ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.wr_sfr ;
  wire [2:0] \oc8051_top_1.op1_cur ;
  wire [7:0] \oc8051_top_1.op1_n ;
  wire [7:0] \oc8051_top_1.op2_n ;
  wire [7:0] \oc8051_top_1.op3_n ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire \oc8051_top_1.pc_wr ;
  wire [2:0] \oc8051_top_1.pc_wr_sel ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire [7:0] \oc8051_top_1.ram_out ;
  wire [2:0] \oc8051_top_1.ram_rd_sel ;
  wire [2:0] \oc8051_top_1.ram_wr_sel ;
  wire \oc8051_top_1.rd ;
  wire [7:0] \oc8051_top_1.rd_addr ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire [7:0] \oc8051_top_1.ri ;
  wire \oc8051_top_1.rmw ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire [7:0] \oc8051_top_1.sp ;
  wire [7:0] \oc8051_top_1.sp_w ;
  wire [7:0] \oc8051_top_1.src1 ;
  wire [7:0] \oc8051_top_1.src2 ;
  wire [7:0] \oc8051_top_1.src3 ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire [7:0] \oc8051_top_1.sub_result ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire \oc8051_top_1.wr ;
  wire [7:0] \oc8051_top_1.wr_addr ;
  wire [7:0] \oc8051_top_1.wr_dat ;
  wire \oc8051_top_1.wr_ind ;
  wire \oc8051_top_1.wr_o ;
  wire [1:0] \oc8051_top_1.wr_sfr ;
  wire [7:0] op_out;
  wire op_valid;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pcp1;
  wire pcp2;
  wire pcp3;
  output property_invalid;
  wire property_invalid_pcp1;
  wire property_invalid_pcp2;
  wire property_invalid_pcp3;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  nand (_18557_, _14799_, _13651_);
  nand (_18558_, _13653_, _28364_);
  nand (_28366_, _18558_, _18557_);
  nand (_18559_, _14802_, _13651_);
  nand (_18560_, _13653_, _28368_);
  nand (_28370_, _18560_, _18559_);
  nand (_18561_, _14805_, _13651_);
  nand (_18562_, _13653_, _28372_);
  nand (_28374_, _18562_, _18561_);
  nand (_18563_, _14808_, _13651_);
  nand (_18564_, _13653_, _28376_);
  nand (_28378_, _18564_, _18563_);
  nand (_18565_, _13642_, _14789_);
  nand (_18566_, _13644_, _28380_);
  nand (_28382_, _18566_, _18565_);
  nand (_18567_, _14792_, _13642_);
  nand (_18568_, _13644_, _28384_);
  nand (_28386_, _18568_, _18567_);
  nand (_18569_, _14795_, _13642_);
  nand (_18570_, _13644_, _28388_);
  nand (_28390_, _18570_, _18569_);
  nand (_18571_, _14799_, _13642_);
  nand (_18572_, _13644_, _28392_);
  nand (_28394_, _18572_, _18571_);
  nand (_18574_, _14802_, _13642_);
  nand (_18575_, _13644_, _28396_);
  nand (_28398_, _18575_, _18574_);
  nand (_18576_, _14805_, _13642_);
  nand (_18577_, _13644_, _28400_);
  nand (_28402_, _18577_, _18576_);
  nand (_18578_, _14808_, _13642_);
  nand (_18579_, _13644_, _28404_);
  nand (_28406_, _18579_, _18578_);
  nor (_18581_, _13619_, _28408_);
  nor (_28410_, _18581_, _00914_);
  nor (_18582_, _13619_, _28412_);
  nor (_28414_, _18582_, _00911_);
  nor (_18583_, _13619_, _28416_);
  nor (_28418_, _18583_, _00907_);
  nor (_18584_, _13619_, _28420_);
  nor (_28422_, _18584_, _00903_);
  nor (_18585_, _13619_, _28424_);
  nor (_28426_, _18585_, _00899_);
  nor (_18586_, _13619_, _28428_);
  nor (_28430_, _18586_, _00896_);
  nor (_18587_, _13619_, _28433_);
  nor (_28435_, _18587_, _00892_);
  nand (_18588_, _14805_, _13780_);
  nand (_18589_, _13782_, _28437_);
  nand (_28439_, _18589_, _18588_);
  nand (_18590_, _14802_, _13780_);
  nand (_18591_, _13782_, _28441_);
  nand (_28443_, _18591_, _18590_);
  nand (_18592_, _14799_, _13780_);
  nand (_18593_, _13782_, _28445_);
  nand (_28447_, _18593_, _18592_);
  nand (_18594_, _14808_, _13780_);
  nand (_18595_, _13782_, _28449_);
  nand (_28451_, _18595_, _18594_);
  nand (_18596_, _14795_, _13780_);
  nand (_18597_, _13782_, _28453_);
  nand (_28455_, _18597_, _18596_);
  nand (_18598_, _14792_, _13780_);
  nand (_18600_, _13782_, _28457_);
  nand (_28459_, _18600_, _18598_);
  nand (_18601_, _25613_, _03355_);
  nor (_18602_, _18601_, _28271_);
  not (_18603_, _04466_);
  not (_18604_, _18601_);
  nor (_18605_, _18604_, _18603_);
  nor (_18606_, _18605_, _18602_);
  nor (_04469_, _18606_, _23698_);
  nor (_18607_, _18601_, _18603_);
  not (_18609_, _04471_);
  nor (_18610_, _18604_, _18609_);
  nor (_18611_, _18610_, _18607_);
  nor (_04473_, _18611_, _23698_);
  nand (_18612_, _13780_, _14789_);
  nand (_18613_, _13782_, _29296_);
  nand (_04678_, _18613_, _18612_);
  nor (_18614_, _18601_, _27231_);
  not (_18615_, _05028_);
  nor (_18616_, _18604_, _18615_);
  nor (_18617_, _18616_, _18614_);
  nor (_05072_, _18617_, _23698_);
  nor (_18618_, _18601_, _27281_);
  not (_18619_, _05031_);
  nor (_18620_, _18604_, _18619_);
  nor (_18621_, _18620_, _18618_);
  nor (_05074_, _18621_, _23698_);
  nor (_18622_, _18601_, _28503_);
  not (_18623_, _05034_);
  nor (_18624_, _18604_, _18623_);
  nor (_18625_, _18624_, _18622_);
  nor (_05076_, _18625_, _23698_);
  nor (_18626_, _18601_, _27364_);
  not (_18627_, _05036_);
  nor (_18628_, _18604_, _18627_);
  nor (_18629_, _18628_, _18626_);
  nor (_05078_, _18629_, _23698_);
  nor (_18630_, _18601_, _26929_);
  not (_18631_, _05040_);
  nor (_18632_, _18604_, _18631_);
  nor (_18634_, _18632_, _18630_);
  nor (_05079_, _18634_, _23698_);
  nor (_18635_, _18601_, _28347_);
  not (_18636_, _05043_);
  nor (_18637_, _18604_, _18636_);
  nor (_18638_, _18637_, _18635_);
  nor (_05081_, _18638_, _23698_);
  nor (_18639_, _18601_, _28407_);
  not (_18640_, _05046_);
  nor (_18641_, _18604_, _18640_);
  nor (_18643_, _18641_, _18639_);
  nor (_05083_, _18643_, _23698_);
  nor (_18644_, _18601_, _28266_);
  not (_18645_, _05048_);
  nor (_18646_, _18604_, _18645_);
  nor (_18647_, _18646_, _18644_);
  nor (_05085_, _18647_, _23698_);
  nor (_18648_, _18601_, _27227_);
  not (_18649_, _05051_);
  nor (_18650_, _18604_, _18649_);
  nor (_18651_, _18650_, _18648_);
  nor (_05087_, _18651_, _23698_);
  nor (_18652_, _18601_, _27306_);
  not (_18653_, _05054_);
  nor (_18654_, _18604_, _18653_);
  nor (_18655_, _18654_, _18652_);
  nor (_05089_, _18655_, _23698_);
  nor (_18656_, _18601_, _27346_);
  not (_18657_, _05057_);
  nor (_18658_, _18604_, _18657_);
  nor (_18659_, _18658_, _18656_);
  nor (_05091_, _18659_, _23698_);
  nor (_18660_, _18601_, _27368_);
  not (_18661_, _05060_);
  nor (_18662_, _18604_, _18661_);
  nor (_18663_, _18662_, _18660_);
  nor (_05093_, _18663_, _23698_);
  nor (_18664_, _18601_, _26939_);
  not (_18665_, _05063_);
  nor (_18666_, _18604_, _18665_);
  nor (_18668_, _18666_, _18664_);
  nor (_05095_, _18668_, _23698_);
  nor (_18669_, _18601_, _28353_);
  not (_18670_, _05066_);
  nor (_18671_, _18604_, _18670_);
  nor (_18672_, _18671_, _18669_);
  nor (_05097_, _18672_, _23698_);
  nor (_18673_, _18601_, _28411_);
  not (_18674_, _05069_);
  nor (_18675_, _18604_, _18674_);
  nor (_18677_, _18675_, _18673_);
  nor (_05099_, _18677_, _23698_);
  nor (_18678_, _18601_, _18615_);
  not (_18679_, _05101_);
  nor (_18680_, _18604_, _18679_);
  nor (_18681_, _18680_, _18678_);
  nor (_05145_, _18681_, _23698_);
  nor (_18682_, _18601_, _18619_);
  not (_18683_, _05104_);
  nor (_18684_, _18604_, _18683_);
  nor (_18685_, _18684_, _18682_);
  nor (_05147_, _18685_, _23698_);
  nor (_18686_, _18601_, _18623_);
  not (_18687_, _05107_);
  nor (_18688_, _18604_, _18687_);
  nor (_18689_, _18688_, _18686_);
  nor (_05149_, _18689_, _23698_);
  nor (_18690_, _18601_, _18627_);
  not (_18691_, _05110_);
  nor (_18692_, _18604_, _18691_);
  nor (_18693_, _18692_, _18690_);
  nor (_05151_, _18693_, _23698_);
  nor (_18694_, _18601_, _18631_);
  not (_18695_, _05112_);
  nor (_18696_, _18604_, _18695_);
  nor (_18697_, _18696_, _18694_);
  nor (_05153_, _18697_, _23698_);
  nor (_18698_, _18601_, _18636_);
  not (_18699_, _05115_);
  nor (_18700_, _18604_, _18699_);
  nor (_18702_, _18700_, _18698_);
  nor (_05155_, _18702_, _23698_);
  nor (_18703_, _18601_, _18640_);
  not (_18704_, _05118_);
  nor (_18705_, _18604_, _18704_);
  nor (_18706_, _18705_, _18703_);
  nor (_05157_, _18706_, _23698_);
  nor (_18707_, _18601_, _18645_);
  not (_18708_, _05121_);
  nor (_18709_, _18604_, _18708_);
  nor (_18711_, _18709_, _18707_);
  nor (_05159_, _18711_, _23698_);
  nor (_18712_, _18601_, _18649_);
  not (_18713_, _05124_);
  nor (_18714_, _18604_, _18713_);
  nor (_18715_, _18714_, _18712_);
  nor (_05161_, _18715_, _23698_);
  nor (_18716_, _18601_, _18653_);
  not (_18717_, _05127_);
  nor (_18718_, _18604_, _18717_);
  nor (_18719_, _18718_, _18716_);
  nor (_05163_, _18719_, _23698_);
  nor (_18720_, _18601_, _18657_);
  not (_18721_, _05130_);
  nor (_18722_, _18604_, _18721_);
  nor (_18723_, _18722_, _18720_);
  nor (_05165_, _18723_, _23698_);
  nor (_18724_, _18601_, _18661_);
  not (_18725_, _05133_);
  nor (_18726_, _18604_, _18725_);
  nor (_18727_, _18726_, _18724_);
  nor (_05167_, _18727_, _23698_);
  nor (_18728_, _18601_, _18665_);
  not (_18729_, _05136_);
  nor (_18730_, _18604_, _18729_);
  nor (_18731_, _18730_, _18728_);
  nor (_05170_, _18731_, _23698_);
  nor (_18732_, _18601_, _18670_);
  not (_18733_, _05139_);
  nor (_18734_, _18604_, _18733_);
  nor (_18736_, _18734_, _18732_);
  nor (_05172_, _18736_, _23698_);
  nor (_18737_, _18601_, _18674_);
  not (_18738_, _05142_);
  nor (_18739_, _18604_, _18738_);
  nor (_18740_, _18739_, _18737_);
  nor (_05174_, _18740_, _23698_);
  nor (_18741_, _04680_, _30316_);
  nor (_18742_, _04682_, _02518_);
  nor (_18743_, _18742_, _18741_);
  nor (_18745_, _04684_, _30316_);
  nor (_18746_, _04686_, _02518_);
  nor (_18747_, _18746_, _18745_);
  nor (_18748_, _02453_, _30316_);
  nor (_18749_, _04689_, _02518_);
  nor (_18750_, _18749_, _18748_);
  not (_18751_, _18750_);
  nor (_18752_, _02448_, _30316_);
  nor (_18753_, _04693_, _02518_);
  nor (_18754_, _18753_, _18752_);
  not (_18755_, _18754_);
  nor (_18756_, _18755_, _07880_);
  nor (_18757_, _18754_, _07817_);
  nor (_18758_, _18757_, _18756_);
  not (_18759_, _18758_);
  nor (_18760_, _18759_, _18751_);
  not (_18761_, _07679_);
  nor (_18762_, _18754_, _18750_);
  not (_18763_, _18762_);
  nor (_18764_, _18763_, _18761_);
  not (_18765_, _07731_);
  nor (_18766_, _18755_, _18750_);
  not (_18767_, _18766_);
  nor (_18768_, _18767_, _18765_);
  nor (_18769_, _18768_, _18764_);
  not (_18770_, _18769_);
  nor (_18771_, _18770_, _18760_);
  nor (_18772_, _18771_, _18747_);
  nor (_18773_, _18754_, _07743_);
  not (_18774_, _18747_);
  nor (_18776_, _18750_, _18774_);
  not (_18777_, _18776_);
  nor (_18778_, _18755_, _07546_);
  nor (_18779_, _18778_, _18777_);
  not (_18780_, _18779_);
  nor (_18781_, _18780_, _18773_);
  nor (_18782_, _18751_, _18774_);
  not (_18783_, _18782_);
  nor (_18784_, _18755_, _07902_);
  nor (_18785_, _18754_, _07915_);
  nor (_18787_, _18785_, _18784_);
  not (_18788_, _18787_);
  nor (_18789_, _18788_, _18783_);
  nor (_18790_, _18789_, _18781_);
  not (_18791_, _18790_);
  nor (_18792_, _18791_, _18772_);
  nand (_18793_, _18792_, _18743_);
  not (_18794_, _18743_);
  nor (_18795_, _18755_, _07726_);
  nor (_18796_, _18754_, _07780_);
  nor (_18797_, _18796_, _18795_);
  not (_18798_, _18797_);
  nor (_18799_, _18798_, _18751_);
  not (_18800_, _07658_);
  nor (_18801_, _18763_, _18800_);
  not (_18802_, _07638_);
  nor (_18803_, _18767_, _18802_);
  nor (_18804_, _18803_, _18801_);
  not (_18805_, _18804_);
  nor (_18806_, _18805_, _18799_);
  nor (_18807_, _18806_, _18747_);
  nor (_18808_, _18755_, _07835_);
  nor (_18809_, _18754_, _07708_);
  nor (_18810_, _18809_, _18777_);
  not (_18811_, _18810_);
  nor (_18812_, _18811_, _18808_);
  nor (_18813_, _18755_, _07690_);
  nor (_18814_, _18754_, _07863_);
  nor (_18815_, _18814_, _18813_);
  not (_18816_, _18815_);
  nor (_18818_, _18816_, _18783_);
  nor (_18819_, _18818_, _18812_);
  not (_18820_, _18819_);
  nor (_18821_, _18820_, _18807_);
  nand (_18822_, _18821_, _18794_);
  nand (_18823_, _18822_, _18793_);
  not (_18824_, _18823_);
  nor (_18825_, _18794_, _08008_);
  nor (_18826_, _18743_, _08006_);
  nor (_18827_, _18826_, _18825_);
  nor (_18829_, _18827_, _18747_);
  nor (_18830_, _18794_, _08012_);
  nor (_18831_, _18743_, _08010_);
  nor (_18832_, _18831_, _18830_);
  nor (_18833_, _18832_, _18774_);
  nor (_18834_, _18833_, _18829_);
  nand (_18835_, _18834_, _18751_);
  nor (_18836_, _18751_, _18747_);
  nor (_18837_, _18794_, _08016_);
  nor (_18838_, _18743_, _08014_);
  nor (_18839_, _18838_, _18837_);
  nand (_18840_, _18839_, _18836_);
  nand (_18841_, _18840_, _18835_);
  nand (_18842_, _18841_, _18755_);
  not (_18843_, _08037_);
  nand (_18844_, _18743_, _18843_);
  not (_18845_, _08035_);
  nand (_18846_, _18794_, _18845_);
  nand (_18847_, _18846_, _18844_);
  nor (_18848_, _18847_, _18783_);
  not (_18849_, _18836_);
  not (_18850_, _08033_);
  nand (_18851_, _18743_, _18850_);
  not (_18852_, _08031_);
  nand (_18853_, _18794_, _18852_);
  nand (_18854_, _18853_, _18851_);
  nor (_18855_, _18854_, _18849_);
  nor (_18856_, _18855_, _18848_);
  nor (_18857_, _18856_, _18755_);
  nor (_18858_, _18794_, _08020_);
  nor (_18860_, _18743_, _08018_);
  nor (_18861_, _18860_, _18858_);
  nor (_18862_, _18783_, _18754_);
  nand (_18863_, _18862_, _18861_);
  nor (_18864_, _18794_, _08029_);
  nor (_18865_, _18743_, _08027_);
  nor (_18866_, _18865_, _18864_);
  nand (_18867_, _18866_, _18747_);
  nor (_18868_, _18794_, _08025_);
  nor (_18869_, _18743_, _08022_);
  nor (_18871_, _18869_, _18868_);
  nand (_18872_, _18871_, _18774_);
  nand (_18873_, _18872_, _18867_);
  nand (_18874_, _18873_, _18766_);
  nand (_18875_, _18874_, _18863_);
  nor (_18876_, _18875_, _18857_);
  nand (_18877_, _18876_, _18842_);
  nand (_18878_, _18877_, _18824_);
  nand (_18879_, _18823_, _07539_);
  nand (_07543_, _18879_, _18878_);
  nor (_18880_, _18794_, _18747_);
  not (_18881_, _18880_);
  nor (_18882_, _18794_, _18774_);
  not (_18883_, _18882_);
  nor (_18884_, _18883_, _18751_);
  nor (_18885_, _18882_, _18750_);
  nor (_18886_, _18885_, _18884_);
  not (_18887_, _07708_);
  not (_18888_, _18884_);
  nor (_18889_, _18888_, _18755_);
  nor (_18890_, _18884_, _18754_);
  nor (_18891_, _18890_, _18889_);
  nor (_18892_, _18891_, _18887_);
  not (_18893_, _07835_);
  not (_18894_, _18891_);
  nor (_18895_, _18894_, _18893_);
  nor (_18896_, _18895_, _18892_);
  nor (_18897_, _18896_, _18886_);
  not (_18898_, _18886_);
  not (_18899_, _07863_);
  nor (_18901_, _18891_, _18899_);
  not (_18902_, _07690_);
  nor (_18903_, _18894_, _18902_);
  nor (_18904_, _18903_, _18901_);
  nor (_18905_, _18904_, _18898_);
  nor (_18906_, _18905_, _18897_);
  nor (_18907_, _18906_, _18881_);
  nor (_18908_, _18743_, _18774_);
  not (_18909_, _18908_);
  not (_18910_, _07743_);
  nor (_18913_, _18891_, _18910_);
  not (_18914_, _07546_);
  nor (_18915_, _18894_, _18914_);
  nor (_18916_, _18915_, _18913_);
  nor (_18917_, _18916_, _18886_);
  not (_18918_, _07915_);
  nor (_18919_, _18891_, _18918_);
  not (_18920_, _07902_);
  nor (_18921_, _18894_, _18920_);
  nor (_18922_, _18921_, _18919_);
  nor (_18923_, _18922_, _18898_);
  nor (_18924_, _18923_, _18917_);
  nor (_18925_, _18924_, _18909_);
  nor (_18926_, _18925_, _18907_);
  nor (_18927_, _18891_, _18800_);
  nor (_18928_, _18894_, _18802_);
  nor (_18929_, _18928_, _18927_);
  nor (_18930_, _18929_, _18886_);
  not (_18931_, _07780_);
  nor (_18932_, _18891_, _18931_);
  not (_18933_, _07726_);
  nor (_18934_, _18894_, _18933_);
  nor (_18935_, _18934_, _18932_);
  nor (_18936_, _18935_, _18898_);
  nor (_18937_, _18936_, _18930_);
  nor (_18938_, _18937_, _18883_);
  nor (_18939_, _18743_, _18747_);
  not (_18940_, _18939_);
  nor (_18941_, _18891_, _18761_);
  nor (_18942_, _18894_, _18765_);
  nor (_18944_, _18942_, _18941_);
  nor (_18945_, _18944_, _18886_);
  not (_18946_, _07817_);
  nor (_18947_, _18891_, _18946_);
  not (_18948_, _07880_);
  nor (_18949_, _18894_, _18948_);
  nor (_18950_, _18949_, _18947_);
  nor (_18951_, _18950_, _18898_);
  nor (_18952_, _18951_, _18945_);
  nor (_18953_, _18952_, _18940_);
  nor (_18955_, _18953_, _18938_);
  nand (_18956_, _18955_, _18926_);
  nor (_18957_, _18908_, _18880_);
  nor (_18958_, _18794_, _08022_);
  nor (_18959_, _18743_, _08025_);
  nor (_18960_, _18959_, _18958_);
  nand (_18961_, _18960_, _18957_);
  not (_18962_, _18957_);
  nor (_18963_, _18794_, _08027_);
  nor (_18964_, _18743_, _08029_);
  nor (_18965_, _18964_, _18963_);
  nand (_18966_, _18965_, _18962_);
  nand (_18967_, _18966_, _18961_);
  nand (_18968_, _18967_, _18898_);
  nor (_18969_, _18794_, _08031_);
  nor (_18970_, _18743_, _08033_);
  nor (_18971_, _18970_, _18969_);
  nand (_18972_, _18971_, _18957_);
  nor (_18973_, _18794_, _08035_);
  nor (_18974_, _18743_, _08037_);
  nor (_18975_, _18974_, _18973_);
  nand (_18976_, _18975_, _18962_);
  nand (_18977_, _18976_, _18972_);
  nand (_18978_, _18977_, _18886_);
  nand (_18979_, _18978_, _18968_);
  nand (_18980_, _18979_, _18891_);
  nor (_18981_, _18794_, _08006_);
  nor (_18982_, _18743_, _08008_);
  nor (_18983_, _18982_, _18981_);
  nand (_18984_, _18983_, _18957_);
  nor (_18986_, _18794_, _08010_);
  nor (_18987_, _18743_, _08012_);
  nor (_18988_, _18987_, _18986_);
  nand (_18989_, _18988_, _18962_);
  nand (_18990_, _18989_, _18984_);
  nand (_18991_, _18990_, _18898_);
  nor (_18992_, _18794_, _08014_);
  nor (_18993_, _18743_, _08016_);
  nor (_18994_, _18993_, _18992_);
  nand (_18995_, _18994_, _18957_);
  nor (_18997_, _18794_, _08018_);
  nor (_18998_, _18743_, _08020_);
  nor (_18999_, _18998_, _18997_);
  nand (_19000_, _18999_, _18962_);
  nand (_19001_, _19000_, _18995_);
  nand (_19002_, _19001_, _18886_);
  nand (_19003_, _19002_, _18991_);
  nand (_19004_, _19003_, _18894_);
  nand (_19005_, _19004_, _18980_);
  nand (_19006_, _19005_, _18956_);
  not (_19007_, _18956_);
  nand (_19008_, _19007_, _07549_);
  nand (_07552_, _19008_, _19006_);
  nor (_19009_, _18782_, _18755_);
  nor (_19010_, _19009_, _18862_);
  not (_19011_, _19010_);
  nor (_19012_, _19011_, _07780_);
  nor (_19013_, _18836_, _18776_);
  nor (_19014_, _19013_, _18795_);
  not (_19015_, _19014_);
  nor (_19016_, _19015_, _19012_);
  not (_19017_, _19013_);
  nor (_19018_, _19017_, _19011_);
  not (_19019_, _19018_);
  nor (_19020_, _19019_, _18800_);
  nor (_19021_, _19017_, _19010_);
  not (_19022_, _19021_);
  nor (_19023_, _19022_, _18802_);
  nor (_19024_, _19023_, _19020_);
  not (_19025_, _19024_);
  nor (_19027_, _19025_, _19016_);
  nor (_19028_, _19027_, _18909_);
  nor (_19029_, _18883_, _18750_);
  nor (_19030_, _19010_, _07880_);
  nor (_19031_, _19011_, _07817_);
  nor (_19032_, _19031_, _19030_);
  nand (_19033_, _19032_, _19029_);
  not (_19034_, _19033_);
  nor (_19035_, _19022_, _18765_);
  nor (_19036_, _19019_, _18761_);
  nor (_19038_, _19036_, _19035_);
  nor (_19039_, _19038_, _18883_);
  nor (_19040_, _19039_, _19034_);
  not (_19041_, _19040_);
  nor (_19042_, _19041_, _19028_);
  nor (_19043_, _19011_, _07863_);
  nor (_19044_, _19013_, _18813_);
  not (_19045_, _19044_);
  nor (_19046_, _19045_, _19043_);
  nor (_19047_, _19019_, _18887_);
  nor (_19048_, _19022_, _18893_);
  nor (_19049_, _19048_, _19047_);
  not (_19050_, _19049_);
  nor (_19051_, _19050_, _19046_);
  nor (_19052_, _19051_, _18940_);
  nor (_19053_, _19011_, _07915_);
  nor (_19054_, _19013_, _18784_);
  not (_19055_, _19054_);
  nor (_19056_, _19055_, _19053_);
  nor (_19057_, _19022_, _18914_);
  nor (_19058_, _19019_, _18910_);
  nor (_19059_, _19058_, _19057_);
  not (_19060_, _19059_);
  nor (_19061_, _19060_, _19056_);
  nor (_19062_, _19061_, _18881_);
  nor (_19063_, _19062_, _19052_);
  nand (_19064_, _19063_, _19042_);
  nor (_19065_, _18832_, _18747_);
  nor (_19066_, _18827_, _18774_);
  nor (_19067_, _19066_, _19065_);
  nand (_19069_, _19067_, _19013_);
  nand (_19070_, _18839_, _18747_);
  nand (_19071_, _18861_, _18774_);
  nand (_19072_, _19071_, _19070_);
  nand (_19073_, _19072_, _19017_);
  nand (_19074_, _19073_, _19069_);
  nand (_19075_, _19074_, _19010_);
  nor (_19076_, _18866_, _18747_);
  nor (_19077_, _18871_, _18774_);
  nor (_19078_, _19077_, _19076_);
  nand (_19080_, _19078_, _19013_);
  nor (_19081_, _18847_, _18849_);
  nor (_19082_, _18854_, _18777_);
  nor (_19083_, _19082_, _19081_);
  nand (_19084_, _19083_, _19080_);
  nand (_19085_, _19084_, _19011_);
  nand (_19086_, _19085_, _19075_);
  nand (_19087_, _19086_, _19064_);
  not (_19088_, _19064_);
  nand (_19089_, _19088_, _07558_);
  nand (_07561_, _19089_, _19087_);
  nor (_19090_, _18939_, _18751_);
  nor (_19091_, _18940_, _18750_);
  nor (_19092_, _19091_, _19090_);
  not (_19093_, _19090_);
  nor (_19094_, _19093_, _18754_);
  nor (_19095_, _19090_, _18755_);
  nor (_19096_, _19095_, _19094_);
  not (_19097_, _19096_);
  nor (_19098_, _19097_, _19092_);
  not (_19099_, _19098_);
  nor (_19100_, _19099_, _18761_);
  not (_19101_, _19092_);
  nor (_19102_, _19101_, _18759_);
  nor (_19103_, _19096_, _19092_);
  not (_19104_, _19103_);
  nor (_19105_, _19104_, _18765_);
  nor (_19106_, _19105_, _19102_);
  not (_19107_, _19106_);
  nor (_19108_, _19107_, _19100_);
  nor (_19110_, _19108_, _18909_);
  nor (_19111_, _19104_, _18914_);
  nor (_19112_, _19101_, _18788_);
  nor (_19113_, _19099_, _18910_);
  nor (_19114_, _19113_, _19112_);
  not (_19115_, _19114_);
  nor (_19116_, _19115_, _19111_);
  nor (_19117_, _19116_, _18940_);
  nor (_19118_, _19117_, _19110_);
  nor (_19119_, _19104_, _18802_);
  nor (_19121_, _19101_, _18798_);
  nor (_19122_, _19099_, _18800_);
  nor (_19123_, _19122_, _19121_);
  not (_19124_, _19123_);
  nor (_19125_, _19124_, _19119_);
  nor (_19126_, _19125_, _18881_);
  nor (_19127_, _19099_, _18887_);
  nor (_19128_, _19101_, _18816_);
  nor (_19129_, _19104_, _18893_);
  nor (_19130_, _19129_, _19128_);
  not (_19131_, _19130_);
  nor (_19132_, _19131_, _19127_);
  nor (_19133_, _19132_, _18883_);
  nor (_19134_, _19133_, _19126_);
  nand (_19135_, _19134_, _19118_);
  nand (_19136_, _18971_, _18962_);
  nand (_19137_, _18975_, _18957_);
  nand (_19138_, _19137_, _19136_);
  nor (_19139_, _19101_, _18755_);
  nand (_19140_, _19139_, _19138_);
  not (_19141_, _18960_);
  nor (_19142_, _19141_, _18957_);
  not (_19143_, _18965_);
  nor (_19144_, _19143_, _18962_);
  nor (_19145_, _19144_, _19142_);
  nor (_19146_, _19145_, _19104_);
  nand (_19147_, _18983_, _18962_);
  nand (_19148_, _18988_, _18957_);
  nand (_19149_, _19148_, _19147_);
  nand (_19150_, _19149_, _19098_);
  nand (_19151_, _18994_, _18962_);
  nand (_19152_, _18999_, _18957_);
  nand (_19153_, _19152_, _19151_);
  nor (_19154_, _19101_, _18754_);
  nand (_19155_, _19154_, _19153_);
  nand (_19156_, _19155_, _19150_);
  nor (_19157_, _19156_, _19146_);
  nand (_19158_, _19157_, _19140_);
  nand (_19159_, _19158_, _19135_);
  not (_19160_, _19135_);
  nand (_19162_, _19160_, _07569_);
  nand (_07572_, _19162_, _19159_);
  nor (_19163_, _19135_, _23698_);
  not (_19164_, _19163_);
  nor (_19165_, _19164_, _19101_);
  not (_19166_, _19165_);
  nor (_19167_, _19166_, _19096_);
  not (_19168_, _19167_);
  nor (_19169_, _19168_, _18940_);
  not (_19170_, _19169_);
  nor (_19172_, _19064_, _23698_);
  not (_19173_, _19172_);
  nor (_19174_, _19173_, _19013_);
  not (_19175_, _19174_);
  nor (_19176_, _19175_, _19010_);
  not (_19177_, _19176_);
  nor (_19178_, _19177_, _18881_);
  not (_19179_, _19178_);
  nor (_19180_, _18793_, _23698_);
  not (_19181_, _19180_);
  nor (_19182_, _19181_, _18774_);
  not (_19183_, _19182_);
  nor (_19184_, _18824_, _23698_);
  not (_19185_, _19184_);
  nand (_19186_, _18754_, _18750_);
  nor (_19187_, _19186_, _19185_);
  not (_19188_, _19187_);
  nor (_19189_, _19188_, _19183_);
  nor (_19190_, _18879_, _23698_);
  not (_19191_, _19190_);
  nand (_19192_, _19191_, _19189_);
  nor (_19193_, _18956_, _23698_);
  not (_19194_, _19193_);
  nor (_19195_, _19194_, _18894_);
  not (_19196_, _19195_);
  nor (_19197_, _19196_, _18898_);
  not (_19198_, _19197_);
  nor (_19199_, _19198_, _18909_);
  nor (_19200_, _19189_, _08037_);
  nor (_19201_, _19200_, _19199_);
  nand (_19203_, _19201_, _19192_);
  not (_19204_, _07549_);
  nor (_19205_, _19194_, _19204_);
  nand (_19206_, _19205_, _19199_);
  nand (_19207_, _19206_, _19203_);
  nand (_19208_, _19207_, _19179_);
  nor (_19209_, _19089_, _23698_);
  nand (_19210_, _19209_, _19178_);
  nand (_19211_, _19210_, _19208_);
  nand (_19212_, _19211_, _19170_);
  nor (_19214_, _19162_, _23698_);
  nand (_19215_, _19214_, _19169_);
  nand (_07650_, _19215_, _19212_);
  nor (_19216_, _19099_, _18881_);
  not (_19217_, _19216_);
  nor (_19218_, _18940_, _18763_);
  nor (_19219_, _19218_, _07658_);
  nand (_19220_, _19219_, _19217_);
  nor (_19221_, _18783_, _18755_);
  nor (_19222_, _19221_, _19220_);
  nor (_07676_, _19222_, _23698_);
  nor (_19223_, _19013_, _19010_);
  nor (_19224_, _19223_, _07880_);
  nor (_07683_, _19224_, _23698_);
  nand (_19225_, _18762_, _18774_);
  nand (_19226_, _19225_, _18761_);
  nor (_19227_, _19226_, _19221_);
  nor (_07704_, _19227_, _23698_);
  nor (_19228_, _18766_, _07546_);
  nor (_07718_, _19228_, _23698_);
  nor (_19229_, _19103_, _07638_);
  nor (_07724_, _19229_, _23698_);
  nor (_19230_, _18882_, _18763_);
  not (_19231_, _18889_);
  nand (_19232_, _19231_, _18887_);
  nor (_19233_, _19232_, _19230_);
  nor (_07740_, _19233_, _23698_);
  nor (_19234_, _18762_, _07743_);
  nor (_07777_, _19234_, _23698_);
  nor (_19235_, _19019_, _18909_);
  not (_19237_, _19235_);
  nor (_19238_, _18940_, _18751_);
  nand (_19239_, _19238_, _18754_);
  nand (_19240_, _19239_, _19237_);
  nor (_19241_, _18889_, _07902_);
  nand (_19242_, _19241_, _19217_);
  nor (_19243_, _19242_, _19240_);
  nor (_07787_, _19243_, _23698_);
  nor (_19244_, _18957_, _18763_);
  nand (_19245_, _18882_, _18762_);
  nor (_19247_, _18754_, _18751_);
  not (_19248_, _19247_);
  nor (_19249_, _19248_, _18940_);
  nor (_19250_, _19249_, _07780_);
  nand (_19251_, _19250_, _19245_);
  nor (_19252_, _19251_, _19244_);
  nor (_07814_, _19252_, _23698_);
  nand (_19253_, _18766_, _18774_);
  nand (_19254_, _19253_, _18765_);
  nor (_19255_, _19254_, _18862_);
  nor (_07832_, _19255_, _23698_);
  nor (_19256_, _19104_, _18881_);
  not (_19257_, _19249_);
  nor (_19258_, _18777_, _18754_);
  nor (_19259_, _19258_, _07817_);
  nand (_19260_, _19259_, _19257_);
  nor (_19261_, _19260_, _19256_);
  nor (_07860_, _19261_, _23698_);
  nor (_19262_, _18883_, _18767_);
  not (_19263_, _19262_);
  nand (_19264_, _19239_, _19263_);
  nand (_19265_, _18962_, _18766_);
  nand (_19266_, _19265_, _18933_);
  nor (_19267_, _19266_, _19264_);
  nor (_07873_, _19267_, _23698_);
  nor (_19268_, _18862_, _07915_);
  nand (_19269_, _19268_, _19257_);
  nor (_19270_, _19269_, _19256_);
  nor (_07878_, _19270_, _23698_);
  nor (_19271_, _19264_, _07690_);
  nand (_19273_, _19271_, _19217_);
  nor (_19274_, _19273_, _19235_);
  nor (_07897_, _19274_, _23698_);
  nand (_19275_, _19247_, _18962_);
  nand (_19276_, _19275_, _18899_);
  nand (_19277_, _19257_, _19245_);
  nor (_19278_, _19277_, _19276_);
  nor (_07911_, _19278_, _23698_);
  nor (_19279_, _18882_, _18767_);
  nand (_19280_, _18884_, _18755_);
  nand (_19282_, _19280_, _18893_);
  nor (_19283_, _19282_, _19279_);
  nor (_07929_, _19283_, _23698_);
  nor (_19284_, _19217_, _19164_);
  not (_19285_, _19284_);
  nor (_19286_, _19237_, _19173_);
  not (_19287_, _19286_);
  nor (_19288_, _19194_, _18898_);
  nor (_19289_, _19288_, _19195_);
  not (_19290_, _19289_);
  nor (_19291_, _19290_, _18883_);
  nand (_19292_, _19291_, _19193_);
  nor (_19293_, _19185_, _18774_);
  nor (_19294_, _19293_, _19180_);
  not (_19295_, _19294_);
  nor (_19296_, _19295_, _18763_);
  nand (_19297_, _19296_, _19184_);
  nand (_19298_, _19297_, _08006_);
  nand (_19299_, _19296_, _19190_);
  nand (_19300_, _19299_, _19298_);
  nand (_19301_, _19300_, _19292_);
  nand (_19302_, _19291_, _19205_);
  nand (_19303_, _19302_, _19301_);
  nand (_19304_, _19303_, _19287_);
  nand (_19305_, _19286_, _19209_);
  nand (_19306_, _19305_, _19304_);
  nand (_19307_, _19306_, _19285_);
  nand (_19308_, _19284_, _07569_);
  nand (_08109_, _19308_, _19307_);
  nor (_19309_, _19173_, _18883_);
  not (_19312_, _19309_);
  nor (_19313_, _19312_, _19019_);
  not (_19314_, _19313_);
  nor (_19315_, _19194_, _18940_);
  nand (_19316_, _19315_, _19289_);
  not (_19317_, _08008_);
  nand (_19318_, _19184_, _18763_);
  not (_19319_, _19318_);
  nor (_19320_, _19181_, _18747_);
  not (_19321_, _19320_);
  nor (_19323_, _19321_, _19319_);
  not (_19324_, _19323_);
  nand (_19325_, _19324_, _19317_);
  nand (_19326_, _19323_, _19191_);
  nand (_19327_, _19326_, _19325_);
  nand (_19328_, _19327_, _19316_);
  not (_19329_, _19316_);
  nand (_19330_, _19329_, _19204_);
  nand (_19331_, _19330_, _19328_);
  nand (_19332_, _19331_, _19314_);
  nor (_19333_, _19164_, _18909_);
  nand (_19334_, _19333_, _19098_);
  not (_19335_, _19334_);
  nor (_19336_, _19314_, _19209_);
  nor (_19337_, _19336_, _19335_);
  nand (_19338_, _19337_, _19332_);
  nand (_19339_, _19335_, _19214_);
  nand (_08135_, _19339_, _19338_);
  nor (_19340_, _19164_, _18883_);
  not (_19341_, _19340_);
  nor (_19342_, _19341_, _19099_);
  not (_19343_, _19342_);
  nor (_19344_, _19290_, _18881_);
  nand (_19345_, _19344_, _19193_);
  not (_19346_, _19345_);
  nand (_19347_, _19293_, _19181_);
  nor (_19348_, _19347_, _18763_);
  not (_19349_, _19348_);
  nor (_19350_, _19349_, _19191_);
  not (_19351_, _08010_);
  nor (_19353_, _19348_, _19351_);
  nor (_19354_, _19353_, _19350_);
  nor (_19355_, _19354_, _19346_);
  nor (_19356_, _19173_, _18940_);
  not (_19357_, _19356_);
  nor (_19358_, _19357_, _19019_);
  not (_19359_, _19358_);
  nand (_19360_, _19344_, _19205_);
  nand (_19361_, _19360_, _19359_);
  nor (_19362_, _19361_, _19355_);
  nor (_19364_, _19359_, _19209_);
  nor (_19365_, _19364_, _19362_);
  nand (_19366_, _19365_, _19343_);
  nand (_19367_, _19342_, _19214_);
  nand (_08161_, _19367_, _19366_);
  nor (_19368_, _19194_, _18909_);
  nand (_19369_, _19289_, _19368_);
  not (_19370_, _19369_);
  nor (_19371_, _19319_, _19183_);
  not (_19372_, _19371_);
  nand (_19373_, _19372_, _08012_);
  nand (_19374_, _19371_, _19190_);
  nand (_19375_, _19374_, _19373_);
  nor (_19376_, _19375_, _19370_);
  nor (_19377_, _19173_, _18881_);
  not (_19378_, _19377_);
  nor (_19379_, _19378_, _19019_);
  not (_19380_, _19379_);
  nand (_19381_, _19370_, _19204_);
  nand (_19382_, _19381_, _19380_);
  nor (_19383_, _19382_, _19376_);
  nand (_19384_, _19218_, _19163_);
  nand (_19385_, _19379_, _19209_);
  nand (_19386_, _19385_, _19384_);
  nor (_19387_, _19386_, _19383_);
  nor (_19388_, _19384_, _19214_);
  nor (_08178_, _19388_, _19387_);
  nor (_19389_, _19166_, _19097_);
  not (_19390_, _19389_);
  nor (_19391_, _19390_, _18881_);
  nor (_19393_, _19175_, _19011_);
  not (_19394_, _19393_);
  nor (_19395_, _19394_, _18909_);
  not (_19396_, _19395_);
  nor (_19397_, _19396_, _19209_);
  nor (_19398_, _19248_, _19185_);
  not (_19399_, _19398_);
  nor (_19400_, _19399_, _19295_);
  nand (_19401_, _19400_, _19191_);
  nand (_19402_, _19288_, _18894_);
  nor (_19404_, _19402_, _18883_);
  nor (_19405_, _19400_, _08014_);
  nor (_19406_, _19405_, _19404_);
  nand (_19407_, _19406_, _19401_);
  nand (_19408_, _19404_, _19205_);
  nand (_19409_, _19408_, _19407_);
  nor (_19410_, _19409_, _19395_);
  nor (_19411_, _19410_, _19397_);
  nor (_19412_, _19411_, _19391_);
  not (_19413_, _19391_);
  nor (_19414_, _19413_, _19214_);
  nor (_08204_, _19414_, _19412_);
  nor (_19415_, _19390_, _18909_);
  nor (_19416_, _19394_, _18883_);
  nor (_19417_, _19399_, _19321_);
  nand (_19418_, _19417_, _19191_);
  nor (_19419_, _19402_, _18940_);
  nor (_19420_, _19417_, _08016_);
  nor (_19421_, _19420_, _19419_);
  nand (_19422_, _19421_, _19418_);
  nand (_19423_, _19419_, _19205_);
  nand (_19424_, _19423_, _19422_);
  nor (_19425_, _19424_, _19416_);
  not (_19426_, _19416_);
  nor (_19427_, _19426_, _19209_);
  nor (_19428_, _19427_, _19425_);
  nor (_19429_, _19428_, _19415_);
  not (_19430_, _19415_);
  nor (_19431_, _19430_, _19214_);
  nor (_08217_, _19431_, _19429_);
  nor (_19433_, _19390_, _18883_);
  nor (_19434_, _19394_, _18940_);
  not (_19435_, _19434_);
  nor (_19436_, _19435_, _19209_);
  nor (_19437_, _19347_, _19248_);
  nand (_19438_, _19437_, _19191_);
  nor (_19439_, _19402_, _18881_);
  nor (_19440_, _19437_, _08018_);
  nor (_19441_, _19440_, _19439_);
  nand (_19442_, _19441_, _19438_);
  nand (_19444_, _19439_, _19205_);
  nand (_19445_, _19444_, _19442_);
  nor (_19446_, _19445_, _19434_);
  nor (_19447_, _19446_, _19436_);
  nor (_19448_, _19447_, _19433_);
  not (_19449_, _19433_);
  nor (_19450_, _19449_, _19214_);
  nor (_08230_, _19450_, _19448_);
  nor (_19451_, _19390_, _18940_);
  nor (_19452_, _19394_, _18881_);
  nor (_19453_, _19399_, _19183_);
  nand (_19454_, _19453_, _19191_);
  nor (_19455_, _19402_, _18909_);
  nor (_19456_, _19453_, _08020_);
  nor (_19457_, _19456_, _19455_);
  nand (_19458_, _19457_, _19454_);
  nand (_19459_, _19455_, _19205_);
  nand (_19460_, _19459_, _19458_);
  nor (_19461_, _19460_, _19452_);
  not (_19462_, _19452_);
  nor (_19463_, _19462_, _19209_);
  nor (_19464_, _19463_, _19461_);
  nor (_19465_, _19464_, _19451_);
  not (_19466_, _19451_);
  nor (_19467_, _19466_, _19214_);
  nor (_08244_, _19467_, _19465_);
  nand (_19468_, _19256_, _19163_);
  not (_19469_, _18862_);
  nor (_19470_, _19469_, _18743_);
  nand (_19471_, _19470_, _19172_);
  not (_19473_, _19471_);
  nor (_19474_, _19185_, _18767_);
  not (_19475_, _19474_);
  nor (_19476_, _19475_, _19295_);
  nand (_19477_, _19476_, _19191_);
  nor (_19478_, _19196_, _18888_);
  nor (_19479_, _19476_, _08022_);
  nor (_19480_, _19479_, _19478_);
  nand (_19481_, _19480_, _19477_);
  nand (_19482_, _19478_, _19205_);
  nand (_19484_, _19482_, _19481_);
  nor (_19485_, _19484_, _19473_);
  nor (_19486_, _19471_, _07558_);
  nor (_19487_, _19486_, _19485_);
  nand (_19488_, _19487_, _19468_);
  not (_19489_, _19468_);
  nand (_19490_, _19489_, _07569_);
  nand (_08269_, _19490_, _19488_);
  nor (_19491_, _19312_, _19022_);
  nor (_19492_, _19196_, _18886_);
  not (_19493_, _19492_);
  nor (_19494_, _19493_, _18940_);
  not (_19495_, _08025_);
  nor (_19496_, _19475_, _19321_);
  nor (_19497_, _19496_, _19495_);
  not (_19498_, _19496_);
  nor (_19499_, _19498_, _19191_);
  nor (_19500_, _19499_, _19497_);
  nor (_19501_, _19500_, _19494_);
  not (_19502_, _19494_);
  nor (_19503_, _19502_, _19204_);
  nor (_19504_, _19503_, _19501_);
  nor (_19505_, _19504_, _19491_);
  nand (_19506_, _19333_, _19103_);
  nand (_19507_, _19491_, _19209_);
  nand (_19508_, _19507_, _19506_);
  nor (_19509_, _19508_, _19505_);
  nor (_19510_, _19506_, _19214_);
  nor (_08282_, _19510_, _19509_);
  nor (_19511_, _19341_, _19104_);
  not (_19513_, _19511_);
  nor (_19514_, _19493_, _18881_);
  not (_19515_, _08027_);
  nor (_19516_, _19347_, _18767_);
  nor (_19517_, _19516_, _19515_);
  not (_19518_, _19516_);
  nor (_19519_, _19518_, _19191_);
  nor (_19520_, _19519_, _19517_);
  nor (_19521_, _19520_, _19514_);
  nor (_19522_, _19357_, _19022_);
  not (_19524_, _19522_);
  nand (_19525_, _19514_, _19205_);
  nand (_19526_, _19525_, _19524_);
  nor (_19527_, _19526_, _19521_);
  nor (_19528_, _19524_, _19209_);
  nor (_19529_, _19528_, _19527_);
  nand (_19530_, _19529_, _19513_);
  nand (_19531_, _19511_, _19214_);
  nand (_08297_, _19531_, _19530_);
  nor (_19532_, _19493_, _18909_);
  not (_19533_, _19532_);
  nor (_19534_, _19533_, _19205_);
  nor (_19535_, _19378_, _19022_);
  not (_19536_, _19535_);
  not (_19537_, _08029_);
  nor (_19538_, _19475_, _19183_);
  not (_19539_, _19538_);
  nand (_19540_, _19539_, _19537_);
  nand (_19541_, _19538_, _19191_);
  nand (_19542_, _19541_, _19540_);
  nand (_19543_, _19542_, _19533_);
  nand (_19544_, _19543_, _19536_);
  nor (_19545_, _19544_, _19534_);
  nor (_19546_, _19104_, _18940_);
  nand (_19547_, _19546_, _19163_);
  nand (_19548_, _19535_, _19209_);
  nand (_19549_, _19548_, _19547_);
  nor (_19550_, _19549_, _19545_);
  nor (_19551_, _19547_, _07569_);
  nor (_08310_, _19551_, _19550_);
  nor (_19553_, _19168_, _18881_);
  not (_19554_, _19553_);
  nor (_19555_, _19177_, _18909_);
  not (_19556_, _19555_);
  nor (_19557_, _19295_, _19188_);
  nand (_19558_, _19557_, _19191_);
  nor (_19559_, _19263_, _19194_);
  nor (_19560_, _19557_, _08031_);
  nor (_19561_, _19560_, _19559_);
  nand (_19562_, _19561_, _19558_);
  nand (_19564_, _19559_, _19205_);
  nand (_19565_, _19564_, _19562_);
  nand (_19566_, _19565_, _19556_);
  nand (_19567_, _19555_, _19209_);
  nand (_19568_, _19567_, _19566_);
  nand (_19569_, _19568_, _19554_);
  nand (_19570_, _19553_, _19214_);
  nand (_08327_, _19570_, _19569_);
  nor (_19571_, _19168_, _18909_);
  nor (_19572_, _19177_, _18883_);
  nor (_19573_, _19321_, _19188_);
  nand (_19574_, _19573_, _19191_);
  nor (_19575_, _19198_, _18940_);
  nor (_19576_, _19573_, _08033_);
  nor (_19577_, _19576_, _19575_);
  nand (_19578_, _19577_, _19574_);
  nand (_19579_, _19575_, _19205_);
  nand (_19580_, _19579_, _19578_);
  nor (_19581_, _19580_, _19572_);
  not (_19582_, _19572_);
  nor (_19583_, _19582_, _07558_);
  nor (_19584_, _19583_, _19581_);
  nor (_19585_, _19584_, _19571_);
  not (_19586_, _19571_);
  nor (_19587_, _19586_, _19214_);
  nor (_08341_, _19587_, _19585_);
  nor (_19588_, _19168_, _18883_);
  nor (_19589_, _19177_, _18940_);
  nor (_19590_, _19347_, _19188_);
  nand (_19591_, _19590_, _19191_);
  nor (_19593_, _19198_, _18881_);
  nor (_19594_, _19590_, _08035_);
  nor (_19595_, _19594_, _19593_);
  nand (_19596_, _19595_, _19591_);
  nand (_19597_, _19593_, _19205_);
  nand (_19598_, _19597_, _19596_);
  nor (_19599_, _19598_, _19589_);
  not (_19600_, _19589_);
  nor (_19601_, _19600_, _19209_);
  nor (_19602_, _19601_, _19599_);
  nor (_19604_, _19602_, _19588_);
  not (_19605_, _19588_);
  nor (_19606_, _19605_, _19214_);
  nor (_08354_, _19606_, _19604_);
  nand (_19607_, _18823_, _08395_);
  nor (_19608_, _19607_, _23698_);
  not (_19609_, _19608_);
  nand (_19610_, _19609_, _19189_);
  nor (_19611_, _19189_, _08699_);
  nor (_19612_, _19611_, _19199_);
  nand (_19613_, _19612_, _19610_);
  not (_19614_, _08426_);
  nor (_19615_, _19194_, _19614_);
  nand (_19616_, _19615_, _19199_);
  nand (_19617_, _19616_, _19613_);
  nor (_19618_, _19617_, _19178_);
  nand (_19619_, _19088_, _08469_);
  nor (_19620_, _19619_, _23698_);
  nor (_19621_, _19620_, _19179_);
  nor (_19622_, _19621_, _19618_);
  nor (_19623_, _19622_, _19169_);
  nand (_19624_, _19160_, _08520_);
  nor (_19625_, _19624_, _23698_);
  nor (_19626_, _19625_, _19170_);
  nor (_08367_, _19626_, _19623_);
  nand (_19627_, _18823_, _08400_);
  nor (_19628_, _19627_, _23698_);
  not (_19629_, _19628_);
  nand (_19630_, _19629_, _19189_);
  nor (_19631_, _19189_, _08704_);
  nor (_19633_, _19631_, _19199_);
  nand (_19634_, _19633_, _19630_);
  not (_19635_, _08431_);
  nor (_19636_, _19194_, _19635_);
  nand (_19637_, _19636_, _19199_);
  nand (_19638_, _19637_, _19634_);
  nor (_19639_, _19638_, _19178_);
  nand (_19640_, _19088_, _08474_);
  nor (_19641_, _19640_, _23698_);
  nor (_19642_, _19641_, _19179_);
  nor (_19644_, _19642_, _19639_);
  nor (_19645_, _19644_, _19169_);
  nand (_19646_, _19160_, _08525_);
  nor (_19647_, _19646_, _23698_);
  nor (_19648_, _19647_, _19170_);
  nor (_08371_, _19648_, _19645_);
  nand (_19649_, _18823_, _08405_);
  nor (_19650_, _19649_, _23698_);
  not (_19651_, _19650_);
  nand (_19652_, _19651_, _19189_);
  nor (_19653_, _19189_, _08709_);
  nor (_19654_, _19653_, _19199_);
  nand (_19655_, _19654_, _19652_);
  not (_19656_, _08436_);
  nor (_19657_, _19194_, _19656_);
  nand (_19658_, _19657_, _19199_);
  nand (_19659_, _19658_, _19655_);
  nor (_19660_, _19659_, _19178_);
  nand (_19661_, _19088_, _08479_);
  nor (_19662_, _19661_, _23698_);
  nor (_19663_, _19662_, _19179_);
  nor (_19664_, _19663_, _19660_);
  nor (_19665_, _19664_, _19169_);
  nand (_19666_, _19160_, _08530_);
  nor (_19667_, _19666_, _23698_);
  nor (_19668_, _19667_, _19170_);
  nor (_08375_, _19668_, _19665_);
  nand (_19669_, _18823_, _08410_);
  nor (_19670_, _19669_, _23698_);
  not (_19671_, _19670_);
  nand (_19673_, _19671_, _19189_);
  nor (_19674_, _19189_, _08713_);
  nor (_19675_, _19674_, _19199_);
  nand (_19676_, _19675_, _19673_);
  not (_19677_, _08441_);
  nor (_19678_, _19194_, _19677_);
  nand (_19679_, _19678_, _19199_);
  nand (_19680_, _19679_, _19676_);
  nor (_19681_, _19680_, _19178_);
  nand (_19682_, _19088_, _08484_);
  nor (_19684_, _19682_, _23698_);
  nor (_19685_, _19684_, _19179_);
  nor (_19686_, _19685_, _19681_);
  nor (_19687_, _19686_, _19169_);
  nand (_19688_, _19160_, _08535_);
  nor (_19689_, _19688_, _23698_);
  nor (_19690_, _19689_, _19170_);
  nor (_08380_, _19690_, _19687_);
  nand (_19691_, _18823_, _08414_);
  nor (_19692_, _19691_, _23698_);
  not (_19693_, _19692_);
  nand (_19694_, _19693_, _19189_);
  nor (_19695_, _19189_, _08558_);
  nor (_19696_, _19695_, _19199_);
  nand (_19697_, _19696_, _19694_);
  not (_19698_, _08447_);
  nor (_19699_, _19194_, _19698_);
  nand (_19700_, _19699_, _19199_);
  nand (_19701_, _19700_, _19697_);
  nor (_19702_, _19701_, _19178_);
  nand (_19703_, _19088_, _08489_);
  nor (_19704_, _19703_, _23698_);
  nor (_19705_, _19704_, _19179_);
  nor (_19706_, _19705_, _19702_);
  nor (_19707_, _19706_, _19169_);
  nand (_19708_, _19160_, _08540_);
  nor (_19709_, _19708_, _23698_);
  nor (_19710_, _19709_, _19170_);
  nor (_08384_, _19710_, _19707_);
  nand (_19711_, _18823_, _08418_);
  nor (_19714_, _19711_, _23698_);
  not (_19715_, _19714_);
  nand (_19716_, _19715_, _19189_);
  nor (_19717_, _19189_, _08731_);
  nor (_19718_, _19717_, _19199_);
  nand (_19719_, _19718_, _19716_);
  not (_19720_, _08452_);
  nor (_19721_, _19194_, _19720_);
  nand (_19722_, _19721_, _19199_);
  nand (_19723_, _19722_, _19719_);
  nor (_19725_, _19723_, _19178_);
  nand (_19726_, _19088_, _08494_);
  nor (_19727_, _19726_, _23698_);
  nor (_19728_, _19727_, _19179_);
  nor (_19729_, _19728_, _19725_);
  nor (_19730_, _19729_, _19169_);
  nand (_19731_, _19160_, _08545_);
  nor (_19732_, _19731_, _23698_);
  nor (_19733_, _19732_, _19170_);
  nor (_08388_, _19733_, _19730_);
  nand (_19734_, _18823_, _08422_);
  nor (_19735_, _19734_, _23698_);
  not (_19736_, _19735_);
  nand (_19737_, _19736_, _19189_);
  nor (_19738_, _19189_, _08736_);
  nor (_19739_, _19738_, _19199_);
  nand (_19740_, _19739_, _19737_);
  not (_19741_, _08457_);
  nor (_19742_, _19194_, _19741_);
  nand (_19743_, _19742_, _19199_);
  nand (_19744_, _19743_, _19740_);
  nor (_19745_, _19744_, _19178_);
  nand (_19746_, _19088_, _08499_);
  nor (_19747_, _19746_, _23698_);
  nor (_19748_, _19747_, _19179_);
  nor (_19749_, _19748_, _19745_);
  nor (_19750_, _19749_, _19169_);
  nand (_19751_, _19160_, _08550_);
  nor (_19752_, _19751_, _23698_);
  nor (_19753_, _19752_, _19170_);
  nor (_08392_, _19753_, _19750_);
  nor (_19755_, _18794_, _08902_);
  nor (_19756_, _18743_, _08900_);
  nor (_19757_, _19756_, _19755_);
  nor (_19758_, _19757_, _18747_);
  nor (_19759_, _18794_, _08849_);
  nor (_19760_, _18743_, _08847_);
  nor (_19761_, _19760_, _19759_);
  nor (_19762_, _19761_, _18774_);
  nor (_19763_, _19762_, _19758_);
  nand (_19765_, _19763_, _18751_);
  not (_19766_, _08567_);
  nand (_19767_, _18743_, _19766_);
  not (_19768_, _08565_);
  nand (_19769_, _18794_, _19768_);
  nand (_19770_, _19769_, _19767_);
  nor (_19771_, _19770_, _18849_);
  not (_19772_, _08699_);
  nand (_19773_, _18743_, _19772_);
  not (_19774_, _08696_);
  nand (_19775_, _18794_, _19774_);
  nand (_19776_, _19775_, _19773_);
  nor (_19777_, _19776_, _18783_);
  nor (_19778_, _19777_, _19771_);
  nand (_19779_, _19778_, _19765_);
  nand (_19780_, _19779_, _18754_);
  nor (_19781_, _18794_, _09060_);
  nor (_19782_, _18743_, _09058_);
  nor (_19783_, _19782_, _19781_);
  nor (_19784_, _19783_, _18747_);
  nor (_19785_, _18794_, _08512_);
  nor (_19786_, _18743_, _08510_);
  nor (_19787_, _19786_, _19785_);
  nor (_19788_, _19787_, _18774_);
  nor (_19789_, _19788_, _19784_);
  nand (_19790_, _19789_, _18751_);
  nor (_19791_, _18794_, _08988_);
  nor (_19792_, _18743_, _08986_);
  nor (_19793_, _19792_, _19791_);
  nand (_19794_, _19793_, _18774_);
  nor (_19795_, _18794_, _08938_);
  nor (_19796_, _18743_, _08936_);
  nor (_19797_, _19796_, _19795_);
  nand (_19798_, _19797_, _18747_);
  nand (_19799_, _19798_, _19794_);
  nand (_19800_, _19799_, _18750_);
  nand (_19801_, _19800_, _19790_);
  nand (_19802_, _19801_, _18755_);
  nand (_19803_, _19802_, _19780_);
  nand (_19804_, _19803_, _18824_);
  nand (_08398_, _19804_, _19607_);
  nor (_19805_, _18794_, _08907_);
  nor (_19806_, _18743_, _08905_);
  nor (_19807_, _19806_, _19805_);
  nor (_19808_, _19807_, _18747_);
  nor (_19809_, _18794_, _08854_);
  nor (_19810_, _18743_, _08852_);
  nor (_19811_, _19810_, _19809_);
  nor (_19812_, _19811_, _18774_);
  nor (_19813_, _19812_, _19808_);
  nand (_19814_, _19813_, _18751_);
  nor (_19815_, _18794_, _08704_);
  nor (_19816_, _18743_, _08702_);
  nor (_19817_, _19816_, _19815_);
  not (_19818_, _19817_);
  nor (_19819_, _19818_, _18783_);
  nor (_19820_, _18794_, _08811_);
  nor (_19821_, _18743_, _08809_);
  nor (_19822_, _19821_, _19820_);
  not (_19823_, _19822_);
  nor (_19824_, _19823_, _18849_);
  nor (_19825_, _19824_, _19819_);
  nand (_19826_, _19825_, _19814_);
  nand (_19827_, _19826_, _18754_);
  nor (_19828_, _18794_, _08506_);
  nor (_19829_, _18743_, _08504_);
  nor (_19830_, _19829_, _19828_);
  nor (_19831_, _19830_, _18747_);
  nor (_19832_, _18794_, _09034_);
  nor (_19833_, _18743_, _09032_);
  nor (_19834_, _19833_, _19832_);
  nor (_19835_, _19834_, _18774_);
  nor (_19836_, _19835_, _19831_);
  nand (_19837_, _19836_, _18751_);
  nor (_19838_, _18794_, _08995_);
  nor (_19839_, _18743_, _08993_);
  nor (_19840_, _19839_, _19838_);
  nand (_19841_, _19840_, _18774_);
  nor (_19842_, _18794_, _08944_);
  nor (_19843_, _18743_, _08942_);
  nor (_19845_, _19843_, _19842_);
  nand (_19846_, _19845_, _18747_);
  nand (_19847_, _19846_, _19841_);
  nand (_19848_, _19847_, _18750_);
  nand (_19849_, _19848_, _19837_);
  nand (_19850_, _19849_, _18755_);
  nand (_19851_, _19850_, _19827_);
  nand (_19852_, _19851_, _18824_);
  nand (_08403_, _19852_, _19627_);
  nor (_19853_, _18794_, _08913_);
  nor (_19855_, _18743_, _08911_);
  nor (_19856_, _19855_, _19853_);
  nor (_19857_, _19856_, _18747_);
  nor (_19858_, _18794_, _08861_);
  nor (_19859_, _18743_, _08859_);
  nor (_19860_, _19859_, _19858_);
  nor (_19861_, _19860_, _18774_);
  nor (_19862_, _19861_, _19857_);
  nand (_19863_, _19862_, _18751_);
  not (_19864_, _08816_);
  nand (_19865_, _18743_, _19864_);
  not (_19866_, _08814_);
  nand (_19867_, _18794_, _19866_);
  nand (_19868_, _19867_, _19865_);
  nor (_19869_, _19868_, _18849_);
  not (_19870_, _08709_);
  nand (_19871_, _18743_, _19870_);
  not (_19872_, _08707_);
  nand (_19873_, _18794_, _19872_);
  nand (_19874_, _19873_, _19871_);
  nor (_19875_, _19874_, _18783_);
  nor (_19876_, _19875_, _19869_);
  nand (_19877_, _19876_, _19863_);
  nand (_19878_, _19877_, _18754_);
  nor (_19879_, _18794_, _09644_);
  nor (_19880_, _18743_, _09696_);
  nor (_19881_, _19880_, _19879_);
  nor (_19882_, _19881_, _18747_);
  nor (_19883_, _18794_, _09039_);
  nor (_19884_, _18743_, _09037_);
  nor (_19886_, _19884_, _19883_);
  nor (_19887_, _19886_, _18774_);
  nor (_19888_, _19887_, _19882_);
  nand (_19889_, _19888_, _18751_);
  nor (_19890_, _18794_, _09000_);
  nor (_19891_, _18743_, _08998_);
  nor (_19892_, _19891_, _19890_);
  nand (_19893_, _19892_, _18774_);
  nor (_19894_, _18794_, _08952_);
  nor (_19895_, _18743_, _08950_);
  nor (_19897_, _19895_, _19894_);
  nand (_19898_, _19897_, _18747_);
  nand (_19899_, _19898_, _19893_);
  nand (_19900_, _19899_, _18750_);
  nand (_19901_, _19900_, _19889_);
  nand (_19902_, _19901_, _18755_);
  nand (_19903_, _19902_, _19878_);
  nand (_19904_, _19903_, _18824_);
  nand (_08408_, _19904_, _19649_);
  nor (_19905_, _18794_, _08918_);
  nor (_19906_, _18743_, _08916_);
  nor (_19907_, _19906_, _19905_);
  nor (_19908_, _19907_, _18747_);
  nor (_19909_, _18794_, _08866_);
  nor (_19910_, _18743_, _08864_);
  nor (_19911_, _19910_, _19909_);
  nor (_19912_, _19911_, _18774_);
  nor (_19913_, _19912_, _19908_);
  nand (_19914_, _19913_, _18751_);
  nor (_19915_, _18794_, _08713_);
  nor (_19916_, _18743_, _08711_);
  nor (_19917_, _19916_, _19915_);
  not (_19918_, _19917_);
  nor (_19919_, _19918_, _18783_);
  nor (_19920_, _18794_, _08820_);
  nor (_19921_, _18743_, _08818_);
  nor (_19922_, _19921_, _19920_);
  not (_19923_, _19922_);
  nor (_19924_, _19923_, _18849_);
  nor (_19925_, _19924_, _19919_);
  nand (_19927_, _19925_, _19914_);
  nand (_19928_, _19927_, _18754_);
  nor (_19929_, _18794_, _09646_);
  nor (_19930_, _18743_, _09698_);
  nor (_19931_, _19930_, _19929_);
  nor (_19932_, _19931_, _18747_);
  nor (_19933_, _18794_, _09045_);
  nor (_19934_, _18743_, _09043_);
  nor (_19935_, _19934_, _19933_);
  nor (_19936_, _19935_, _18774_);
  nor (_19938_, _19936_, _19932_);
  nand (_19939_, _19938_, _18751_);
  nor (_19940_, _18794_, _09005_);
  nor (_19941_, _18743_, _09003_);
  nor (_19942_, _19941_, _19940_);
  nand (_19943_, _19942_, _18774_);
  nor (_19944_, _18794_, _08517_);
  nor (_19945_, _18743_, _08515_);
  nor (_19946_, _19945_, _19944_);
  nand (_19947_, _19946_, _18747_);
  nand (_19948_, _19947_, _19943_);
  nand (_19949_, _19948_, _18750_);
  nand (_19950_, _19949_, _19939_);
  nand (_19951_, _19950_, _18755_);
  nand (_19952_, _19951_, _19928_);
  nand (_19953_, _19952_, _18824_);
  nand (_08412_, _19953_, _19669_);
  nor (_19954_, _18794_, _08923_);
  nor (_19955_, _18743_, _08921_);
  nor (_19956_, _19955_, _19954_);
  nor (_19957_, _19956_, _18747_);
  nor (_19958_, _18794_, _08878_);
  nor (_19959_, _18743_, _08876_);
  nor (_19960_, _19959_, _19958_);
  nor (_19961_, _19960_, _18774_);
  nor (_19962_, _19961_, _19957_);
  nand (_19963_, _19962_, _18751_);
  nor (_19964_, _18794_, _08558_);
  nor (_19965_, _18743_, _08556_);
  nor (_19966_, _19965_, _19964_);
  not (_19968_, _19966_);
  nor (_19969_, _19968_, _18783_);
  nor (_19970_, _18794_, _08827_);
  nor (_19971_, _18743_, _08825_);
  nor (_19972_, _19971_, _19970_);
  not (_19973_, _19972_);
  nor (_19974_, _19973_, _18849_);
  nor (_19975_, _19974_, _19969_);
  nand (_19976_, _19975_, _19963_);
  nand (_19977_, _19976_, _18754_);
  nor (_19979_, _18794_, _09648_);
  nor (_19980_, _18743_, _09700_);
  nor (_19981_, _19980_, _19979_);
  nor (_19982_, _19981_, _18747_);
  nor (_19983_, _18794_, _09050_);
  nor (_19984_, _18743_, _09048_);
  nor (_19985_, _19984_, _19983_);
  nor (_19986_, _19985_, _18774_);
  nor (_19987_, _19986_, _19982_);
  nand (_19988_, _19987_, _18751_);
  nor (_19989_, _18794_, _09012_);
  nor (_19990_, _18743_, _09010_);
  nor (_19991_, _19990_, _19989_);
  nand (_19992_, _19991_, _18774_);
  nor (_19993_, _18794_, _08971_);
  nor (_19994_, _18743_, _08969_);
  nor (_19995_, _19994_, _19993_);
  nand (_19996_, _19995_, _18747_);
  nand (_19997_, _19996_, _19992_);
  nand (_19998_, _19997_, _18750_);
  nand (_19999_, _19998_, _19988_);
  nand (_20000_, _19999_, _18755_);
  nand (_20001_, _20000_, _19977_);
  nand (_20002_, _20001_, _18824_);
  nand (_08416_, _20002_, _19691_);
  nor (_20003_, _18794_, _09056_);
  nor (_20004_, _18743_, _09054_);
  nor (_20005_, _20004_, _20003_);
  nand (_20006_, _20005_, _18747_);
  nor (_20007_, _18794_, _09649_);
  nor (_20009_, _18743_, _09702_);
  nor (_20010_, _20009_, _20007_);
  nand (_20011_, _20010_, _18774_);
  nand (_20012_, _20011_, _20006_);
  nand (_20013_, _20012_, _18751_);
  nor (_20014_, _18794_, _09018_);
  nor (_20015_, _18743_, _09016_);
  nor (_20016_, _20015_, _20014_);
  nand (_20017_, _20016_, _18836_);
  nand (_20018_, _20017_, _20013_);
  nand (_20020_, _20018_, _18755_);
  not (_20021_, _07607_);
  nand (_20022_, _18743_, _20021_);
  not (_20023_, _07605_);
  nand (_20024_, _18794_, _20023_);
  nand (_20025_, _20024_, _20022_);
  nor (_20026_, _20025_, _19469_);
  nor (_20027_, _18794_, _08928_);
  nor (_20028_, _18743_, _08926_);
  nor (_20029_, _20028_, _20027_);
  not (_20030_, _20029_);
  nand (_20031_, _20030_, _18774_);
  nor (_20032_, _18794_, _08573_);
  nor (_20033_, _18743_, _08570_);
  nor (_20034_, _20033_, _20032_);
  not (_20035_, _20034_);
  nand (_20036_, _20035_, _18747_);
  nand (_20037_, _20036_, _20031_);
  nor (_20038_, _20037_, _18750_);
  nor (_20039_, _18794_, _08832_);
  nor (_20040_, _18743_, _08830_);
  nor (_20041_, _20040_, _20039_);
  nand (_20042_, _20041_, _18836_);
  nor (_20043_, _18794_, _08731_);
  nor (_20044_, _18743_, _08729_);
  nor (_20045_, _20044_, _20043_);
  nand (_20046_, _20045_, _18782_);
  nand (_20047_, _20046_, _20042_);
  nor (_20048_, _20047_, _20038_);
  nor (_20049_, _20048_, _18755_);
  nor (_20051_, _20049_, _20026_);
  nand (_20052_, _20051_, _20020_);
  nand (_20053_, _20052_, _18824_);
  nand (_08420_, _20053_, _19711_);
  nor (_20054_, _18794_, _08578_);
  nor (_20055_, _18743_, _08576_);
  nor (_20056_, _20055_, _20054_);
  nand (_20057_, _20056_, _18747_);
  nor (_20058_, _18794_, _09651_);
  nor (_20059_, _18743_, _09704_);
  nor (_20061_, _20059_, _20058_);
  nand (_20062_, _20061_, _18774_);
  nand (_20063_, _20062_, _20057_);
  nand (_20064_, _20063_, _18751_);
  nor (_20065_, _18794_, _09023_);
  nor (_20066_, _18743_, _09021_);
  nor (_20067_, _20066_, _20065_);
  nand (_20068_, _20067_, _18836_);
  nand (_20069_, _20068_, _20064_);
  nand (_20070_, _20069_, _18755_);
  not (_20071_, _08982_);
  nand (_20072_, _18743_, _20071_);
  not (_20073_, _08980_);
  nand (_20074_, _18794_, _20073_);
  nand (_20075_, _20074_, _20072_);
  nor (_20076_, _20075_, _19469_);
  nor (_20077_, _18794_, _08934_);
  nor (_20078_, _18743_, _08932_);
  nor (_20079_, _20078_, _20077_);
  not (_20080_, _20079_);
  nand (_20081_, _20080_, _18774_);
  nor (_20082_, _18794_, _08898_);
  nor (_20083_, _18743_, _08895_);
  nor (_20084_, _20083_, _20082_);
  not (_20085_, _20084_);
  nand (_20086_, _20085_, _18747_);
  nand (_20087_, _20086_, _20081_);
  nor (_20088_, _20087_, _18750_);
  nor (_20089_, _18794_, _08837_);
  nor (_20090_, _18743_, _08835_);
  nor (_20092_, _20090_, _20089_);
  nand (_20093_, _20092_, _18836_);
  nor (_20094_, _18794_, _08736_);
  nor (_20095_, _18743_, _08734_);
  nor (_20096_, _20095_, _20094_);
  nand (_20097_, _20096_, _18782_);
  nand (_20098_, _20097_, _20093_);
  nor (_20099_, _20098_, _20088_);
  nor (_20100_, _20099_, _18755_);
  nor (_20101_, _20100_, _20076_);
  nand (_20103_, _20101_, _20070_);
  nand (_20104_, _20103_, _18824_);
  nand (_08424_, _20104_, _19734_);
  nand (_20105_, _19007_, _08426_);
  nor (_20106_, _18794_, _08847_);
  nor (_20107_, _18743_, _08849_);
  nor (_20108_, _20107_, _20106_);
  nand (_20109_, _20108_, _18962_);
  nor (_20110_, _18794_, _08900_);
  nor (_20111_, _18743_, _08902_);
  nor (_20112_, _20111_, _20110_);
  nand (_20113_, _20112_, _18957_);
  nand (_20114_, _20113_, _20109_);
  nand (_20115_, _20114_, _18898_);
  nor (_20116_, _18794_, _08565_);
  nor (_20117_, _18743_, _08567_);
  nor (_20118_, _20117_, _20116_);
  nand (_20119_, _20118_, _18957_);
  nor (_20120_, _18794_, _08696_);
  nor (_20121_, _18743_, _08699_);
  nor (_20123_, _20121_, _20120_);
  nand (_20124_, _20123_, _18962_);
  nand (_20125_, _20124_, _20119_);
  nand (_20126_, _20125_, _18886_);
  nand (_20127_, _20126_, _20115_);
  nand (_20128_, _20127_, _18891_);
  nor (_20129_, _18794_, _08510_);
  nor (_20130_, _18743_, _08512_);
  nor (_20131_, _20130_, _20129_);
  nand (_20132_, _20131_, _18962_);
  nor (_20134_, _18794_, _09058_);
  nor (_20135_, _18743_, _09060_);
  nor (_20136_, _20135_, _20134_);
  nand (_20137_, _20136_, _18957_);
  nand (_20138_, _20137_, _20132_);
  nand (_20139_, _20138_, _18898_);
  nor (_20140_, _18794_, _08986_);
  nor (_20141_, _18743_, _08988_);
  nor (_20142_, _20141_, _20140_);
  nand (_20143_, _20142_, _18957_);
  nor (_20145_, _18794_, _08936_);
  nor (_20146_, _18743_, _08938_);
  nor (_20147_, _20146_, _20145_);
  nand (_20148_, _20147_, _18962_);
  nand (_20149_, _20148_, _20143_);
  nand (_20150_, _20149_, _18886_);
  nand (_20151_, _20150_, _20139_);
  nand (_20152_, _20151_, _18894_);
  nand (_20153_, _20152_, _20128_);
  nand (_20154_, _20153_, _18956_);
  nand (_08429_, _20154_, _20105_);
  nand (_20155_, _19007_, _08431_);
  nor (_20156_, _18794_, _08852_);
  nor (_20157_, _18743_, _08854_);
  nor (_20158_, _20157_, _20156_);
  nand (_20159_, _20158_, _18962_);
  nor (_20160_, _18794_, _08905_);
  nor (_20161_, _18743_, _08907_);
  nor (_20162_, _20161_, _20160_);
  nand (_20163_, _20162_, _18957_);
  nand (_20164_, _20163_, _20159_);
  nand (_20165_, _20164_, _18898_);
  nor (_20166_, _18794_, _08809_);
  nor (_20167_, _18743_, _08811_);
  nor (_20168_, _20167_, _20166_);
  nand (_20169_, _20168_, _18957_);
  nor (_20170_, _18794_, _08702_);
  nor (_20171_, _18743_, _08704_);
  nor (_20172_, _20171_, _20170_);
  nand (_20173_, _20172_, _18962_);
  nand (_20175_, _20173_, _20169_);
  nand (_20176_, _20175_, _18886_);
  nand (_20177_, _20176_, _20165_);
  nand (_20178_, _20177_, _18891_);
  nor (_20179_, _18794_, _09032_);
  nor (_20180_, _18743_, _09034_);
  nor (_20181_, _20180_, _20179_);
  nand (_20182_, _20181_, _18962_);
  nor (_20183_, _18794_, _08504_);
  nor (_20184_, _18743_, _08506_);
  nor (_20186_, _20184_, _20183_);
  nand (_20187_, _20186_, _18957_);
  nand (_20188_, _20187_, _20182_);
  nand (_20189_, _20188_, _18898_);
  nor (_20190_, _18794_, _08993_);
  nor (_20191_, _18743_, _08995_);
  nor (_20192_, _20191_, _20190_);
  nand (_20193_, _20192_, _18957_);
  nor (_20194_, _18794_, _08942_);
  nor (_20195_, _18743_, _08944_);
  nor (_20196_, _20195_, _20194_);
  nand (_20197_, _20196_, _18962_);
  nand (_20198_, _20197_, _20193_);
  nand (_20199_, _20198_, _18886_);
  nand (_20200_, _20199_, _20189_);
  nand (_20201_, _20200_, _18894_);
  nand (_20202_, _20201_, _20178_);
  nand (_20203_, _20202_, _18956_);
  nand (_08434_, _20203_, _20155_);
  nand (_20204_, _19007_, _08436_);
  nor (_20205_, _18794_, _08859_);
  nor (_20206_, _18743_, _08861_);
  nor (_20207_, _20206_, _20205_);
  nand (_20208_, _20207_, _18962_);
  nor (_20209_, _18794_, _08911_);
  nor (_20210_, _18743_, _08913_);
  nor (_20211_, _20210_, _20209_);
  nand (_20212_, _20211_, _18957_);
  nand (_20213_, _20212_, _20208_);
  nand (_20214_, _20213_, _18898_);
  nor (_20216_, _18794_, _08814_);
  nor (_20217_, _18743_, _08816_);
  nor (_20218_, _20217_, _20216_);
  nand (_20219_, _20218_, _18957_);
  nor (_20220_, _18794_, _08707_);
  nor (_20221_, _18743_, _08709_);
  nor (_20222_, _20221_, _20220_);
  nand (_20223_, _20222_, _18962_);
  nand (_20224_, _20223_, _20219_);
  nand (_20225_, _20224_, _18886_);
  nand (_20227_, _20225_, _20214_);
  nand (_20228_, _20227_, _18891_);
  nor (_20229_, _18794_, _09037_);
  nor (_20230_, _18743_, _09039_);
  nor (_20231_, _20230_, _20229_);
  nand (_20232_, _20231_, _18962_);
  nor (_20233_, _18794_, _09696_);
  nor (_20234_, _18743_, _09644_);
  nor (_20235_, _20234_, _20233_);
  nand (_20236_, _20235_, _18957_);
  nand (_20237_, _20236_, _20232_);
  nand (_20238_, _20237_, _18898_);
  nor (_20239_, _18794_, _08998_);
  nor (_20240_, _18743_, _09000_);
  nor (_20241_, _20240_, _20239_);
  nand (_20242_, _20241_, _18957_);
  nor (_20243_, _18794_, _08950_);
  nor (_20244_, _18743_, _08952_);
  nor (_20245_, _20244_, _20243_);
  nand (_20246_, _20245_, _18962_);
  nand (_20247_, _20246_, _20242_);
  nand (_20248_, _20247_, _18886_);
  nand (_20249_, _20248_, _20238_);
  nand (_20250_, _20249_, _18894_);
  nand (_20251_, _20250_, _20228_);
  nand (_20252_, _20251_, _18956_);
  nand (_08439_, _20252_, _20204_);
  nand (_20253_, _19007_, _08441_);
  nor (_20254_, _18794_, _08864_);
  nor (_20255_, _18743_, _08866_);
  nor (_20257_, _20255_, _20254_);
  nand (_20258_, _20257_, _18962_);
  nor (_20259_, _18794_, _08916_);
  nor (_20260_, _18743_, _08918_);
  nor (_20261_, _20260_, _20259_);
  nand (_20262_, _20261_, _18957_);
  nand (_20263_, _20262_, _20258_);
  nand (_20264_, _20263_, _18898_);
  nor (_20265_, _18794_, _08818_);
  nor (_20266_, _18743_, _08820_);
  nor (_20268_, _20266_, _20265_);
  nand (_20269_, _20268_, _18957_);
  nor (_20270_, _18794_, _08711_);
  nor (_20271_, _18743_, _08713_);
  nor (_20272_, _20271_, _20270_);
  nand (_20273_, _20272_, _18962_);
  nand (_20274_, _20273_, _20269_);
  nand (_20275_, _20274_, _18886_);
  nand (_20276_, _20275_, _20264_);
  nand (_20277_, _20276_, _18891_);
  nor (_20278_, _18794_, _09043_);
  nor (_20279_, _18743_, _09045_);
  nor (_20280_, _20279_, _20278_);
  nand (_20281_, _20280_, _18962_);
  nor (_20282_, _18794_, _09698_);
  nor (_20283_, _18743_, _09646_);
  nor (_20284_, _20283_, _20282_);
  nand (_20285_, _20284_, _18957_);
  nand (_20286_, _20285_, _20281_);
  nand (_20287_, _20286_, _18898_);
  nor (_20288_, _18794_, _09003_);
  nor (_20289_, _18743_, _09005_);
  nor (_20290_, _20289_, _20288_);
  nand (_20291_, _20290_, _18957_);
  nor (_20292_, _18794_, _08515_);
  nor (_20293_, _18743_, _08517_);
  nor (_20294_, _20293_, _20292_);
  nand (_20295_, _20294_, _18962_);
  nand (_20296_, _20295_, _20291_);
  nand (_20297_, _20296_, _18886_);
  nand (_20299_, _20297_, _20287_);
  nand (_20300_, _20299_, _18894_);
  nand (_20301_, _20300_, _20277_);
  nand (_20302_, _20301_, _18956_);
  nand (_08445_, _20302_, _20253_);
  nand (_20303_, _19007_, _08447_);
  nor (_20304_, _18794_, _08876_);
  nor (_20305_, _18743_, _08878_);
  nor (_20306_, _20305_, _20304_);
  nand (_20307_, _20306_, _18962_);
  nor (_20309_, _18794_, _08921_);
  nor (_20310_, _18743_, _08923_);
  nor (_20311_, _20310_, _20309_);
  nand (_20312_, _20311_, _18957_);
  nand (_20313_, _20312_, _20307_);
  nand (_20314_, _20313_, _18898_);
  nor (_20315_, _18794_, _08825_);
  nor (_20316_, _18743_, _08827_);
  nor (_20317_, _20316_, _20315_);
  nand (_20318_, _20317_, _18957_);
  nor (_20319_, _18794_, _08556_);
  nor (_20320_, _18743_, _08558_);
  nor (_20321_, _20320_, _20319_);
  nand (_20322_, _20321_, _18962_);
  nand (_20323_, _20322_, _20318_);
  nand (_20324_, _20323_, _18886_);
  nand (_20325_, _20324_, _20314_);
  nand (_20326_, _20325_, _18891_);
  nor (_20327_, _18794_, _09700_);
  nor (_20328_, _18743_, _09648_);
  nor (_20329_, _20328_, _20327_);
  nand (_20330_, _20329_, _18957_);
  nor (_20331_, _18794_, _09048_);
  nor (_20332_, _18743_, _09050_);
  nor (_20333_, _20332_, _20331_);
  nand (_20334_, _20333_, _18962_);
  nand (_20335_, _20334_, _20330_);
  nand (_20336_, _20335_, _18898_);
  nor (_20337_, _18794_, _08969_);
  nor (_20338_, _18743_, _08971_);
  nor (_20340_, _20338_, _20337_);
  nand (_20341_, _20340_, _18962_);
  nor (_20342_, _18794_, _09010_);
  nor (_20343_, _18743_, _09012_);
  nor (_20344_, _20343_, _20342_);
  nand (_20345_, _20344_, _18957_);
  nand (_20346_, _20345_, _20341_);
  nand (_20347_, _20346_, _18886_);
  nand (_20348_, _20347_, _20336_);
  nand (_20349_, _20348_, _18894_);
  nand (_20351_, _20349_, _20326_);
  nand (_20352_, _20351_, _18956_);
  nand (_08450_, _20352_, _20303_);
  nand (_20353_, _19007_, _08452_);
  nor (_20354_, _18794_, _08570_);
  nor (_20355_, _18743_, _08573_);
  nor (_20356_, _20355_, _20354_);
  nand (_20357_, _20356_, _18962_);
  nor (_20358_, _18794_, _08926_);
  nor (_20359_, _18743_, _08928_);
  nor (_20360_, _20359_, _20358_);
  nand (_20361_, _20360_, _18957_);
  nand (_20362_, _20361_, _20357_);
  nand (_20363_, _20362_, _18898_);
  nor (_20364_, _18794_, _08830_);
  nor (_20365_, _18743_, _08832_);
  nor (_20366_, _20365_, _20364_);
  nand (_20367_, _20366_, _18957_);
  nor (_20368_, _18794_, _08729_);
  nor (_20369_, _18743_, _08731_);
  nor (_20370_, _20369_, _20368_);
  nand (_20371_, _20370_, _18962_);
  nand (_20372_, _20371_, _20367_);
  nand (_20373_, _20372_, _18886_);
  nand (_20374_, _20373_, _20363_);
  nand (_20375_, _20374_, _18891_);
  nor (_20376_, _18794_, _09054_);
  nor (_20377_, _18743_, _09056_);
  nor (_20378_, _20377_, _20376_);
  nand (_20379_, _20378_, _18962_);
  nor (_20381_, _18794_, _09702_);
  nor (_20382_, _18743_, _09649_);
  nor (_20383_, _20382_, _20381_);
  nand (_20384_, _20383_, _18957_);
  nand (_20385_, _20384_, _20379_);
  nand (_20386_, _20385_, _18898_);
  nor (_20387_, _18794_, _09016_);
  nor (_20388_, _18743_, _09018_);
  nor (_20389_, _20388_, _20387_);
  nand (_20390_, _20389_, _18957_);
  nor (_20392_, _18794_, _07605_);
  nor (_20393_, _18743_, _07607_);
  nor (_20394_, _20393_, _20392_);
  nand (_20395_, _20394_, _18962_);
  nand (_20396_, _20395_, _20390_);
  nand (_20397_, _20396_, _18886_);
  nand (_20398_, _20397_, _20386_);
  nand (_20399_, _20398_, _18894_);
  nand (_20400_, _20399_, _20375_);
  nand (_20401_, _20400_, _18956_);
  nand (_08455_, _20401_, _20353_);
  nand (_20402_, _19007_, _08457_);
  nor (_20403_, _18794_, _08895_);
  nor (_20404_, _18743_, _08898_);
  nor (_20405_, _20404_, _20403_);
  nand (_20406_, _20405_, _18962_);
  nor (_20407_, _18794_, _08932_);
  nor (_20408_, _18743_, _08934_);
  nor (_20409_, _20408_, _20407_);
  nand (_20410_, _20409_, _18957_);
  nand (_20411_, _20410_, _20406_);
  nand (_20412_, _20411_, _18898_);
  nor (_20413_, _18794_, _08835_);
  nor (_20414_, _18743_, _08837_);
  nor (_20415_, _20414_, _20413_);
  nand (_20416_, _20415_, _18957_);
  nor (_20417_, _18794_, _08734_);
  nor (_20418_, _18743_, _08736_);
  nor (_20419_, _20418_, _20417_);
  nand (_20420_, _20419_, _18962_);
  nand (_20422_, _20420_, _20416_);
  nand (_20423_, _20422_, _18886_);
  nand (_20424_, _20423_, _20412_);
  nand (_20425_, _20424_, _18891_);
  nor (_20426_, _18794_, _08576_);
  nor (_20427_, _18743_, _08578_);
  nor (_20428_, _20427_, _20426_);
  nand (_20429_, _20428_, _18962_);
  nor (_20430_, _18794_, _09704_);
  nor (_20431_, _18743_, _09651_);
  nor (_20433_, _20431_, _20430_);
  nand (_20434_, _20433_, _18957_);
  nand (_20435_, _20434_, _20429_);
  nand (_20436_, _20435_, _18898_);
  nor (_20437_, _18794_, _09021_);
  nor (_20438_, _18743_, _09023_);
  nor (_20439_, _20438_, _20437_);
  nand (_20440_, _20439_, _18957_);
  nor (_20441_, _18794_, _08980_);
  nor (_20442_, _18743_, _08982_);
  nor (_20443_, _20442_, _20441_);
  nand (_20444_, _20443_, _18962_);
  nand (_20445_, _20444_, _20440_);
  nand (_20446_, _20445_, _18886_);
  nand (_20447_, _20446_, _20436_);
  nand (_20448_, _20447_, _18894_);
  nand (_20449_, _20448_, _20425_);
  nand (_20450_, _20449_, _18956_);
  nand (_08460_, _20450_, _20402_);
  nand (_20451_, _19783_, _18747_);
  nand (_20452_, _19787_, _18774_);
  nand (_20453_, _20452_, _20451_);
  nand (_20454_, _20453_, _19013_);
  nand (_20455_, _19793_, _18747_);
  nand (_20456_, _19797_, _18774_);
  nand (_20457_, _20456_, _20455_);
  nand (_20458_, _20457_, _19017_);
  nand (_20459_, _20458_, _20454_);
  nand (_20460_, _20459_, _19010_);
  nor (_20461_, _19761_, _18747_);
  nor (_20463_, _19757_, _18774_);
  nor (_20464_, _20463_, _20461_);
  nand (_20465_, _20464_, _19013_);
  nor (_20466_, _19770_, _18777_);
  nor (_20467_, _19776_, _18849_);
  nor (_20468_, _20467_, _20466_);
  nand (_20469_, _20468_, _20465_);
  nand (_20470_, _20469_, _19011_);
  nand (_20471_, _20470_, _20460_);
  nand (_20472_, _20471_, _19064_);
  nand (_08472_, _20472_, _19619_);
  nor (_20474_, _19834_, _18747_);
  nor (_20475_, _19830_, _18774_);
  nor (_20476_, _20475_, _20474_);
  nand (_20477_, _20476_, _19013_);
  nand (_20478_, _19840_, _18747_);
  nand (_20479_, _19845_, _18774_);
  nand (_20480_, _20479_, _20478_);
  nand (_20481_, _20480_, _19017_);
  nand (_20482_, _20481_, _20477_);
  nand (_20483_, _20482_, _19010_);
  nor (_20484_, _19811_, _18747_);
  nor (_20485_, _19807_, _18774_);
  nor (_20486_, _20485_, _20484_);
  nand (_20487_, _20486_, _19013_);
  nor (_20488_, _19818_, _18849_);
  nor (_20489_, _19823_, _18777_);
  nor (_20490_, _20489_, _20488_);
  nand (_20491_, _20490_, _20487_);
  nand (_20492_, _20491_, _19011_);
  nand (_20493_, _20492_, _20483_);
  nand (_20494_, _20493_, _19064_);
  nand (_08477_, _20494_, _19640_);
  nor (_20495_, _19886_, _18747_);
  nor (_20496_, _19881_, _18774_);
  nor (_20497_, _20496_, _20495_);
  nand (_20498_, _20497_, _19013_);
  nand (_20499_, _19897_, _18836_);
  nand (_20500_, _19892_, _18776_);
  nand (_20501_, _20500_, _20499_);
  nor (_20502_, _20501_, _19011_);
  nand (_20503_, _20502_, _20498_);
  nor (_20504_, _19860_, _18747_);
  nor (_20505_, _19856_, _18774_);
  nor (_20506_, _20505_, _20504_);
  nand (_20507_, _20506_, _19013_);
  nor (_20508_, _19874_, _18849_);
  nor (_20509_, _19868_, _18777_);
  nor (_20510_, _20509_, _20508_);
  nand (_20511_, _20510_, _20507_);
  nor (_20513_, _20511_, _19010_);
  nor (_20514_, _20513_, _19088_);
  nand (_20515_, _20514_, _20503_);
  nand (_08482_, _20515_, _19661_);
  nand (_20516_, _19931_, _18747_);
  nand (_20517_, _19935_, _18774_);
  nand (_20518_, _20517_, _20516_);
  nand (_20519_, _20518_, _19013_);
  nand (_20520_, _19942_, _18747_);
  nand (_20521_, _19946_, _18774_);
  nand (_20523_, _20521_, _20520_);
  nand (_20524_, _20523_, _19017_);
  nand (_20525_, _20524_, _20519_);
  nand (_20526_, _20525_, _19010_);
  nand (_20527_, _19907_, _18747_);
  nand (_20528_, _19911_, _18774_);
  nand (_20529_, _20528_, _20527_);
  nand (_20530_, _20529_, _19013_);
  nor (_20531_, _19918_, _18849_);
  nor (_20532_, _19923_, _18777_);
  nor (_20534_, _20532_, _20531_);
  nand (_20535_, _20534_, _20530_);
  nand (_20536_, _20535_, _19011_);
  nand (_20537_, _20536_, _20526_);
  nand (_20538_, _20537_, _19064_);
  nand (_08487_, _20538_, _19682_);
  nand (_20539_, _19981_, _18747_);
  nand (_20540_, _19985_, _18774_);
  nand (_20541_, _20540_, _20539_);
  nand (_20542_, _20541_, _19013_);
  nand (_20543_, _19991_, _18747_);
  nand (_20544_, _19995_, _18774_);
  nand (_20545_, _20544_, _20543_);
  nand (_20546_, _20545_, _19017_);
  nand (_20547_, _20546_, _20542_);
  nand (_20548_, _20547_, _19010_);
  nand (_20549_, _19956_, _18747_);
  nand (_20550_, _19960_, _18774_);
  nand (_20551_, _20550_, _20549_);
  nand (_20552_, _20551_, _19013_);
  nor (_20554_, _19968_, _18849_);
  nor (_20555_, _19973_, _18777_);
  nor (_20556_, _20555_, _20554_);
  nand (_20557_, _20556_, _20552_);
  nand (_20558_, _20557_, _19011_);
  nand (_20559_, _20558_, _20548_);
  nand (_20560_, _20559_, _19064_);
  nand (_08492_, _20560_, _19703_);
  nand (_20561_, _20010_, _18747_);
  nand (_20562_, _20005_, _18774_);
  nand (_20564_, _20562_, _20561_);
  nand (_20565_, _20564_, _19013_);
  nor (_20566_, _20025_, _18849_);
  not (_20567_, _20016_);
  nor (_20568_, _20567_, _18777_);
  nor (_20569_, _20568_, _20566_);
  nand (_20570_, _20569_, _20565_);
  nand (_20571_, _20570_, _19010_);
  nand (_20572_, _20029_, _18747_);
  nand (_20573_, _20034_, _18774_);
  nand (_20574_, _20573_, _20572_);
  nand (_20575_, _20574_, _19013_);
  nand (_20576_, _20041_, _18747_);
  nand (_20577_, _20045_, _18774_);
  nand (_20578_, _20577_, _20576_);
  nand (_20579_, _20578_, _19017_);
  nand (_20580_, _20579_, _20575_);
  nand (_20581_, _20580_, _19011_);
  nand (_20582_, _20581_, _20571_);
  nand (_20583_, _20582_, _19064_);
  nand (_08497_, _20583_, _19726_);
  nand (_20584_, _20061_, _18747_);
  nand (_20585_, _20056_, _18774_);
  nand (_20586_, _20585_, _20584_);
  nand (_20587_, _20586_, _19013_);
  not (_20588_, _20067_);
  nor (_20589_, _20588_, _18777_);
  nor (_20590_, _20075_, _18849_);
  nor (_20591_, _20590_, _20589_);
  nand (_20592_, _20591_, _20587_);
  nand (_20594_, _20592_, _19010_);
  nor (_20595_, _20084_, _18747_);
  nor (_20596_, _20079_, _18774_);
  nor (_20597_, _20596_, _20595_);
  nand (_20598_, _20597_, _19013_);
  nand (_20599_, _20092_, _18747_);
  nand (_20600_, _20096_, _18774_);
  nand (_20601_, _20600_, _20599_);
  nand (_20602_, _20601_, _19017_);
  nand (_20603_, _20602_, _20598_);
  nand (_20605_, _20603_, _19011_);
  nand (_20606_, _20605_, _20594_);
  nand (_20607_, _20606_, _19064_);
  nand (_08502_, _20607_, _19746_);
  nand (_20608_, _20118_, _18962_);
  nand (_20609_, _20123_, _18957_);
  nand (_20610_, _20609_, _20608_);
  nand (_20611_, _20610_, _19139_);
  not (_20612_, _20112_);
  nor (_20613_, _20612_, _18957_);
  not (_20614_, _20108_);
  nor (_20615_, _20614_, _18962_);
  nor (_20616_, _20615_, _20613_);
  nor (_20617_, _20616_, _19104_);
  nand (_20618_, _20136_, _18962_);
  nand (_20619_, _20131_, _18957_);
  nand (_20620_, _20619_, _20618_);
  nand (_20621_, _20620_, _19098_);
  nand (_20622_, _20142_, _18962_);
  nand (_20623_, _20147_, _18957_);
  nand (_20624_, _20623_, _20622_);
  nand (_20625_, _20624_, _19154_);
  nand (_20626_, _20625_, _20621_);
  nor (_20627_, _20626_, _20617_);
  nand (_20628_, _20627_, _20611_);
  nand (_20629_, _20628_, _19135_);
  nand (_08523_, _20629_, _19624_);
  nand (_20630_, _20168_, _18962_);
  nand (_20631_, _20172_, _18957_);
  nand (_20632_, _20631_, _20630_);
  nand (_20634_, _20632_, _19139_);
  not (_20635_, _20162_);
  nor (_20636_, _20635_, _18957_);
  not (_20637_, _20158_);
  nor (_20638_, _20637_, _18962_);
  nor (_20639_, _20638_, _20636_);
  nor (_20640_, _20639_, _19104_);
  nand (_20641_, _20186_, _18962_);
  nand (_20642_, _20181_, _18957_);
  nand (_20643_, _20642_, _20641_);
  nand (_20645_, _20643_, _19098_);
  nand (_20646_, _20192_, _18962_);
  nand (_20647_, _20196_, _18957_);
  nand (_20648_, _20647_, _20646_);
  nand (_20649_, _20648_, _19154_);
  nand (_20650_, _20649_, _20645_);
  nor (_20651_, _20650_, _20640_);
  nand (_20652_, _20651_, _20634_);
  nand (_20653_, _20652_, _19135_);
  nand (_08528_, _20653_, _19646_);
  nand (_20654_, _20218_, _18962_);
  nand (_20655_, _20222_, _18957_);
  nand (_20656_, _20655_, _20654_);
  nand (_20657_, _20656_, _19139_);
  not (_20658_, _20211_);
  nor (_20659_, _20658_, _18957_);
  not (_20660_, _20207_);
  nor (_20661_, _20660_, _18962_);
  nor (_20662_, _20661_, _20659_);
  nor (_20663_, _20662_, _19104_);
  nand (_20664_, _20235_, _18962_);
  nand (_20665_, _20231_, _18957_);
  nand (_20666_, _20665_, _20664_);
  nand (_20667_, _20666_, _19098_);
  nand (_20668_, _20241_, _18962_);
  nand (_20669_, _20245_, _18957_);
  nand (_20670_, _20669_, _20668_);
  nand (_20671_, _20670_, _19154_);
  nand (_20672_, _20671_, _20667_);
  nor (_20673_, _20672_, _20663_);
  nand (_20675_, _20673_, _20657_);
  nand (_20676_, _20675_, _19135_);
  nand (_08533_, _20676_, _19666_);
  nand (_20677_, _20268_, _18962_);
  nand (_20678_, _20272_, _18957_);
  nand (_20679_, _20678_, _20677_);
  nand (_20680_, _20679_, _19139_);
  not (_20681_, _20261_);
  nor (_20682_, _20681_, _18957_);
  not (_20683_, _20257_);
  nor (_20685_, _20683_, _18962_);
  nor (_20686_, _20685_, _20682_);
  nor (_20687_, _20686_, _19104_);
  nand (_20688_, _20284_, _18962_);
  nand (_20689_, _20280_, _18957_);
  nand (_20690_, _20689_, _20688_);
  nand (_20691_, _20690_, _19098_);
  nand (_20692_, _20290_, _18962_);
  nand (_20693_, _20294_, _18957_);
  nand (_20694_, _20693_, _20692_);
  nand (_20695_, _20694_, _19154_);
  nand (_20696_, _20695_, _20691_);
  nor (_20697_, _20696_, _20687_);
  nand (_20698_, _20697_, _20680_);
  nand (_20699_, _20698_, _19135_);
  nand (_08538_, _20699_, _19688_);
  nand (_20700_, _20317_, _18962_);
  nand (_20701_, _20321_, _18957_);
  nand (_20702_, _20701_, _20700_);
  nand (_20703_, _20702_, _19139_);
  not (_20704_, _20311_);
  nor (_20705_, _20704_, _18957_);
  not (_20706_, _20306_);
  nor (_20707_, _20706_, _18962_);
  nor (_20708_, _20707_, _20705_);
  nor (_20709_, _20708_, _19104_);
  nand (_20710_, _20329_, _18962_);
  nand (_20711_, _20333_, _18957_);
  nand (_20712_, _20711_, _20710_);
  nand (_20713_, _20712_, _19098_);
  nand (_20715_, _20344_, _18962_);
  nand (_20716_, _20340_, _18957_);
  nand (_20717_, _20716_, _20715_);
  nand (_20718_, _20717_, _19154_);
  nand (_20719_, _20718_, _20713_);
  nor (_20720_, _20719_, _20709_);
  nand (_20721_, _20720_, _20703_);
  nand (_20722_, _20721_, _19135_);
  nand (_08543_, _20722_, _19708_);
  nand (_20723_, _20366_, _18962_);
  nand (_20725_, _20370_, _18957_);
  nand (_20726_, _20725_, _20723_);
  nand (_20727_, _20726_, _19139_);
  not (_20728_, _20360_);
  nor (_20729_, _20728_, _18957_);
  not (_20730_, _20356_);
  nor (_20731_, _20730_, _18962_);
  nor (_20732_, _20731_, _20729_);
  nor (_20733_, _20732_, _19104_);
  nand (_20734_, _20383_, _18962_);
  nand (_20735_, _20378_, _18957_);
  nand (_20736_, _20735_, _20734_);
  nand (_20737_, _20736_, _19098_);
  nand (_20738_, _20389_, _18962_);
  nand (_20739_, _20394_, _18957_);
  nand (_20740_, _20739_, _20738_);
  nand (_20741_, _20740_, _19154_);
  nand (_20742_, _20741_, _20737_);
  nor (_20743_, _20742_, _20733_);
  nand (_20744_, _20743_, _20727_);
  nand (_20745_, _20744_, _19135_);
  nand (_08548_, _20745_, _19731_);
  nand (_20746_, _20415_, _18962_);
  nand (_20747_, _20419_, _18957_);
  nand (_20748_, _20747_, _20746_);
  nand (_20749_, _20748_, _19139_);
  not (_20750_, _20409_);
  nor (_20751_, _20750_, _18957_);
  not (_20752_, _20405_);
  nor (_20753_, _20752_, _18962_);
  nor (_20755_, _20753_, _20751_);
  nor (_20756_, _20755_, _19104_);
  nand (_20757_, _20433_, _18962_);
  nand (_20758_, _20428_, _18957_);
  nand (_20759_, _20758_, _20757_);
  nand (_20760_, _20759_, _19098_);
  nand (_20761_, _20439_, _18962_);
  nand (_20762_, _20443_, _18957_);
  nand (_20763_, _20762_, _20761_);
  nand (_20764_, _20763_, _19154_);
  nand (_20766_, _20764_, _20760_);
  nor (_20767_, _20766_, _20756_);
  nand (_20768_, _20767_, _20749_);
  nand (_20769_, _20768_, _19135_);
  nand (_08553_, _20769_, _19751_);
  nand (_20770_, _19609_, _19590_);
  nor (_20771_, _19590_, _08696_);
  nor (_20772_, _20771_, _19593_);
  nand (_20773_, _20772_, _20770_);
  nand (_20774_, _19615_, _19593_);
  nand (_20775_, _20774_, _20773_);
  nor (_20776_, _20775_, _19589_);
  nor (_20777_, _19620_, _19600_);
  nor (_20778_, _20777_, _20776_);
  nor (_20779_, _20778_, _19588_);
  nor (_20780_, _19625_, _19605_);
  nor (_09144_, _20780_, _20779_);
  nand (_20781_, _19629_, _19590_);
  nor (_20782_, _19590_, _08702_);
  nor (_20783_, _20782_, _19593_);
  nand (_20784_, _20783_, _20781_);
  nand (_20785_, _19636_, _19593_);
  nand (_20786_, _20785_, _20784_);
  nor (_20787_, _20786_, _19589_);
  nor (_20788_, _19641_, _19600_);
  nor (_20789_, _20788_, _20787_);
  nor (_20790_, _20789_, _19588_);
  nor (_20791_, _19647_, _19605_);
  nor (_09147_, _20791_, _20790_);
  nor (_20792_, _19662_, _19600_);
  nand (_20794_, _19651_, _19590_);
  nor (_20795_, _19590_, _08707_);
  nor (_20796_, _20795_, _19593_);
  nand (_20797_, _20796_, _20794_);
  nand (_20798_, _19657_, _19593_);
  nand (_20799_, _20798_, _20797_);
  nor (_20800_, _20799_, _19589_);
  nor (_20801_, _20800_, _20792_);
  nor (_20802_, _20801_, _19588_);
  nor (_20803_, _19667_, _19605_);
  nor (_09150_, _20803_, _20802_);
  nand (_20805_, _19671_, _19590_);
  nor (_20806_, _19590_, _08711_);
  nor (_20807_, _20806_, _19593_);
  nand (_20808_, _20807_, _20805_);
  nand (_20809_, _19678_, _19593_);
  nand (_20810_, _20809_, _20808_);
  nor (_20811_, _20810_, _19589_);
  nor (_20812_, _19684_, _19600_);
  nor (_20813_, _20812_, _20811_);
  nor (_20814_, _20813_, _19588_);
  nor (_20815_, _19689_, _19605_);
  nor (_09153_, _20815_, _20814_);
  nand (_20816_, _19693_, _19590_);
  nor (_20817_, _19590_, _08556_);
  nor (_20818_, _20817_, _19593_);
  nand (_20819_, _20818_, _20816_);
  nand (_20820_, _19699_, _19593_);
  nand (_20821_, _20820_, _20819_);
  nor (_20822_, _20821_, _19589_);
  nor (_20823_, _19704_, _19600_);
  nor (_20824_, _20823_, _20822_);
  nor (_20825_, _20824_, _19588_);
  nor (_20826_, _19709_, _19605_);
  nor (_09156_, _20826_, _20825_);
  nand (_20827_, _19715_, _19590_);
  nor (_20828_, _19590_, _08729_);
  nor (_20829_, _20828_, _19593_);
  nand (_20830_, _20829_, _20827_);
  nand (_20831_, _19721_, _19593_);
  nand (_20833_, _20831_, _20830_);
  nor (_20834_, _20833_, _19589_);
  nor (_20835_, _19727_, _19600_);
  nor (_20836_, _20835_, _20834_);
  nor (_20837_, _20836_, _19588_);
  nor (_20838_, _19732_, _19605_);
  nor (_09160_, _20838_, _20837_);
  nand (_20839_, _19736_, _19590_);
  nor (_20840_, _19590_, _08734_);
  nor (_20841_, _20840_, _19593_);
  nand (_20843_, _20841_, _20839_);
  nand (_20844_, _19742_, _19593_);
  nand (_20845_, _20844_, _20843_);
  nor (_20846_, _20845_, _19589_);
  nor (_20847_, _19747_, _19600_);
  nor (_20848_, _20847_, _20846_);
  nor (_20849_, _20848_, _19588_);
  nor (_20850_, _19752_, _19605_);
  nor (_09163_, _20850_, _20849_);
  nand (_20851_, _19609_, _19573_);
  nor (_20852_, _19573_, _08567_);
  nor (_20853_, _20852_, _19575_);
  nand (_20854_, _20853_, _20851_);
  nand (_20855_, _19615_, _19575_);
  nand (_20856_, _20855_, _20854_);
  nor (_20857_, _20856_, _19572_);
  nor (_20858_, _19582_, _08469_);
  nor (_20859_, _20858_, _20857_);
  nor (_20860_, _20859_, _19571_);
  nor (_20861_, _19625_, _19586_);
  nor (_09180_, _20861_, _20860_);
  nand (_20862_, _19629_, _19573_);
  nor (_20863_, _19573_, _08811_);
  nor (_20864_, _20863_, _19575_);
  nand (_20865_, _20864_, _20862_);
  nand (_20866_, _19636_, _19575_);
  nand (_20867_, _20866_, _20865_);
  nor (_20868_, _20867_, _19572_);
  nor (_20869_, _19582_, _08474_);
  nor (_20870_, _20869_, _20868_);
  nor (_20872_, _20870_, _19571_);
  nor (_20873_, _19647_, _19586_);
  nor (_09183_, _20873_, _20872_);
  nand (_20874_, _19651_, _19573_);
  nor (_20875_, _19573_, _08816_);
  nor (_20876_, _20875_, _19575_);
  nand (_20877_, _20876_, _20874_);
  nand (_20878_, _19657_, _19575_);
  nand (_20879_, _20878_, _20877_);
  nor (_20880_, _20879_, _19572_);
  nor (_20882_, _19582_, _08479_);
  nor (_20883_, _20882_, _20880_);
  nor (_20884_, _20883_, _19571_);
  nor (_20885_, _19667_, _19586_);
  nor (_09186_, _20885_, _20884_);
  nand (_20886_, _19671_, _19573_);
  nor (_20887_, _19573_, _08820_);
  nor (_20888_, _20887_, _19575_);
  nand (_20889_, _20888_, _20886_);
  nand (_20890_, _19678_, _19575_);
  nand (_20891_, _20890_, _20889_);
  nor (_20892_, _20891_, _19572_);
  nor (_20893_, _19582_, _08484_);
  nor (_20894_, _20893_, _20892_);
  nor (_20895_, _20894_, _19571_);
  nor (_20896_, _19689_, _19586_);
  nor (_09189_, _20896_, _20895_);
  nand (_20897_, _19693_, _19573_);
  nor (_20898_, _19573_, _08827_);
  nor (_20899_, _20898_, _19575_);
  nand (_20900_, _20899_, _20897_);
  nand (_20901_, _19699_, _19575_);
  nand (_20902_, _20901_, _20900_);
  nor (_20903_, _20902_, _19572_);
  nor (_20904_, _19582_, _08489_);
  nor (_20905_, _20904_, _20903_);
  nor (_20906_, _20905_, _19571_);
  nor (_20907_, _19709_, _19586_);
  nor (_09192_, _20907_, _20906_);
  nand (_20908_, _19715_, _19573_);
  nor (_20910_, _19573_, _08832_);
  nor (_20911_, _20910_, _19575_);
  nand (_20912_, _20911_, _20908_);
  nand (_20913_, _19721_, _19575_);
  nand (_20914_, _20913_, _20912_);
  nor (_20915_, _20914_, _19572_);
  nor (_20916_, _19582_, _08494_);
  nor (_20917_, _20916_, _20915_);
  nor (_20918_, _20917_, _19571_);
  nor (_20919_, _19732_, _19586_);
  nor (_09195_, _20919_, _20918_);
  nand (_20921_, _19736_, _19573_);
  nor (_20922_, _19573_, _08837_);
  nor (_20923_, _20922_, _19575_);
  nand (_20924_, _20923_, _20921_);
  nand (_20925_, _19742_, _19575_);
  nand (_20926_, _20925_, _20924_);
  nor (_20927_, _20926_, _19572_);
  nor (_20928_, _19582_, _08499_);
  nor (_20929_, _20928_, _20927_);
  nor (_20932_, _20929_, _19571_);
  nor (_20933_, _19752_, _19586_);
  nor (_09198_, _20933_, _20932_);
  nor (_20934_, _19620_, _19556_);
  not (_20935_, _19557_);
  nor (_20936_, _19608_, _20935_);
  not (_20937_, _19559_);
  nand (_20938_, _20935_, _19768_);
  nand (_20939_, _20938_, _20937_);
  nor (_20940_, _20939_, _20936_);
  nand (_20941_, _19615_, _19559_);
  nand (_20942_, _20941_, _19556_);
  nor (_20943_, _20942_, _20940_);
  nor (_20944_, _20943_, _20934_);
  nor (_20945_, _20944_, _19553_);
  nor (_20946_, _19625_, _19554_);
  nor (_09216_, _20946_, _20945_);
  nor (_20947_, _19641_, _19556_);
  nor (_20948_, _19628_, _20935_);
  not (_20949_, _08809_);
  nand (_20951_, _20935_, _20949_);
  nand (_20952_, _20951_, _20937_);
  nor (_20953_, _20952_, _20948_);
  nand (_20954_, _19636_, _19559_);
  nand (_20955_, _20954_, _19556_);
  nor (_20956_, _20955_, _20953_);
  nor (_20957_, _20956_, _20947_);
  nor (_20958_, _20957_, _19553_);
  nor (_20959_, _19647_, _19554_);
  nor (_09219_, _20959_, _20958_);
  nand (_20961_, _19651_, _19557_);
  nor (_20962_, _19557_, _08814_);
  nor (_20963_, _20962_, _19559_);
  nand (_20964_, _20963_, _20961_);
  nand (_20965_, _19657_, _19559_);
  nand (_20966_, _20965_, _20964_);
  nand (_20967_, _20966_, _19556_);
  nand (_20968_, _19662_, _19555_);
  nand (_20969_, _20968_, _20967_);
  nand (_20970_, _20969_, _19554_);
  nand (_20971_, _19667_, _19553_);
  nand (_09222_, _20971_, _20970_);
  nand (_20972_, _19671_, _19557_);
  nor (_20973_, _19557_, _08818_);
  nor (_20974_, _20973_, _19559_);
  nand (_20975_, _20974_, _20972_);
  nand (_20976_, _19678_, _19559_);
  nand (_20977_, _20976_, _20975_);
  nand (_20978_, _20977_, _19556_);
  nand (_20979_, _19684_, _19555_);
  nand (_20980_, _20979_, _20978_);
  nand (_20981_, _20980_, _19554_);
  nand (_20982_, _19689_, _19553_);
  nand (_09225_, _20982_, _20981_);
  nor (_20983_, _19704_, _19556_);
  nor (_20984_, _19692_, _20935_);
  not (_20985_, _08825_);
  nand (_20986_, _20935_, _20985_);
  nand (_20987_, _20986_, _20937_);
  nor (_20988_, _20987_, _20984_);
  nand (_20990_, _19699_, _19559_);
  nand (_20991_, _20990_, _19556_);
  nor (_20992_, _20991_, _20988_);
  nor (_20993_, _20992_, _20983_);
  nor (_20994_, _20993_, _19553_);
  nor (_20995_, _19709_, _19554_);
  nor (_09228_, _20995_, _20994_);
  nand (_20996_, _19715_, _19557_);
  nor (_20997_, _19557_, _08830_);
  nor (_20998_, _20997_, _19559_);
  nand (_21000_, _20998_, _20996_);
  nand (_21001_, _19721_, _19559_);
  nand (_21002_, _21001_, _21000_);
  nand (_21003_, _21002_, _19556_);
  nand (_21004_, _19727_, _19555_);
  nand (_21005_, _21004_, _21003_);
  nand (_21006_, _21005_, _19554_);
  nand (_21007_, _19732_, _19553_);
  nand (_09231_, _21007_, _21006_);
  nor (_21008_, _19747_, _19556_);
  nor (_21009_, _19735_, _20935_);
  not (_21010_, _08835_);
  nand (_21011_, _20935_, _21010_);
  nand (_21012_, _21011_, _20937_);
  nor (_21013_, _21012_, _21009_);
  nand (_21014_, _19742_, _19559_);
  nand (_21015_, _21014_, _19556_);
  nor (_21016_, _21015_, _21013_);
  nor (_21017_, _21016_, _21008_);
  nor (_21018_, _21017_, _19553_);
  nor (_21019_, _19752_, _19554_);
  nor (_09234_, _21019_, _21018_);
  nor (_21020_, _19615_, _19533_);
  nor (_21021_, _19609_, _19539_);
  not (_21022_, _08849_);
  nor (_21023_, _19538_, _21022_);
  nor (_21024_, _21023_, _21021_);
  nand (_21025_, _21024_, _19533_);
  nand (_21026_, _21025_, _19536_);
  nor (_21027_, _21026_, _21020_);
  nand (_21029_, _19620_, _19535_);
  nand (_21030_, _21029_, _19547_);
  nor (_21031_, _21030_, _21027_);
  nor (_21032_, _19625_, _19547_);
  nor (_09251_, _21032_, _21031_);
  nor (_21033_, _19629_, _19539_);
  not (_21034_, _08854_);
  nor (_21035_, _19538_, _21034_);
  nor (_21036_, _21035_, _21033_);
  nor (_21037_, _21036_, _19532_);
  not (_21039_, _19636_);
  nor (_21040_, _21039_, _19533_);
  nor (_21041_, _21040_, _21037_);
  nor (_21042_, _21041_, _19535_);
  nand (_21043_, _19641_, _19535_);
  nand (_21044_, _21043_, _19547_);
  nor (_21045_, _21044_, _21042_);
  nor (_21046_, _19647_, _19547_);
  nor (_09254_, _21046_, _21045_);
  nor (_21047_, _19651_, _19539_);
  not (_21048_, _08861_);
  nor (_21049_, _19538_, _21048_);
  nor (_21050_, _21049_, _21047_);
  nor (_21051_, _21050_, _19532_);
  not (_21052_, _19657_);
  nor (_21053_, _21052_, _19533_);
  nor (_21054_, _21053_, _21051_);
  nor (_21055_, _21054_, _19535_);
  nand (_21056_, _19662_, _19535_);
  nand (_21057_, _21056_, _19547_);
  nor (_21058_, _21057_, _21055_);
  nor (_21059_, _19667_, _19547_);
  nor (_09257_, _21059_, _21058_);
  nor (_21060_, _19671_, _19539_);
  not (_21061_, _08866_);
  nor (_21062_, _19538_, _21061_);
  nor (_21063_, _21062_, _21060_);
  nor (_21064_, _21063_, _19532_);
  not (_21065_, _19678_);
  nor (_21066_, _21065_, _19533_);
  nor (_21068_, _21066_, _21064_);
  nor (_21069_, _21068_, _19535_);
  nand (_21070_, _19684_, _19535_);
  nand (_21071_, _21070_, _19547_);
  nor (_21072_, _21071_, _21069_);
  nor (_21073_, _19689_, _19547_);
  nor (_09261_, _21073_, _21072_);
  nor (_21074_, _19693_, _19539_);
  not (_21075_, _08878_);
  nor (_21076_, _19538_, _21075_);
  nor (_21078_, _21076_, _21074_);
  nor (_21079_, _21078_, _19532_);
  not (_21080_, _19699_);
  nor (_21081_, _21080_, _19533_);
  nor (_21082_, _21081_, _21079_);
  nor (_21083_, _21082_, _19535_);
  nand (_21084_, _19704_, _19535_);
  nand (_21085_, _21084_, _19547_);
  nor (_21086_, _21085_, _21083_);
  nor (_21087_, _19709_, _19547_);
  nor (_09264_, _21087_, _21086_);
  nor (_21088_, _19721_, _19533_);
  nor (_21089_, _19715_, _19539_);
  not (_21090_, _08573_);
  nor (_21091_, _19538_, _21090_);
  nor (_21092_, _21091_, _21089_);
  nand (_21093_, _21092_, _19533_);
  nand (_21094_, _21093_, _19536_);
  nor (_21095_, _21094_, _21088_);
  nand (_21096_, _19727_, _19535_);
  nand (_21097_, _21096_, _19547_);
  nor (_21098_, _21097_, _21095_);
  nor (_21099_, _19732_, _19547_);
  nor (_09267_, _21099_, _21098_);
  nor (_21100_, _19742_, _19533_);
  nor (_21101_, _19736_, _19539_);
  not (_21102_, _08898_);
  nor (_21103_, _19538_, _21102_);
  nor (_21104_, _21103_, _21101_);
  nand (_21105_, _21104_, _19533_);
  nand (_21107_, _21105_, _19536_);
  nor (_21108_, _21107_, _21100_);
  nand (_21109_, _19747_, _19535_);
  nand (_21110_, _21109_, _19547_);
  nor (_21111_, _21110_, _21108_);
  nor (_21112_, _19752_, _19547_);
  nor (_09270_, _21112_, _21111_);
  not (_21113_, _08847_);
  nor (_21114_, _19516_, _21113_);
  nor (_21115_, _19609_, _19518_);
  nor (_21117_, _21115_, _21114_);
  nor (_21118_, _21117_, _19514_);
  nand (_21119_, _19615_, _19514_);
  nand (_21120_, _21119_, _19524_);
  nor (_21121_, _21120_, _21118_);
  nor (_21122_, _19620_, _19524_);
  nor (_21123_, _21122_, _21121_);
  nand (_21124_, _21123_, _19513_);
  nand (_21125_, _19625_, _19511_);
  nand (_09287_, _21125_, _21124_);
  not (_21126_, _08852_);
  nor (_21127_, _19516_, _21126_);
  nor (_21128_, _19629_, _19518_);
  nor (_21129_, _21128_, _21127_);
  nor (_21130_, _21129_, _19514_);
  nand (_21131_, _19636_, _19514_);
  nand (_21132_, _21131_, _19524_);
  nor (_21133_, _21132_, _21130_);
  nor (_21134_, _19641_, _19524_);
  nor (_21135_, _21134_, _21133_);
  nand (_21136_, _21135_, _19513_);
  nand (_21137_, _19647_, _19511_);
  nand (_09290_, _21137_, _21136_);
  not (_21138_, _08859_);
  nor (_21139_, _19516_, _21138_);
  nor (_21140_, _19651_, _19518_);
  nor (_21141_, _21140_, _21139_);
  nor (_21142_, _21141_, _19514_);
  nand (_21143_, _19657_, _19514_);
  nand (_21144_, _21143_, _19524_);
  nor (_21145_, _21144_, _21142_);
  nor (_21146_, _19662_, _19524_);
  nor (_21147_, _21146_, _21145_);
  nand (_21148_, _21147_, _19513_);
  nand (_21149_, _19667_, _19511_);
  nand (_09293_, _21149_, _21148_);
  not (_21150_, _08864_);
  nor (_21151_, _19516_, _21150_);
  nor (_21152_, _19671_, _19518_);
  nor (_21153_, _21152_, _21151_);
  nor (_21155_, _21153_, _19514_);
  nand (_21156_, _19678_, _19514_);
  nand (_21157_, _21156_, _19524_);
  nor (_21158_, _21157_, _21155_);
  nor (_21159_, _19684_, _19524_);
  nor (_21160_, _21159_, _21158_);
  nand (_21161_, _21160_, _19513_);
  nand (_21162_, _19689_, _19511_);
  nand (_09296_, _21162_, _21161_);
  not (_21163_, _08876_);
  nor (_21165_, _19516_, _21163_);
  nor (_21166_, _19693_, _19518_);
  nor (_21167_, _21166_, _21165_);
  nor (_21168_, _21167_, _19514_);
  nand (_21169_, _19699_, _19514_);
  nand (_21170_, _21169_, _19524_);
  nor (_21171_, _21170_, _21168_);
  nor (_21172_, _19704_, _19524_);
  nor (_21173_, _21172_, _21171_);
  nand (_21174_, _21173_, _19513_);
  nand (_21175_, _19709_, _19511_);
  nand (_09299_, _21175_, _21174_);
  not (_21176_, _08570_);
  nor (_21177_, _19516_, _21176_);
  nor (_21178_, _19715_, _19518_);
  nor (_21179_, _21178_, _21177_);
  nor (_21180_, _21179_, _19514_);
  nand (_21181_, _19721_, _19514_);
  nand (_21182_, _21181_, _19524_);
  nor (_21183_, _21182_, _21180_);
  nor (_21184_, _19727_, _19524_);
  nor (_21185_, _21184_, _21183_);
  nand (_21186_, _21185_, _19513_);
  nand (_21187_, _19732_, _19511_);
  nand (_09302_, _21187_, _21186_);
  not (_21188_, _08895_);
  nor (_21189_, _19516_, _21188_);
  nor (_21190_, _19736_, _19518_);
  nor (_21191_, _21190_, _21189_);
  nor (_21192_, _21191_, _19514_);
  nand (_21194_, _19742_, _19514_);
  nand (_21195_, _21194_, _19524_);
  nor (_21196_, _21195_, _21192_);
  nor (_21197_, _19747_, _19524_);
  nor (_21198_, _21197_, _21196_);
  nand (_21199_, _21198_, _19513_);
  nand (_21200_, _19752_, _19511_);
  nand (_09305_, _21200_, _21199_);
  not (_21201_, _08902_);
  nor (_21202_, _19496_, _21201_);
  nor (_21204_, _19609_, _19498_);
  nor (_21205_, _21204_, _21202_);
  nor (_21206_, _21205_, _19494_);
  nor (_21207_, _19502_, _19614_);
  nor (_21208_, _21207_, _21206_);
  nor (_21209_, _21208_, _19491_);
  nand (_21210_, _19620_, _19491_);
  nand (_21211_, _21210_, _19506_);
  nor (_21212_, _21211_, _21209_);
  nor (_21213_, _19625_, _19506_);
  nor (_09324_, _21213_, _21212_);
  not (_21214_, _08907_);
  nor (_21215_, _19496_, _21214_);
  nor (_21216_, _19629_, _19498_);
  nor (_21217_, _21216_, _21215_);
  nor (_21218_, _21217_, _19494_);
  nor (_21219_, _19502_, _19635_);
  nor (_21220_, _21219_, _21218_);
  nor (_21221_, _21220_, _19491_);
  nand (_21222_, _19641_, _19491_);
  nand (_21223_, _21222_, _19506_);
  nor (_21224_, _21223_, _21221_);
  nor (_21225_, _19647_, _19506_);
  nor (_09327_, _21225_, _21224_);
  not (_21226_, _08913_);
  nor (_21227_, _19496_, _21226_);
  nor (_21228_, _19651_, _19498_);
  nor (_21229_, _21228_, _21227_);
  nor (_21230_, _21229_, _19494_);
  nor (_21231_, _19502_, _19656_);
  nor (_21233_, _21231_, _21230_);
  nor (_21234_, _21233_, _19491_);
  nand (_21235_, _19662_, _19491_);
  nand (_21236_, _21235_, _19506_);
  nor (_21237_, _21236_, _21234_);
  nor (_21238_, _19667_, _19506_);
  nor (_09330_, _21238_, _21237_);
  not (_21239_, _08918_);
  nor (_21240_, _19496_, _21239_);
  nor (_21241_, _19671_, _19498_);
  nor (_21243_, _21241_, _21240_);
  nor (_21244_, _21243_, _19494_);
  nor (_21245_, _19502_, _19677_);
  nor (_21246_, _21245_, _21244_);
  nor (_21247_, _21246_, _19491_);
  nand (_21248_, _19684_, _19491_);
  nand (_21249_, _21248_, _19506_);
  nor (_21250_, _21249_, _21247_);
  nor (_21251_, _19689_, _19506_);
  nor (_09333_, _21251_, _21250_);
  not (_21252_, _08923_);
  nor (_21253_, _19496_, _21252_);
  nor (_21254_, _19693_, _19498_);
  nor (_21255_, _21254_, _21253_);
  nor (_21256_, _21255_, _19494_);
  nor (_21257_, _19502_, _19698_);
  nor (_21258_, _21257_, _21256_);
  nor (_21259_, _21258_, _19491_);
  nand (_21260_, _19704_, _19491_);
  nand (_21261_, _21260_, _19506_);
  nor (_21262_, _21261_, _21259_);
  nor (_21263_, _19709_, _19506_);
  nor (_09336_, _21263_, _21262_);
  not (_21264_, _08928_);
  nor (_21265_, _19496_, _21264_);
  nor (_21266_, _19715_, _19498_);
  nor (_21267_, _21266_, _21265_);
  nor (_21268_, _21267_, _19494_);
  nor (_21269_, _19502_, _19720_);
  nor (_21270_, _21269_, _21268_);
  nor (_21272_, _21270_, _19491_);
  nand (_21273_, _19727_, _19491_);
  nand (_21274_, _21273_, _19506_);
  nor (_21275_, _21274_, _21272_);
  nor (_21276_, _19732_, _19506_);
  nor (_09339_, _21276_, _21275_);
  not (_21277_, _08934_);
  nor (_21278_, _19496_, _21277_);
  nor (_21279_, _19736_, _19498_);
  nor (_21280_, _21279_, _21278_);
  nor (_21282_, _21280_, _19494_);
  nor (_21283_, _19502_, _19741_);
  nor (_21284_, _21283_, _21282_);
  nor (_21285_, _21284_, _19491_);
  nand (_21286_, _19747_, _19491_);
  nand (_21287_, _21286_, _19506_);
  nor (_21288_, _21287_, _21285_);
  nor (_21289_, _19752_, _19506_);
  nor (_09342_, _21289_, _21288_);
  nor (_21290_, _19471_, _08469_);
  not (_21291_, _19476_);
  nor (_21292_, _21291_, _08395_);
  not (_21293_, _19478_);
  not (_21294_, _08900_);
  nand (_21295_, _21291_, _21294_);
  nand (_21296_, _21295_, _21293_);
  nor (_21297_, _21296_, _21292_);
  nand (_21298_, _19615_, _19478_);
  nand (_21299_, _21298_, _19471_);
  nor (_21300_, _21299_, _21297_);
  nor (_21301_, _21300_, _21290_);
  nand (_21302_, _21301_, _19468_);
  nand (_21303_, _19489_, _08520_);
  nand (_09359_, _21303_, _21302_);
  nor (_21304_, _19476_, _08905_);
  nor (_21305_, _21291_, _08400_);
  nor (_21306_, _21305_, _21304_);
  nand (_21307_, _21306_, _21293_);
  nor (_21308_, _21039_, _21293_);
  nor (_21309_, _21308_, _19473_);
  nand (_21311_, _21309_, _21307_);
  nor (_21312_, _19471_, _08474_);
  nor (_21313_, _21312_, _19489_);
  nand (_21314_, _21313_, _21311_);
  nand (_21315_, _19489_, _08525_);
  nand (_09363_, _21315_, _21314_);
  nand (_21316_, _19489_, _08530_);
  nor (_21317_, _19476_, _08911_);
  nor (_21318_, _21291_, _08405_);
  nor (_21319_, _21318_, _21317_);
  nand (_21322_, _21319_, _21293_);
  nor (_21323_, _21052_, _21293_);
  nor (_21324_, _21323_, _19473_);
  nand (_21325_, _21324_, _21322_);
  nor (_21326_, _19471_, _08479_);
  nor (_21327_, _21326_, _19489_);
  nand (_21328_, _21327_, _21325_);
  nand (_09366_, _21328_, _21316_);
  nor (_21329_, _19476_, _08916_);
  nor (_21330_, _21291_, _08410_);
  nor (_21331_, _21330_, _21329_);
  nand (_21332_, _21331_, _21293_);
  nor (_21333_, _21065_, _21293_);
  nor (_21334_, _21333_, _19473_);
  nand (_21335_, _21334_, _21332_);
  nor (_21336_, _19471_, _08484_);
  nor (_21337_, _21336_, _19489_);
  nand (_21338_, _21337_, _21335_);
  nand (_21339_, _19489_, _08535_);
  nand (_09369_, _21339_, _21338_);
  nand (_21340_, _19489_, _08540_);
  nor (_21341_, _19476_, _08921_);
  nor (_21342_, _21291_, _08414_);
  nor (_21343_, _21342_, _21341_);
  nand (_21344_, _21343_, _21293_);
  nor (_21345_, _21080_, _21293_);
  nor (_21346_, _21345_, _19473_);
  nand (_21347_, _21346_, _21344_);
  nor (_21348_, _19471_, _08489_);
  nor (_21349_, _21348_, _19489_);
  nand (_21351_, _21349_, _21347_);
  nand (_09372_, _21351_, _21340_);
  nor (_21352_, _19471_, _08494_);
  nor (_21353_, _21291_, _08418_);
  not (_21354_, _08926_);
  nand (_21355_, _21291_, _21354_);
  nand (_21356_, _21355_, _21293_);
  nor (_21357_, _21356_, _21353_);
  nand (_21358_, _19721_, _19478_);
  nand (_21359_, _21358_, _19471_);
  nor (_21361_, _21359_, _21357_);
  nor (_21362_, _21361_, _21352_);
  nand (_21363_, _21362_, _19468_);
  nand (_21364_, _19489_, _08545_);
  nand (_09375_, _21364_, _21363_);
  nor (_21365_, _19471_, _08499_);
  nor (_21366_, _21291_, _08422_);
  not (_21367_, _08932_);
  nand (_21368_, _21291_, _21367_);
  nand (_21369_, _21368_, _21293_);
  nor (_21370_, _21369_, _21366_);
  nand (_21371_, _19742_, _19478_);
  nand (_21372_, _21371_, _19471_);
  nor (_21373_, _21372_, _21370_);
  nor (_21374_, _21373_, _21365_);
  nand (_21375_, _21374_, _19468_);
  nand (_21376_, _19489_, _08550_);
  nand (_09378_, _21376_, _21375_);
  nor (_21377_, _19620_, _19462_);
  nand (_21378_, _19609_, _19453_);
  nor (_21379_, _19453_, _08938_);
  nor (_21380_, _21379_, _19455_);
  nand (_21381_, _21380_, _21378_);
  nand (_21382_, _19615_, _19455_);
  nand (_21383_, _21382_, _21381_);
  nor (_21384_, _21383_, _19452_);
  nor (_21385_, _21384_, _21377_);
  nor (_21386_, _21385_, _19451_);
  nor (_21387_, _19625_, _19466_);
  nor (_09395_, _21387_, _21386_);
  nand (_21389_, _19629_, _19453_);
  nor (_21390_, _19453_, _08944_);
  nor (_21391_, _21390_, _19455_);
  nand (_21392_, _21391_, _21389_);
  nand (_21393_, _19636_, _19455_);
  nand (_21394_, _21393_, _21392_);
  nor (_21395_, _21394_, _19452_);
  nor (_21396_, _19641_, _19462_);
  nor (_21397_, _21396_, _21395_);
  nor (_21398_, _21397_, _19451_);
  nor (_21400_, _19647_, _19466_);
  nor (_09398_, _21400_, _21398_);
  nand (_21401_, _19651_, _19453_);
  nor (_21402_, _19453_, _08952_);
  nor (_21403_, _21402_, _19455_);
  nand (_21404_, _21403_, _21401_);
  nand (_21405_, _19657_, _19455_);
  nand (_21406_, _21405_, _21404_);
  nor (_21407_, _21406_, _19452_);
  nor (_21408_, _19662_, _19462_);
  nor (_21409_, _21408_, _21407_);
  nor (_21410_, _21409_, _19451_);
  nor (_21411_, _19667_, _19466_);
  nor (_09401_, _21411_, _21410_);
  nor (_21412_, _19684_, _19462_);
  nand (_21413_, _19671_, _19453_);
  nor (_21414_, _19453_, _08517_);
  nor (_21415_, _21414_, _19455_);
  nand (_21416_, _21415_, _21413_);
  nand (_21417_, _19678_, _19455_);
  nand (_21418_, _21417_, _21416_);
  nor (_21419_, _21418_, _19452_);
  nor (_21420_, _21419_, _21412_);
  nor (_21421_, _21420_, _19451_);
  nor (_21422_, _19689_, _19466_);
  nor (_09404_, _21422_, _21421_);
  nand (_21423_, _19693_, _19453_);
  nor (_21424_, _19453_, _08971_);
  nor (_21425_, _21424_, _19455_);
  nand (_21426_, _21425_, _21423_);
  nand (_21428_, _19699_, _19455_);
  nand (_21429_, _21428_, _21426_);
  nand (_21430_, _21429_, _19462_);
  nand (_21431_, _19704_, _19452_);
  nand (_21432_, _21431_, _21430_);
  nand (_21433_, _21432_, _19466_);
  nand (_21434_, _19709_, _19451_);
  nand (_09407_, _21434_, _21433_);
  nor (_21435_, _19727_, _19462_);
  nand (_21436_, _19715_, _19453_);
  nor (_21438_, _19453_, _07607_);
  nor (_21439_, _21438_, _19455_);
  nand (_21440_, _21439_, _21436_);
  nand (_21441_, _19721_, _19455_);
  nand (_21442_, _21441_, _21440_);
  nor (_21443_, _21442_, _19452_);
  nor (_21444_, _21443_, _21435_);
  nor (_21445_, _21444_, _19451_);
  nor (_21446_, _19732_, _19466_);
  nor (_09410_, _21446_, _21445_);
  nand (_21447_, _19736_, _19453_);
  nor (_21448_, _19453_, _08982_);
  nor (_21449_, _21448_, _19455_);
  nand (_21450_, _21449_, _21447_);
  nand (_21451_, _19742_, _19455_);
  nand (_21452_, _21451_, _21450_);
  nor (_21453_, _21452_, _19452_);
  nor (_21454_, _19747_, _19462_);
  nor (_21455_, _21454_, _21453_);
  nor (_21456_, _21455_, _19451_);
  nor (_21457_, _19752_, _19466_);
  nor (_09413_, _21457_, _21456_);
  nand (_21458_, _19609_, _19437_);
  nor (_21459_, _19437_, _08936_);
  nor (_21460_, _21459_, _19439_);
  nand (_21461_, _21460_, _21458_);
  nand (_21462_, _19615_, _19439_);
  nand (_21463_, _21462_, _21461_);
  nor (_21464_, _21463_, _19434_);
  nor (_21465_, _19620_, _19435_);
  nor (_21467_, _21465_, _21464_);
  nor (_21468_, _21467_, _19433_);
  nor (_21469_, _19625_, _19449_);
  nor (_09431_, _21469_, _21468_);
  nand (_21470_, _19629_, _19437_);
  nor (_21471_, _19437_, _08942_);
  nor (_21472_, _21471_, _19439_);
  nand (_21473_, _21472_, _21470_);
  nand (_21474_, _19636_, _19439_);
  nand (_21475_, _21474_, _21473_);
  nor (_21477_, _21475_, _19434_);
  nor (_21478_, _19641_, _19435_);
  nor (_21479_, _21478_, _21477_);
  nor (_21480_, _21479_, _19433_);
  nor (_21481_, _19647_, _19449_);
  nor (_09434_, _21481_, _21480_);
  nand (_21482_, _19651_, _19437_);
  nor (_21483_, _19437_, _08950_);
  nor (_21484_, _21483_, _19439_);
  nand (_21485_, _21484_, _21482_);
  nand (_21486_, _19657_, _19439_);
  nand (_21487_, _21486_, _21485_);
  nor (_21488_, _21487_, _19434_);
  nor (_21489_, _19662_, _19435_);
  nor (_21490_, _21489_, _21488_);
  nor (_21491_, _21490_, _19433_);
  nor (_21492_, _19667_, _19449_);
  nor (_09437_, _21492_, _21491_);
  nand (_21493_, _19671_, _19437_);
  nor (_21494_, _19437_, _08515_);
  nor (_21495_, _21494_, _19439_);
  nand (_21496_, _21495_, _21493_);
  nand (_21497_, _19678_, _19439_);
  nand (_21498_, _21497_, _21496_);
  nor (_21499_, _21498_, _19434_);
  nor (_21500_, _19684_, _19435_);
  nor (_21501_, _21500_, _21499_);
  nor (_21502_, _21501_, _19433_);
  nor (_21503_, _19689_, _19449_);
  nor (_09440_, _21503_, _21502_);
  nand (_21505_, _19693_, _19437_);
  nor (_21506_, _19437_, _08969_);
  nor (_21507_, _21506_, _19439_);
  nand (_21508_, _21507_, _21505_);
  nand (_21509_, _19699_, _19439_);
  nand (_21510_, _21509_, _21508_);
  nor (_21511_, _21510_, _19434_);
  nor (_21512_, _19704_, _19435_);
  nor (_21513_, _21512_, _21511_);
  nor (_21514_, _21513_, _19433_);
  nor (_21516_, _19709_, _19449_);
  nor (_09443_, _21516_, _21514_);
  nand (_21517_, _19715_, _19437_);
  nor (_21518_, _19437_, _07605_);
  nor (_21519_, _21518_, _19439_);
  nand (_21520_, _21519_, _21517_);
  nand (_21521_, _19721_, _19439_);
  nand (_21522_, _21521_, _21520_);
  nor (_21523_, _21522_, _19434_);
  nor (_21524_, _19727_, _19435_);
  nor (_21525_, _21524_, _21523_);
  nor (_21526_, _21525_, _19433_);
  nor (_21527_, _19732_, _19449_);
  nor (_09446_, _21527_, _21526_);
  nand (_21528_, _19736_, _19437_);
  nor (_21529_, _19437_, _08980_);
  nor (_21530_, _21529_, _19439_);
  nand (_21531_, _21530_, _21528_);
  nand (_21532_, _19742_, _19439_);
  nand (_21533_, _21532_, _21531_);
  nor (_21534_, _21533_, _19434_);
  nor (_21535_, _19747_, _19435_);
  nor (_21536_, _21535_, _21534_);
  nor (_21537_, _21536_, _19433_);
  nor (_21538_, _19752_, _19449_);
  nor (_09449_, _21538_, _21537_);
  nand (_21539_, _19609_, _19417_);
  nor (_21540_, _19417_, _08988_);
  nor (_21541_, _21540_, _19419_);
  nand (_21542_, _21541_, _21539_);
  nand (_21544_, _19615_, _19419_);
  nand (_21545_, _21544_, _21542_);
  nor (_21546_, _21545_, _19416_);
  nor (_21547_, _19620_, _19426_);
  nor (_21548_, _21547_, _21546_);
  nor (_21549_, _21548_, _19415_);
  nor (_21550_, _19625_, _19430_);
  nor (_09467_, _21550_, _21549_);
  nand (_21551_, _19629_, _19417_);
  nor (_21552_, _19417_, _08995_);
  nor (_21554_, _21552_, _19419_);
  nand (_21555_, _21554_, _21551_);
  nand (_21556_, _19636_, _19419_);
  nand (_21557_, _21556_, _21555_);
  nand (_21558_, _21557_, _19426_);
  nand (_21559_, _19641_, _19416_);
  nand (_21560_, _21559_, _21558_);
  nand (_21561_, _21560_, _19430_);
  nand (_21562_, _19647_, _19415_);
  nand (_09470_, _21562_, _21561_);
  nand (_21563_, _19651_, _19417_);
  nor (_21564_, _19417_, _09000_);
  nor (_21565_, _21564_, _19419_);
  nand (_21566_, _21565_, _21563_);
  nand (_21567_, _19657_, _19419_);
  nand (_21568_, _21567_, _21566_);
  nor (_21569_, _21568_, _19416_);
  nor (_21570_, _19662_, _19426_);
  nor (_21571_, _21570_, _21569_);
  nor (_21572_, _21571_, _19415_);
  nor (_21573_, _19667_, _19430_);
  nor (_09473_, _21573_, _21572_);
  nand (_21574_, _19671_, _19417_);
  nor (_21575_, _19417_, _09005_);
  nor (_21576_, _21575_, _19419_);
  nand (_21577_, _21576_, _21574_);
  nand (_21578_, _19678_, _19419_);
  nand (_21579_, _21578_, _21577_);
  nor (_21580_, _21579_, _19416_);
  nor (_21581_, _19684_, _19426_);
  nor (_21583_, _21581_, _21580_);
  nor (_21584_, _21583_, _19415_);
  nor (_21585_, _19689_, _19430_);
  nor (_09476_, _21585_, _21584_);
  nand (_21586_, _19693_, _19417_);
  nor (_21587_, _19417_, _09012_);
  nor (_21588_, _21587_, _19419_);
  nand (_21589_, _21588_, _21586_);
  nand (_21590_, _19699_, _19419_);
  nand (_21591_, _21590_, _21589_);
  nand (_21593_, _21591_, _19426_);
  nand (_21594_, _19704_, _19416_);
  nand (_21595_, _21594_, _21593_);
  nand (_21596_, _21595_, _19430_);
  nand (_21597_, _19709_, _19415_);
  nand (_09479_, _21597_, _21596_);
  nand (_21598_, _19715_, _19417_);
  nor (_21599_, _19417_, _09018_);
  nor (_21600_, _21599_, _19419_);
  nand (_21601_, _21600_, _21598_);
  nand (_21602_, _19721_, _19419_);
  nand (_21603_, _21602_, _21601_);
  nand (_21604_, _21603_, _19426_);
  nand (_21605_, _19727_, _19416_);
  nand (_21606_, _21605_, _21604_);
  nand (_21607_, _21606_, _19430_);
  nand (_21608_, _19732_, _19415_);
  nand (_09482_, _21608_, _21607_);
  nand (_21609_, _19736_, _19417_);
  nor (_21610_, _19417_, _09023_);
  nor (_21611_, _21610_, _19419_);
  nand (_21612_, _21611_, _21609_);
  nand (_21613_, _19742_, _19419_);
  nand (_21614_, _21613_, _21612_);
  nor (_21615_, _21614_, _19416_);
  nor (_21616_, _19747_, _19426_);
  nor (_21617_, _21616_, _21615_);
  nor (_21618_, _21617_, _19415_);
  nor (_21619_, _19752_, _19430_);
  nor (_09485_, _21619_, _21618_);
  nand (_21621_, _19609_, _19400_);
  nor (_21622_, _19400_, _08986_);
  nor (_21623_, _21622_, _19404_);
  nand (_21624_, _21623_, _21621_);
  nand (_21625_, _19615_, _19404_);
  nand (_21626_, _21625_, _21624_);
  nor (_21627_, _21626_, _19395_);
  nor (_21628_, _19620_, _19396_);
  nor (_21629_, _21628_, _21627_);
  nor (_21630_, _21629_, _19391_);
  nor (_21632_, _19625_, _19413_);
  nor (_09502_, _21632_, _21630_);
  nand (_21633_, _19629_, _19400_);
  nor (_21634_, _19400_, _08993_);
  nor (_21635_, _21634_, _19404_);
  nand (_21636_, _21635_, _21633_);
  nand (_21637_, _19636_, _19404_);
  nand (_21638_, _21637_, _21636_);
  nor (_21639_, _21638_, _19395_);
  nor (_21640_, _19641_, _19396_);
  nor (_21641_, _21640_, _21639_);
  nor (_21642_, _21641_, _19391_);
  nor (_21643_, _19647_, _19413_);
  nor (_09505_, _21643_, _21642_);
  nand (_21644_, _19651_, _19400_);
  nor (_21645_, _19400_, _08998_);
  nor (_21646_, _21645_, _19404_);
  nand (_21647_, _21646_, _21644_);
  nand (_21648_, _19657_, _19404_);
  nand (_21649_, _21648_, _21647_);
  nor (_21650_, _21649_, _19395_);
  nor (_21651_, _19662_, _19396_);
  nor (_21652_, _21651_, _21650_);
  nor (_21653_, _21652_, _19391_);
  nor (_21654_, _19667_, _19413_);
  nor (_09508_, _21654_, _21653_);
  nand (_21655_, _19671_, _19400_);
  nor (_21656_, _19400_, _09003_);
  nor (_21657_, _21656_, _19404_);
  nand (_21658_, _21657_, _21655_);
  nand (_21660_, _19678_, _19404_);
  nand (_21661_, _21660_, _21658_);
  nor (_21662_, _21661_, _19395_);
  nor (_21663_, _19684_, _19396_);
  nor (_21664_, _21663_, _21662_);
  nor (_21665_, _21664_, _19391_);
  nor (_21666_, _19689_, _19413_);
  nor (_09511_, _21666_, _21665_);
  nand (_21667_, _19693_, _19400_);
  nor (_21668_, _19400_, _09010_);
  nor (_21670_, _21668_, _19404_);
  nand (_21671_, _21670_, _21667_);
  nand (_21672_, _19699_, _19404_);
  nand (_21673_, _21672_, _21671_);
  nor (_21674_, _21673_, _19395_);
  nor (_21675_, _19704_, _19396_);
  nor (_21676_, _21675_, _21674_);
  nor (_21677_, _21676_, _19391_);
  nor (_21678_, _19709_, _19413_);
  nor (_09514_, _21678_, _21677_);
  nand (_21679_, _19715_, _19400_);
  nor (_21680_, _19400_, _09016_);
  nor (_21681_, _21680_, _19404_);
  nand (_21682_, _21681_, _21679_);
  nand (_21683_, _19721_, _19404_);
  nand (_21684_, _21683_, _21682_);
  nor (_21685_, _21684_, _19395_);
  nor (_21686_, _19727_, _19396_);
  nor (_21687_, _21686_, _21685_);
  nor (_21688_, _21687_, _19391_);
  nor (_21689_, _19732_, _19413_);
  nor (_09518_, _21689_, _21688_);
  nand (_21690_, _19736_, _19400_);
  nor (_21691_, _19400_, _09021_);
  nor (_21692_, _21691_, _19404_);
  nand (_21693_, _21692_, _21690_);
  nand (_21694_, _19742_, _19404_);
  nand (_21695_, _21694_, _21693_);
  nor (_21696_, _21695_, _19395_);
  nor (_21697_, _19747_, _19396_);
  nor (_21699_, _21697_, _21696_);
  nor (_21700_, _21699_, _19391_);
  nor (_21701_, _19752_, _19413_);
  nor (_09521_, _21701_, _21700_);
  nand (_21702_, _19372_, _08512_);
  nand (_21703_, _19608_, _19371_);
  nand (_21704_, _21703_, _21702_);
  nor (_21705_, _21704_, _19370_);
  nand (_21706_, _19370_, _19614_);
  nand (_21707_, _21706_, _19380_);
  nor (_21710_, _21707_, _21705_);
  nand (_21711_, _19620_, _19379_);
  nand (_21712_, _21711_, _19384_);
  nor (_21713_, _21712_, _21710_);
  nor (_21714_, _19625_, _19384_);
  nor (_09538_, _21714_, _21713_);
  nand (_21715_, _19372_, _09034_);
  nand (_21716_, _19628_, _19371_);
  nand (_21717_, _21716_, _21715_);
  nor (_21718_, _21717_, _19370_);
  nand (_21719_, _19370_, _19635_);
  nand (_21720_, _21719_, _19380_);
  nor (_21721_, _21720_, _21718_);
  nand (_21722_, _19641_, _19379_);
  nand (_21723_, _21722_, _19384_);
  nor (_21724_, _21723_, _21721_);
  nor (_21725_, _19647_, _19384_);
  nor (_09541_, _21725_, _21724_);
  nand (_21726_, _19372_, _09039_);
  nand (_21727_, _19650_, _19371_);
  nand (_21728_, _21727_, _21726_);
  nor (_21729_, _21728_, _19370_);
  nand (_21730_, _19370_, _19656_);
  nand (_21731_, _21730_, _19380_);
  nor (_21732_, _21731_, _21729_);
  nand (_21733_, _19662_, _19379_);
  nand (_21734_, _21733_, _19384_);
  nor (_21735_, _21734_, _21732_);
  nor (_21736_, _19667_, _19384_);
  nor (_09544_, _21736_, _21735_);
  nand (_21738_, _19372_, _09045_);
  nand (_21739_, _19670_, _19371_);
  nand (_21740_, _21739_, _21738_);
  nor (_21741_, _21740_, _19370_);
  nand (_21742_, _19370_, _19677_);
  nand (_21743_, _21742_, _19380_);
  nor (_21744_, _21743_, _21741_);
  nand (_21745_, _19684_, _19379_);
  nand (_21746_, _21745_, _19384_);
  nor (_21747_, _21746_, _21744_);
  nor (_21749_, _19689_, _19384_);
  nor (_09547_, _21749_, _21747_);
  not (_21750_, _09050_);
  nand (_21751_, _19372_, _21750_);
  nand (_21752_, _19693_, _19371_);
  nand (_21753_, _21752_, _21751_);
  nand (_21754_, _21753_, _19369_);
  nand (_21755_, _19370_, _19698_);
  nand (_21756_, _21755_, _21754_);
  nand (_21757_, _21756_, _19380_);
  not (_21758_, _19384_);
  nor (_21759_, _19704_, _19380_);
  nor (_21760_, _21759_, _21758_);
  nand (_21761_, _21760_, _21757_);
  nand (_21762_, _19709_, _21758_);
  nand (_09550_, _21762_, _21761_);
  not (_21763_, _09056_);
  nand (_21764_, _19372_, _21763_);
  nand (_21765_, _19715_, _19371_);
  nand (_21766_, _21765_, _21764_);
  nand (_21767_, _21766_, _19369_);
  nand (_21768_, _19370_, _19720_);
  nand (_21769_, _21768_, _21767_);
  nand (_21770_, _21769_, _19380_);
  nor (_21771_, _19727_, _19380_);
  nor (_21772_, _21771_, _21758_);
  nand (_21773_, _21772_, _21770_);
  nand (_21774_, _19732_, _21758_);
  nand (_09553_, _21774_, _21773_);
  not (_21775_, _08578_);
  nand (_21776_, _19372_, _21775_);
  nand (_21777_, _19736_, _19371_);
  nand (_21778_, _21777_, _21776_);
  nand (_21779_, _21778_, _19369_);
  nand (_21780_, _19370_, _19741_);
  nand (_21781_, _21780_, _21779_);
  nand (_21782_, _21781_, _19380_);
  nor (_21783_, _19747_, _19380_);
  nor (_21784_, _21783_, _21758_);
  nand (_21785_, _21784_, _21782_);
  nand (_21787_, _19752_, _21758_);
  nand (_09556_, _21787_, _21785_);
  not (_21788_, _08510_);
  nor (_21789_, _19348_, _21788_);
  nor (_21790_, _19609_, _19349_);
  nor (_21791_, _21790_, _21789_);
  nor (_21792_, _21791_, _19346_);
  nand (_21793_, _19615_, _19344_);
  nand (_21794_, _21793_, _19359_);
  nor (_21795_, _21794_, _21792_);
  nor (_21797_, _19620_, _19359_);
  nor (_21798_, _21797_, _21795_);
  nand (_21799_, _21798_, _19343_);
  nand (_21800_, _19625_, _19342_);
  nand (_09574_, _21800_, _21799_);
  nor (_21801_, _19629_, _19349_);
  not (_21802_, _09032_);
  nor (_21803_, _19348_, _21802_);
  nor (_21804_, _21803_, _21801_);
  nor (_21805_, _21804_, _19346_);
  nand (_21806_, _19636_, _19344_);
  nand (_21807_, _21806_, _19359_);
  nor (_21808_, _21807_, _21805_);
  nor (_21809_, _19641_, _19359_);
  nor (_21810_, _21809_, _21808_);
  nand (_21811_, _21810_, _19343_);
  nand (_21812_, _19647_, _19342_);
  nand (_09577_, _21812_, _21811_);
  nor (_21813_, _19651_, _19349_);
  not (_21814_, _09037_);
  nor (_21815_, _19348_, _21814_);
  nor (_21816_, _21815_, _21813_);
  nor (_21817_, _21816_, _19346_);
  nand (_21818_, _19657_, _19344_);
  nand (_21819_, _21818_, _19359_);
  nor (_21820_, _21819_, _21817_);
  nor (_21821_, _19662_, _19359_);
  nor (_21822_, _21821_, _21820_);
  nand (_21823_, _21822_, _19343_);
  nand (_21824_, _19667_, _19342_);
  nand (_09580_, _21824_, _21823_);
  nor (_21826_, _19671_, _19349_);
  not (_21827_, _09043_);
  nor (_21828_, _19348_, _21827_);
  nor (_21829_, _21828_, _21826_);
  nor (_21830_, _21829_, _19346_);
  nand (_21831_, _19346_, _08441_);
  nand (_21832_, _21831_, _19359_);
  nor (_21833_, _21832_, _21830_);
  nor (_21834_, _19684_, _19359_);
  nor (_21836_, _21834_, _21833_);
  nand (_21837_, _21836_, _19343_);
  nand (_21838_, _19689_, _19342_);
  nand (_09583_, _21838_, _21837_);
  nor (_21839_, _19693_, _19349_);
  not (_21840_, _09048_);
  nor (_21841_, _19348_, _21840_);
  nor (_21842_, _21841_, _21839_);
  nor (_21843_, _21842_, _19346_);
  nand (_21844_, _19699_, _19344_);
  nand (_21845_, _21844_, _19359_);
  nor (_21846_, _21845_, _21843_);
  nor (_21847_, _19704_, _19359_);
  nor (_21848_, _21847_, _21846_);
  nand (_21849_, _21848_, _19343_);
  nand (_21850_, _19709_, _19342_);
  nand (_09586_, _21850_, _21849_);
  not (_21851_, _09054_);
  nor (_21852_, _19348_, _21851_);
  nor (_21853_, _19715_, _19349_);
  nor (_21854_, _21853_, _21852_);
  nor (_21855_, _21854_, _19346_);
  nand (_21856_, _19721_, _19344_);
  nand (_21857_, _21856_, _19359_);
  nor (_21858_, _21857_, _21855_);
  nor (_21859_, _19727_, _19359_);
  nor (_21860_, _21859_, _21858_);
  nand (_21861_, _21860_, _19343_);
  nand (_21862_, _19732_, _19342_);
  nand (_09589_, _21862_, _21861_);
  nor (_21864_, _19736_, _19349_);
  not (_21865_, _08576_);
  nor (_21866_, _19348_, _21865_);
  nor (_21867_, _21866_, _21864_);
  nor (_21868_, _21867_, _19346_);
  nand (_21869_, _19742_, _19344_);
  nand (_21870_, _21869_, _19359_);
  nor (_21871_, _21870_, _21868_);
  nor (_21872_, _19747_, _19359_);
  nor (_21873_, _21872_, _21871_);
  nand (_21875_, _21873_, _19343_);
  nand (_21876_, _19752_, _19342_);
  nand (_09592_, _21876_, _21875_);
  nand (_21877_, _19324_, _09060_);
  nand (_21878_, _19608_, _19323_);
  nand (_21879_, _21878_, _21877_);
  nor (_21880_, _21879_, _19329_);
  nand (_21881_, _19329_, _19614_);
  nand (_21882_, _21881_, _19314_);
  nor (_21883_, _21882_, _21880_);
  nand (_21884_, _19620_, _19313_);
  nand (_21885_, _21884_, _19334_);
  nor (_21886_, _21885_, _21883_);
  nor (_21887_, _19625_, _19334_);
  nor (_09609_, _21887_, _21886_);
  nand (_21888_, _19324_, _08506_);
  nand (_21889_, _19628_, _19323_);
  nand (_21890_, _21889_, _21888_);
  nor (_21891_, _21890_, _19329_);
  nand (_21892_, _19329_, _19635_);
  nand (_21893_, _21892_, _19314_);
  nor (_21894_, _21893_, _21891_);
  nand (_21895_, _19641_, _19313_);
  nand (_21896_, _21895_, _19334_);
  nor (_21897_, _21896_, _21894_);
  nor (_21898_, _19647_, _19334_);
  nor (_09612_, _21898_, _21897_);
  nand (_21899_, _19324_, _09644_);
  nand (_21900_, _19650_, _19323_);
  nand (_21901_, _21900_, _21899_);
  nor (_21903_, _21901_, _19329_);
  nand (_21904_, _19329_, _19656_);
  nand (_21905_, _21904_, _19314_);
  nor (_21906_, _21905_, _21903_);
  nand (_21907_, _19662_, _19313_);
  nand (_21908_, _21907_, _19334_);
  nor (_21909_, _21908_, _21906_);
  nor (_21910_, _19667_, _19334_);
  nor (_09615_, _21910_, _21909_);
  not (_21911_, _09646_);
  nand (_21913_, _19324_, _21911_);
  nand (_21914_, _19671_, _19323_);
  nand (_21915_, _21914_, _21913_);
  nand (_21916_, _21915_, _19316_);
  nor (_21917_, _19316_, _08441_);
  nor (_21918_, _21917_, _19313_);
  nand (_21919_, _21918_, _21916_);
  nand (_21920_, _19684_, _19313_);
  nand (_21921_, _21920_, _21919_);
  nor (_21922_, _21921_, _19335_);
  nor (_21923_, _19689_, _19334_);
  nor (_09619_, _21923_, _21922_);
  nand (_21924_, _19692_, _19323_);
  nand (_21925_, _19324_, _09648_);
  nand (_21926_, _21925_, _21924_);
  nor (_21927_, _21926_, _19329_);
  nand (_21928_, _19329_, _19698_);
  nand (_21929_, _21928_, _19314_);
  nor (_21930_, _21929_, _21927_);
  nand (_21931_, _19704_, _19313_);
  nand (_21932_, _21931_, _19334_);
  nor (_21933_, _21932_, _21930_);
  nor (_21934_, _19709_, _19334_);
  nor (_09622_, _21934_, _21933_);
  nand (_21935_, _19324_, _09649_);
  nand (_21936_, _19714_, _19323_);
  nand (_21937_, _21936_, _21935_);
  nor (_21938_, _21937_, _19329_);
  nand (_21939_, _19329_, _19720_);
  nand (_21940_, _21939_, _19314_);
  nor (_21942_, _21940_, _21938_);
  nand (_21943_, _19727_, _19313_);
  nand (_21944_, _21943_, _19334_);
  nor (_21945_, _21944_, _21942_);
  nor (_21946_, _19732_, _19334_);
  nor (_09625_, _21946_, _21945_);
  nand (_21947_, _19324_, _09651_);
  nand (_21948_, _19735_, _19323_);
  nand (_21949_, _21948_, _21947_);
  nor (_21950_, _21949_, _19329_);
  nand (_21952_, _19329_, _19741_);
  nand (_21953_, _21952_, _19314_);
  nor (_21954_, _21953_, _21950_);
  nand (_21955_, _19747_, _19313_);
  nand (_21956_, _21955_, _19334_);
  nor (_21957_, _21956_, _21954_);
  nor (_21958_, _19752_, _19334_);
  nor (_09628_, _21958_, _21957_);
  nand (_21959_, _19297_, _09058_);
  nand (_21960_, _19608_, _19296_);
  nand (_21961_, _21960_, _21959_);
  nand (_21962_, _21961_, _19292_);
  not (_21963_, _19292_);
  nand (_21964_, _21963_, _08426_);
  nand (_21965_, _21964_, _21962_);
  nand (_21966_, _21965_, _19287_);
  nand (_21967_, _19286_, _08469_);
  nand (_21968_, _21967_, _21966_);
  nand (_21969_, _21968_, _19285_);
  nand (_21970_, _19284_, _08520_);
  nand (_09654_, _21970_, _21969_);
  nor (_21971_, _19287_, _08474_);
  nand (_21972_, _19297_, _08504_);
  nand (_21973_, _19628_, _19296_);
  nand (_21974_, _21973_, _21972_);
  nor (_21975_, _21974_, _21963_);
  nor (_21976_, _19292_, _08431_);
  nor (_21977_, _21976_, _21975_);
  nor (_21978_, _21977_, _19286_);
  nor (_21979_, _21978_, _21971_);
  nand (_21981_, _21979_, _19285_);
  nand (_21982_, _19284_, _08525_);
  nand (_09657_, _21982_, _21981_);
  nand (_21983_, _19286_, _08479_);
  nand (_21984_, _19297_, _09696_);
  nand (_21985_, _19650_, _19296_);
  nand (_21986_, _21985_, _21984_);
  nand (_21987_, _21986_, _19292_);
  nand (_21988_, _21963_, _08436_);
  nand (_21989_, _21988_, _21987_);
  nand (_21991_, _21989_, _19287_);
  nand (_21992_, _21991_, _21983_);
  nand (_21993_, _21992_, _19285_);
  nand (_21994_, _19284_, _08530_);
  nand (_09660_, _21994_, _21993_);
  nor (_21995_, _19287_, _08484_);
  nand (_21996_, _19297_, _09698_);
  nand (_21997_, _19670_, _19296_);
  nand (_21998_, _21997_, _21996_);
  nor (_21999_, _21998_, _21963_);
  nor (_22000_, _19292_, _08441_);
  nor (_22001_, _22000_, _21999_);
  nor (_22002_, _22001_, _19286_);
  nor (_22003_, _22002_, _21995_);
  nand (_22004_, _22003_, _19285_);
  nand (_22005_, _19284_, _08535_);
  nand (_09663_, _22005_, _22004_);
  nand (_22006_, _19297_, _09700_);
  nand (_22007_, _19692_, _19296_);
  nand (_22008_, _22007_, _22006_);
  nand (_22009_, _22008_, _19292_);
  nand (_22010_, _21963_, _08447_);
  nand (_22011_, _22010_, _22009_);
  nand (_22012_, _22011_, _19287_);
  nand (_22013_, _19286_, _08489_);
  nand (_22014_, _22013_, _22012_);
  nand (_22015_, _22014_, _19285_);
  nand (_22016_, _19284_, _08540_);
  nand (_09666_, _22016_, _22015_);
  nor (_22017_, _19287_, _08494_);
  nand (_22019_, _19297_, _09702_);
  nand (_22020_, _19714_, _19296_);
  nand (_22021_, _22020_, _22019_);
  nor (_22022_, _22021_, _21963_);
  nor (_22023_, _19292_, _08452_);
  nor (_22024_, _22023_, _22022_);
  nor (_22025_, _22024_, _19286_);
  nor (_22026_, _22025_, _22017_);
  nand (_22027_, _22026_, _19285_);
  nand (_22028_, _19284_, _08545_);
  nand (_09669_, _22028_, _22027_);
  nand (_22030_, _19286_, _08499_);
  nand (_22031_, _19297_, _09704_);
  nand (_22032_, _19735_, _19296_);
  nand (_22033_, _22032_, _22031_);
  nand (_22034_, _22033_, _19292_);
  nand (_22035_, _21963_, _08457_);
  nand (_22036_, _22035_, _22034_);
  nand (_22037_, _22036_, _19287_);
  nand (_22038_, _22037_, _22030_);
  nand (_22039_, _22038_, _19285_);
  nand (_22040_, _19284_, _08550_);
  nand (_09673_, _22040_, _22039_);
  nor (_22041_, _07863_, _05110_);
  nor (_22042_, _07690_, _18691_);
  nor (_22043_, _22042_, _18687_);
  not (_22044_, _22043_);
  nor (_22045_, _22044_, _22041_);
  nor (_22046_, _07708_, _05110_);
  nor (_22047_, _07835_, _18691_);
  nor (_22048_, _22047_, _05107_);
  not (_22049_, _22048_);
  nor (_22050_, _22049_, _22046_);
  nor (_22051_, _22050_, _22045_);
  nor (_22052_, _22051_, _18683_);
  nor (_22053_, _07726_, _18691_);
  nor (_22054_, _07780_, _05110_);
  nor (_22055_, _22054_, _22053_);
  not (_22056_, _22055_);
  nor (_22057_, _18687_, _05104_);
  not (_22059_, _22057_);
  nor (_22060_, _22059_, _22056_);
  nor (_22061_, _22060_, _05101_);
  nor (_22062_, _05107_, _05104_);
  nor (_22063_, _07658_, _05110_);
  nor (_22064_, _07638_, _18691_);
  nor (_22065_, _22064_, _22063_);
  nand (_22066_, _22065_, _22062_);
  nand (_22067_, _22066_, _22061_);
  nor (_22068_, _22067_, _22052_);
  nor (_22070_, _07902_, _18691_);
  nor (_22071_, _07915_, _05110_);
  nor (_22072_, _22071_, _22070_);
  nor (_22073_, _22072_, _18687_);
  nor (_22074_, _07546_, _18691_);
  nor (_22075_, _07743_, _05110_);
  nor (_22076_, _22075_, _22074_);
  nor (_22077_, _22076_, _05107_);
  nor (_22078_, _22077_, _22073_);
  not (_22079_, _22078_);
  nor (_22080_, _22079_, _18683_);
  nor (_22081_, _07679_, _05110_);
  nor (_22082_, _07731_, _18691_);
  nor (_22083_, _22082_, _22081_);
  nand (_22084_, _22083_, _22062_);
  nor (_22085_, _07880_, _18691_);
  nor (_22086_, _07817_, _05110_);
  nor (_22087_, _22086_, _22085_);
  nand (_22088_, _22087_, _22057_);
  nand (_22089_, _22088_, _22084_);
  nor (_22090_, _22089_, _22080_);
  nand (_22091_, _22090_, _05101_);
  not (_22092_, _22091_);
  nor (_22093_, _22092_, _22068_);
  not (_22094_, _22093_);
  nor (_22095_, _18683_, _05101_);
  not (_22096_, _22095_);
  nor (_22097_, _22096_, _21865_);
  nor (_22098_, _18683_, _18679_);
  not (_22099_, _22098_);
  nor (_22102_, _22099_, _21775_);
  nor (_22103_, _22102_, _22097_);
  not (_22104_, _22103_);
  nor (_22105_, _05104_, _18679_);
  nand (_22106_, _22105_, _09651_);
  nor (_22107_, _05104_, _05101_);
  nand (_22108_, _22107_, _09704_);
  nand (_22109_, _22108_, _22106_);
  nor (_22110_, _22109_, _22104_);
  nor (_22111_, _22110_, _05107_);
  nor (_22113_, _22096_, _20073_);
  nor (_22114_, _22099_, _20071_);
  nor (_22115_, _22114_, _22113_);
  not (_22116_, _22115_);
  nand (_22117_, _22105_, _09023_);
  nand (_22118_, _22107_, _09021_);
  nand (_22119_, _22118_, _22117_);
  nor (_22120_, _22119_, _22116_);
  nor (_22121_, _22120_, _18687_);
  nor (_22122_, _22121_, _22111_);
  nor (_22123_, _22122_, _05110_);
  nor (_22124_, _18691_, _05107_);
  nor (_22125_, _22099_, _21102_);
  not (_22126_, _22107_);
  nor (_22127_, _22126_, _21367_);
  nor (_22128_, _22127_, _22125_);
  nor (_22129_, _22096_, _21188_);
  not (_22130_, _22105_);
  nor (_22131_, _22130_, _21277_);
  nor (_22132_, _22131_, _22129_);
  nand (_22133_, _22132_, _22128_);
  nand (_22134_, _22133_, _22124_);
  not (_22135_, _22134_);
  nor (_22136_, _18691_, _18687_);
  not (_22137_, _22136_);
  nand (_22138_, _22098_, _08736_);
  nand (_22139_, _22095_, _08734_);
  nand (_22140_, _22139_, _22138_);
  nor (_22141_, _22126_, _21010_);
  not (_22142_, _22141_);
  nand (_22144_, _22105_, _08837_);
  nand (_22145_, _22144_, _22142_);
  nor (_22146_, _22145_, _22140_);
  nor (_22147_, _22146_, _22137_);
  nor (_22148_, _22147_, _22135_);
  not (_22149_, _22148_);
  nor (_22150_, _22149_, _22123_);
  nor (_22151_, _22150_, _22094_);
  nand (_22152_, _22095_, _08950_);
  nand (_22153_, _22098_, _08952_);
  nand (_22155_, _22153_, _22152_);
  nand (_22156_, _22105_, _09000_);
  nand (_22157_, _22107_, _08998_);
  nand (_22158_, _22157_, _22156_);
  nor (_22159_, _22158_, _22155_);
  nand (_22160_, _22159_, _05107_);
  nand (_22161_, _22098_, _09039_);
  not (_22162_, _22161_);
  nor (_22163_, _22096_, _21814_);
  nor (_22164_, _22163_, _22162_);
  not (_22165_, _22164_);
  nand (_22166_, _22107_, _09696_);
  nand (_22167_, _22105_, _09644_);
  nand (_22168_, _22167_, _22166_);
  nor (_22169_, _22168_, _22165_);
  nand (_22170_, _22169_, _18687_);
  nand (_22171_, _22170_, _22160_);
  nor (_22172_, _22171_, _05110_);
  nor (_22173_, _22099_, _21048_);
  nand (_22174_, _22107_, _08911_);
  not (_22175_, _22174_);
  nor (_22176_, _22175_, _22173_);
  nor (_22177_, _22096_, _21138_);
  nor (_22178_, _22130_, _21226_);
  nor (_22179_, _22178_, _22177_);
  nand (_22180_, _22179_, _22176_);
  nand (_22181_, _22180_, _22124_);
  nor (_22182_, _22099_, _19870_);
  nor (_22183_, _22126_, _19866_);
  nor (_22184_, _22183_, _22182_);
  nor (_22186_, _22096_, _19872_);
  nor (_22187_, _22130_, _19864_);
  nor (_22188_, _22187_, _22186_);
  nand (_22189_, _22188_, _22184_);
  nand (_22190_, _22189_, _22136_);
  nand (_22191_, _22190_, _22181_);
  nor (_22192_, _22191_, _22172_);
  nor (_22193_, _22192_, _22094_);
  not (_22194_, _22193_);
  nand (_22195_, _22095_, _08936_);
  nand (_22197_, _22098_, _08938_);
  nand (_22198_, _22197_, _22195_);
  nand (_22199_, _22105_, _08988_);
  nand (_22200_, _22107_, _08986_);
  nand (_22201_, _22200_, _22199_);
  nor (_22202_, _22201_, _22198_);
  nand (_22203_, _22202_, _05107_);
  nand (_22204_, _22105_, _09060_);
  not (_22205_, _22204_);
  nor (_22206_, _22205_, _05107_);
  nor (_22207_, _22096_, _21788_);
  nand (_22208_, _22098_, _08512_);
  nand (_22209_, _22107_, _09058_);
  nand (_22210_, _22209_, _22208_);
  nor (_22211_, _22210_, _22207_);
  nand (_22212_, _22211_, _22206_);
  nand (_22213_, _22212_, _22203_);
  nor (_22214_, _22213_, _05110_);
  nor (_22215_, _22099_, _21022_);
  nor (_22216_, _22126_, _21294_);
  nor (_22217_, _22216_, _22215_);
  nor (_22218_, _22096_, _21113_);
  nor (_22219_, _22130_, _21201_);
  nor (_22220_, _22219_, _22218_);
  nand (_22221_, _22220_, _22217_);
  nand (_22222_, _22221_, _22124_);
  nor (_22223_, _22099_, _19772_);
  nor (_22224_, _22126_, _19768_);
  nor (_22225_, _22224_, _22223_);
  nor (_22226_, _22096_, _19774_);
  nor (_22228_, _22130_, _19766_);
  nor (_22229_, _22228_, _22226_);
  nand (_22230_, _22229_, _22225_);
  nand (_22231_, _22230_, _22136_);
  nand (_22232_, _22231_, _22222_);
  nor (_22233_, _22232_, _22214_);
  nor (_22234_, _22233_, _22094_);
  nor (_22235_, _22234_, _22194_);
  nand (_22236_, _22095_, _08969_);
  nand (_22237_, _22098_, _08971_);
  nand (_22239_, _22237_, _22236_);
  nand (_22240_, _22105_, _09012_);
  nand (_22241_, _22107_, _09010_);
  nand (_22242_, _22241_, _22240_);
  nor (_22243_, _22242_, _22239_);
  nand (_22244_, _22243_, _05107_);
  nor (_22245_, _22099_, _21750_);
  nor (_22246_, _22096_, _21840_);
  nor (_22247_, _22246_, _22245_);
  not (_22248_, _22247_);
  nand (_22249_, _22107_, _09700_);
  nand (_22250_, _22105_, _09648_);
  nand (_22251_, _22250_, _22249_);
  nor (_22252_, _22251_, _22248_);
  nand (_22253_, _22252_, _18687_);
  nand (_22254_, _22253_, _22244_);
  nor (_22255_, _22254_, _05110_);
  nor (_22256_, _22099_, _21075_);
  nand (_22257_, _22107_, _08921_);
  not (_22258_, _22257_);
  nor (_22259_, _22258_, _22256_);
  nor (_22260_, _22096_, _21163_);
  nor (_22261_, _22130_, _21252_);
  nor (_22262_, _22261_, _22260_);
  nand (_22263_, _22262_, _22259_);
  nand (_22264_, _22263_, _22124_);
  not (_22265_, _22264_);
  nand (_22266_, _22098_, _08558_);
  nand (_22267_, _22095_, _08556_);
  nand (_22268_, _22267_, _22266_);
  nor (_22270_, _22126_, _20985_);
  not (_22271_, _22270_);
  nand (_22272_, _22105_, _08827_);
  nand (_22273_, _22272_, _22271_);
  nor (_22274_, _22273_, _22268_);
  nor (_22275_, _22274_, _22137_);
  nor (_22276_, _22275_, _22265_);
  not (_22277_, _22276_);
  nor (_22278_, _22277_, _22255_);
  nor (_22279_, _22278_, _22094_);
  nand (_22281_, _22095_, _08942_);
  nand (_22282_, _22098_, _08944_);
  nand (_22283_, _22282_, _22281_);
  nand (_22284_, _22105_, _08995_);
  nand (_22285_, _22107_, _08993_);
  nand (_22286_, _22285_, _22284_);
  nor (_22287_, _22286_, _22283_);
  nand (_22288_, _22287_, _05107_);
  nand (_22289_, _22105_, _08506_);
  not (_22290_, _22289_);
  nor (_22291_, _22290_, _05107_);
  nor (_22292_, _22096_, _21802_);
  nand (_22293_, _22098_, _09034_);
  nand (_22294_, _22107_, _08504_);
  nand (_22295_, _22294_, _22293_);
  nor (_22296_, _22295_, _22292_);
  nand (_22297_, _22296_, _22291_);
  nand (_22298_, _22297_, _22288_);
  nor (_22299_, _22298_, _05110_);
  nor (_22300_, _22099_, _21034_);
  nand (_22301_, _22107_, _08905_);
  not (_22302_, _22301_);
  nor (_22303_, _22302_, _22300_);
  nor (_22304_, _22096_, _21126_);
  nor (_22305_, _22130_, _21214_);
  nor (_22306_, _22305_, _22304_);
  nand (_22307_, _22306_, _22303_);
  nand (_22308_, _22307_, _22124_);
  not (_22309_, _22308_);
  nand (_22310_, _22098_, _08704_);
  nand (_22312_, _22095_, _08702_);
  nand (_22313_, _22312_, _22310_);
  nor (_22314_, _22126_, _20949_);
  not (_22315_, _22314_);
  nand (_22316_, _22105_, _08811_);
  nand (_22317_, _22316_, _22315_);
  nor (_22318_, _22317_, _22313_);
  nor (_22319_, _22318_, _22137_);
  nor (_22320_, _22319_, _22309_);
  not (_22321_, _22320_);
  nor (_22323_, _22321_, _22299_);
  nor (_22324_, _22323_, _22094_);
  not (_22325_, _22324_);
  not (_22326_, _22234_);
  nand (_22327_, _22326_, _22325_);
  nor (_22328_, _22327_, _22279_);
  nor (_22329_, _22328_, _22235_);
  nand (_22330_, _22095_, _08018_);
  nand (_22331_, _22098_, _08020_);
  nand (_22332_, _22331_, _22330_);
  nand (_22333_, _22105_, _08016_);
  nand (_22334_, _22107_, _08014_);
  nand (_22335_, _22334_, _22333_);
  nor (_22336_, _22335_, _22332_);
  nand (_22337_, _22336_, _05107_);
  nand (_22338_, _22098_, _08012_);
  not (_22339_, _22338_);
  nor (_22340_, _22096_, _19351_);
  nor (_22341_, _22340_, _22339_);
  not (_22342_, _08006_);
  nor (_22343_, _22126_, _22342_);
  nor (_22344_, _22130_, _19317_);
  nor (_22345_, _22344_, _22343_);
  nand (_22346_, _22345_, _22341_);
  nor (_22347_, _22346_, _05107_);
  nor (_22348_, _22347_, _05110_);
  nand (_22349_, _22348_, _22337_);
  not (_22350_, _22349_);
  nor (_22351_, _22099_, _19537_);
  nand (_22352_, _22107_, _08022_);
  not (_22354_, _22352_);
  nor (_22355_, _22354_, _22351_);
  nor (_22356_, _22096_, _19515_);
  nor (_22357_, _22130_, _19495_);
  nor (_22358_, _22357_, _22356_);
  nand (_22359_, _22358_, _22355_);
  nand (_22360_, _22359_, _22124_);
  nor (_22361_, _22099_, _18843_);
  nor (_22362_, _22126_, _18852_);
  nor (_22363_, _22362_, _22361_);
  nor (_22365_, _22096_, _18845_);
  nor (_22366_, _22130_, _18850_);
  nor (_22367_, _22366_, _22365_);
  nand (_22368_, _22367_, _22363_);
  nand (_22369_, _22368_, _22136_);
  nand (_22370_, _22369_, _22360_);
  nor (_22371_, _22370_, _22350_);
  nor (_22372_, _22371_, _22094_);
  not (_22373_, _22372_);
  nor (_22374_, _22096_, _20023_);
  nor (_22375_, _22099_, _20021_);
  nor (_22376_, _22375_, _22374_);
  not (_22377_, _22376_);
  nand (_22378_, _22105_, _09018_);
  nand (_22379_, _22107_, _09016_);
  nand (_22380_, _22379_, _22378_);
  nor (_22381_, _22380_, _22377_);
  nand (_22382_, _22381_, _05107_);
  nor (_22383_, _22096_, _21851_);
  nor (_22384_, _22099_, _21763_);
  nor (_22385_, _22384_, _22383_);
  not (_22386_, _22385_);
  nand (_22387_, _22105_, _09649_);
  nand (_22388_, _22107_, _09702_);
  nand (_22389_, _22388_, _22387_);
  nor (_22390_, _22389_, _22386_);
  nand (_22391_, _22390_, _18687_);
  nand (_22392_, _22391_, _22382_);
  nor (_22393_, _22392_, _05110_);
  nor (_22394_, _22099_, _21090_);
  nor (_22396_, _22126_, _21354_);
  nor (_22397_, _22396_, _22394_);
  nor (_22398_, _22096_, _21176_);
  nor (_22399_, _22130_, _21264_);
  nor (_22400_, _22399_, _22398_);
  nand (_22401_, _22400_, _22397_);
  nand (_22402_, _22401_, _22124_);
  not (_22403_, _22402_);
  nand (_22404_, _22098_, _08731_);
  nand (_22405_, _22107_, _08830_);
  nand (_22407_, _22405_, _22404_);
  nand (_22408_, _22095_, _08729_);
  nand (_22409_, _22105_, _08832_);
  nand (_22410_, _22409_, _22408_);
  nor (_22411_, _22410_, _22407_);
  nor (_22412_, _22411_, _22137_);
  nor (_22413_, _22412_, _22403_);
  not (_22414_, _22413_);
  nor (_22415_, _22414_, _22393_);
  nor (_22416_, _22415_, _22094_);
  not (_22417_, _22416_);
  nand (_22418_, _22417_, _22373_);
  nor (_22419_, _22418_, _22329_);
  not (_22420_, _22279_);
  nand (_22421_, _22095_, _08515_);
  nand (_22422_, _22098_, _08517_);
  nand (_22423_, _22422_, _22421_);
  nand (_22424_, _22105_, _09005_);
  nand (_22425_, _22107_, _09003_);
  nand (_22426_, _22425_, _22424_);
  nor (_22427_, _22426_, _22423_);
  nand (_22428_, _22427_, _05107_);
  nor (_22429_, _22096_, _21827_);
  nand (_22430_, _22098_, _09045_);
  not (_22431_, _22430_);
  nor (_22432_, _22431_, _22429_);
  nor (_22433_, _22130_, _21911_);
  nand (_22434_, _22107_, _09698_);
  not (_22435_, _22434_);
  nor (_22436_, _22435_, _22433_);
  nand (_22437_, _22436_, _22432_);
  nor (_22438_, _22437_, _05107_);
  nor (_22439_, _22438_, _05110_);
  nand (_22440_, _22439_, _22428_);
  nor (_22441_, _22099_, _21061_);
  nand (_22442_, _22107_, _08916_);
  not (_22443_, _22442_);
  nor (_22444_, _22443_, _22441_);
  nor (_22445_, _22096_, _21150_);
  nor (_22446_, _22130_, _21239_);
  nor (_22447_, _22446_, _22445_);
  nand (_22448_, _22447_, _22444_);
  nand (_22449_, _22448_, _22124_);
  not (_22450_, _22449_);
  nand (_22451_, _22098_, _08713_);
  nand (_22452_, _22107_, _08818_);
  nand (_22453_, _22452_, _22451_);
  nand (_22454_, _22095_, _08711_);
  nand (_22455_, _22105_, _08820_);
  nand (_22456_, _22455_, _22454_);
  nor (_22458_, _22456_, _22453_);
  nor (_22459_, _22458_, _22137_);
  nor (_22460_, _22459_, _22450_);
  nand (_22461_, _22460_, _22440_);
  nand (_22462_, _22461_, _22093_);
  not (_22463_, _22462_);
  nor (_22464_, _22324_, _22194_);
  not (_22465_, _22464_);
  nor (_22466_, _22465_, _22463_);
  nand (_22467_, _22466_, _22420_);
  nor (_22469_, _22417_, _22373_);
  nor (_22470_, _22234_, _22416_);
  nor (_22471_, _22470_, _22469_);
  nor (_22472_, _22471_, _22467_);
  not (_22473_, _22323_);
  nor (_22474_, _22326_, _22463_);
  nand (_22475_, _22474_, _22473_);
  nor (_22476_, _22475_, _22193_);
  nor (_22477_, _22476_, _22472_);
  nand (_22478_, _22279_, _22415_);
  nor (_22479_, _22478_, _22462_);
  nor (_22480_, _22325_, _22194_);
  nor (_22481_, _22480_, _22463_);
  nor (_22482_, _22481_, _22372_);
  nor (_22483_, _22482_, _22479_);
  nand (_22484_, _22483_, _22477_);
  nor (_22485_, _22484_, _22419_);
  nor (_22486_, _22485_, _22151_);
  nand (_22487_, _22235_, _22462_);
  nand (_22488_, _22487_, _22475_);
  nand (_22489_, _22488_, _22372_);
  not (_22490_, _22469_);
  nor (_22491_, _22474_, _22490_);
  not (_22492_, _22278_);
  nor (_22493_, _22492_, _22481_);
  nor (_22494_, _22493_, _22491_);
  nand (_22495_, _22494_, _22489_);
  nand (_22496_, _22495_, _22151_);
  nor (_22497_, _22418_, _22462_);
  nand (_22498_, _22417_, _22462_);
  nand (_22500_, _22279_, _22480_);
  nor (_22501_, _22500_, _22498_);
  nor (_22502_, _22501_, _22497_);
  nand (_22503_, _22502_, _22496_);
  nor (_22504_, _22503_, _22486_);
  nor (_22505_, _18699_, _18695_);
  nand (_22506_, _22505_, _05118_);
  nor (_22507_, _22506_, _18708_);
  not (_22508_, _22507_);
  nor (_22509_, _22137_, _18683_);
  not (_22511_, _22509_);
  nor (_22512_, _22511_, _22508_);
  not (_22513_, _22512_);
  nor (_22514_, _18717_, _18713_);
  not (_22515_, _22514_);
  nor (_22516_, _22515_, _18721_);
  not (_22517_, _22516_);
  nor (_22518_, _22517_, _18725_);
  not (_22519_, _22518_);
  nor (_22520_, _22519_, _22513_);
  not (_22522_, _22520_);
  nor (_22523_, _22522_, _18729_);
  not (_22524_, _22523_);
  nor (_22525_, _22524_, _18733_);
  not (_22526_, _22525_);
  nor (_22527_, _22526_, _18738_);
  nand (_22528_, _22527_, _05101_);
  not (_22529_, _22528_);
  nor (_22530_, _04471_, _04466_);
  nor (_22531_, _18609_, _18603_);
  nor (_22532_, _22531_, _22530_);
  nor (_22533_, _22526_, _18679_);
  nor (_22534_, _22533_, _05142_);
  nor (_22535_, _22534_, _05069_);
  nor (_22536_, _22535_, _22532_);
  nor (_22537_, _22536_, _22529_);
  nor (_22538_, _22532_, _22528_);
  nor (_22539_, _22137_, _22099_);
  not (_22540_, _22539_);
  nor (_22541_, _22540_, _22508_);
  not (_22543_, _22541_);
  nor (_22544_, _22543_, _22519_);
  not (_22545_, _22544_);
  nor (_22546_, _22545_, _18729_);
  nor (_22547_, _22546_, _18733_);
  not (_22548_, _22546_);
  nor (_22549_, _22548_, _05139_);
  nor (_22550_, _22549_, _22547_);
  not (_22551_, _22550_);
  nand (_22552_, _22551_, _18670_);
  nand (_22554_, _22550_, _05066_);
  nand (_22555_, _22554_, _22552_);
  nor (_22556_, _22555_, _22538_);
  nor (_22557_, _22534_, _22529_);
  nor (_22558_, _22557_, _18674_);
  nand (_22559_, _22545_, _18729_);
  nand (_22560_, _22559_, _22548_);
  nand (_22561_, _22560_, _05063_);
  nor (_22562_, _22560_, _05063_);
  nand (_22563_, _18721_, _18679_);
  nor (_22564_, _22515_, _22513_);
  nor (_22565_, _22564_, _05130_);
  nor (_22566_, _22543_, _22517_);
  nor (_22567_, _22566_, _22565_);
  nand (_22568_, _22567_, _22563_);
  nor (_22569_, _22568_, _05057_);
  nand (_22570_, _22568_, _05057_);
  nand (_22571_, _22509_, _22505_);
  nand (_22572_, _22571_, _18704_);
  nor (_22573_, _22540_, _22506_);
  nor (_22574_, _05118_, _05101_);
  nor (_22575_, _22574_, _22573_);
  nand (_22576_, _22575_, _22572_);
  nor (_22577_, _22576_, _05046_);
  nand (_22578_, _22576_, _05046_);
  nor (_22579_, _22571_, _18679_);
  nor (_22580_, _22540_, _18695_);
  nor (_22581_, _22580_, _05115_);
  nor (_22582_, _22581_, _22579_);
  not (_22583_, _22582_);
  nand (_22585_, _22583_, _05043_);
  nand (_22586_, _22585_, _22578_);
  nor (_22587_, _22586_, _22577_);
  nand (_22588_, _22587_, _22570_);
  nor (_22589_, _22588_, _22569_);
  not (_22590_, _22566_);
  nand (_22591_, _22590_, _18725_);
  nand (_22592_, _22566_, _05133_);
  nand (_22593_, _22592_, _22591_);
  nand (_22594_, _22593_, _05060_);
  nor (_22596_, _22543_, _18713_);
  not (_22597_, _22596_);
  nor (_22598_, _22597_, _05127_);
  nor (_22599_, _22596_, _18717_);
  nor (_22600_, _22599_, _22598_);
  not (_22601_, _22600_);
  nor (_22602_, _22601_, _05054_);
  nor (_22603_, _22600_, _18653_);
  nor (_22604_, _22603_, _22602_);
  nor (_22605_, _22541_, _05124_);
  nor (_22606_, _22605_, _22596_);
  not (_22607_, _22606_);
  nor (_22608_, _22607_, _05051_);
  nor (_22609_, _22608_, _22604_);
  nand (_22610_, _22609_, _22594_);
  not (_22611_, _22573_);
  nand (_22612_, _22611_, _18708_);
  nand (_22613_, _22612_, _22543_);
  nand (_22614_, _22613_, _05048_);
  nor (_22615_, _22099_, _18687_);
  nor (_22616_, _22615_, _05110_);
  nor (_22617_, _22616_, _22539_);
  nor (_22618_, _22617_, _05036_);
  not (_22619_, _22617_);
  nor (_22620_, _22619_, _18627_);
  nor (_22621_, _22620_, _22618_);
  nor (_22622_, _22613_, _05048_);
  nor (_22623_, _22622_, _22621_);
  nand (_22624_, _22623_, _22614_);
  nand (_22625_, _22582_, _18636_);
  nor (_22627_, _05107_, _18683_);
  not (_22628_, _22627_);
  nor (_22629_, _22628_, _18679_);
  nor (_22630_, _22098_, _18687_);
  nor (_22631_, _22630_, _22629_);
  nand (_22632_, _22631_, _05034_);
  not (_22633_, _22631_);
  nand (_22634_, _22633_, _18623_);
  nand (_22635_, _22634_, _22632_);
  nor (_22636_, _22095_, _22105_);
  not (_22638_, _22636_);
  nor (_22639_, _22638_, _18619_);
  nor (_22640_, _22636_, _05031_);
  nor (_22641_, _22640_, _22639_);
  nor (_22642_, _05112_, _05040_);
  nor (_22643_, _18695_, _18631_);
  nor (_22644_, _22643_, _22642_);
  not (_22645_, _22644_);
  nor (_22646_, _22645_, _22539_);
  nor (_22647_, _05101_, _18615_);
  nor (_22648_, _18679_, _05028_);
  nor (_22649_, _22648_, _22647_);
  not (_22650_, _22649_);
  nand (_22651_, _22645_, _22539_);
  nand (_22652_, _22651_, _22650_);
  nor (_22653_, _22652_, _22646_);
  nand (_22654_, _22653_, _22641_);
  nor (_22655_, _22654_, _22635_);
  nand (_22656_, _22655_, _22625_);
  nor (_22657_, _22656_, _22624_);
  nor (_22658_, _22593_, _05060_);
  nor (_22659_, _22606_, _18649_);
  nor (_22660_, _22659_, _22658_);
  nand (_22661_, _22660_, _22657_);
  nor (_22662_, _22661_, _22610_);
  nand (_22663_, _22662_, _22589_);
  nor (_22664_, _22663_, _22562_);
  nand (_22665_, _22664_, _22561_);
  nor (_22666_, _22665_, _22558_);
  nand (_22667_, _22666_, _22556_);
  nor (_22669_, _22667_, _22537_);
  nor (_22670_, _22669_, _22504_);
  nor (_22671_, _22420_, _22417_);
  not (_22672_, _22671_);
  nand (_22673_, _22672_, _22476_);
  nand (_22674_, _22474_, _22464_);
  nor (_22675_, _22674_, _22417_);
  nand (_22676_, _22675_, _22279_);
  nand (_22677_, _22676_, _22673_);
  not (_22678_, _22151_);
  not (_22680_, _22371_);
  nor (_22681_, _22680_, _22678_);
  nand (_22682_, _22681_, _22677_);
  nor (_22683_, _22234_, _22193_);
  nand (_22684_, _22683_, _22462_);
  nor (_22685_, _22684_, _22478_);
  nand (_22686_, _22685_, _22325_);
  nor (_22687_, _22674_, _22279_);
  nand (_22688_, _22687_, _22417_);
  nand (_22689_, _22688_, _22686_);
  not (_22690_, _22150_);
  nor (_22691_, _22373_, _22690_);
  nand (_22692_, _22691_, _22689_);
  nand (_22693_, _22692_, _22682_);
  nor (_22694_, _22137_, _22107_);
  not (_22695_, _22694_);
  nor (_22696_, _22695_, _22508_);
  not (_22697_, _22696_);
  nor (_22698_, _22697_, _22517_);
  not (_22699_, _22698_);
  nor (_22700_, _22699_, _18725_);
  nor (_22701_, _22698_, _05133_);
  nor (_22702_, _22701_, _22700_);
  nand (_22703_, _22702_, _18661_);
  not (_22704_, _22700_);
  nor (_22705_, _22704_, _18729_);
  not (_22706_, _22705_);
  nor (_22707_, _22706_, _18733_);
  nor (_22708_, _22705_, _05139_);
  nor (_22709_, _22708_, _22707_);
  nor (_22711_, _22709_, _18670_);
  nor (_22712_, _22695_, _22506_);
  nor (_22713_, _22695_, _18695_);
  not (_22714_, _22713_);
  nor (_22715_, _22714_, _18699_);
  nor (_22716_, _22715_, _05118_);
  nor (_22717_, _22716_, _22712_);
  not (_22718_, _22717_);
  nor (_22719_, _22718_, _05046_);
  nor (_22720_, _22719_, _22711_);
  nand (_22722_, _22720_, _22703_);
  nor (_22723_, _22107_, _18687_);
  nor (_22724_, _22723_, _05110_);
  nor (_22725_, _22724_, _22644_);
  not (_22726_, _22725_);
  nor (_22727_, _22644_, _05036_);
  nor (_22728_, _22727_, _22694_);
  nor (_22729_, _22728_, _05036_);
  nand (_22730_, _22729_, _22726_);
  nand (_22731_, _22728_, _22725_);
  nand (_22732_, _22731_, _22730_);
  nor (_22733_, _22697_, _22515_);
  nor (_22734_, _22733_, _05130_);
  nor (_22735_, _22734_, _22698_);
  nor (_22736_, _22735_, _18657_);
  not (_22737_, _22712_);
  nand (_22738_, _22737_, _05121_);
  nand (_22739_, _22712_, _18708_);
  nand (_22740_, _22739_, _22738_);
  nand (_22741_, _22740_, _18645_);
  nor (_22742_, _22697_, _18713_);
  nor (_22743_, _22742_, _05127_);
  nor (_22744_, _22743_, _22733_);
  not (_22745_, _22744_);
  nand (_22746_, _22745_, _05054_);
  nand (_22747_, _22746_, _22741_);
  nor (_22748_, _22747_, _22736_);
  nand (_22749_, _22748_, _22732_);
  nor (_22750_, _22749_, _22722_);
  nor (_22751_, _22697_, _22519_);
  not (_22753_, _22751_);
  nor (_22754_, _22753_, _18729_);
  nor (_22755_, _22751_, _05136_);
  nor (_22756_, _22755_, _22754_);
  not (_22757_, _22756_);
  nor (_22758_, _22757_, _18665_);
  nor (_22759_, _22756_, _05063_);
  nor (_22760_, _22759_, _22758_);
  not (_22761_, _22707_);
  nor (_22762_, _22761_, _18738_);
  nor (_22764_, _22762_, _04471_);
  not (_22765_, _22762_);
  nor (_22766_, _22765_, _18609_);
  nor (_22767_, _22766_, _22764_);
  nor (_22768_, _22767_, _18603_);
  nor (_22769_, _22768_, _22760_);
  not (_22770_, _22735_);
  nor (_22771_, _22770_, _05057_);
  not (_22772_, _22767_);
  nor (_22773_, _22772_, _04466_);
  nor (_22774_, _22773_, _22771_);
  nand (_22775_, _22774_, _22769_);
  not (_22776_, _22709_);
  nor (_22777_, _22776_, _05066_);
  nor (_22778_, _22707_, _05142_);
  nor (_22779_, _22778_, _22762_);
  not (_22780_, _22779_);
  nor (_22781_, _22780_, _18674_);
  nor (_22782_, _22779_, _05069_);
  nor (_22783_, _22782_, _22781_);
  nor (_22784_, _22783_, _22777_);
  not (_22785_, _22702_);
  nand (_22786_, _22785_, _05060_);
  nor (_22787_, _22696_, _05124_);
  nor (_22788_, _22787_, _22742_);
  nand (_22789_, _22788_, _05051_);
  not (_22790_, _22788_);
  nand (_22791_, _22790_, _18649_);
  nand (_22792_, _22791_, _22789_);
  nand (_22793_, _22792_, _22786_);
  nand (_22795_, _22744_, _18653_);
  nor (_22796_, _22740_, _18645_);
  nor (_22797_, _22714_, _05115_);
  nor (_22798_, _22713_, _18699_);
  nor (_22799_, _22798_, _22797_);
  nor (_22800_, _22799_, _05043_);
  nand (_22801_, _22799_, _05043_);
  not (_22802_, _22062_);
  nor (_22803_, _22105_, _22802_);
  nor (_22804_, _22803_, _22723_);
  nor (_22806_, _22804_, _18623_);
  nor (_22807_, _22806_, _22641_);
  nand (_22808_, _22807_, _22801_);
  nor (_22809_, _22808_, _22800_);
  nor (_22810_, _22717_, _18640_);
  nand (_22811_, _22804_, _18623_);
  nand (_22812_, _22811_, _22650_);
  nor (_22813_, _22812_, _22810_);
  nand (_22814_, _22813_, _22809_);
  nor (_22815_, _22814_, _22796_);
  nand (_22816_, _22815_, _22795_);
  nor (_22817_, _22816_, _22793_);
  nand (_22818_, _22817_, _22784_);
  nor (_22819_, _22818_, _22775_);
  nand (_22820_, _22819_, _22750_);
  nand (_22821_, _22820_, _22693_);
  nand (_22822_, _22466_, _22416_);
  nand (_22823_, _22822_, _22678_);
  nor (_22824_, _22687_, _22678_);
  nor (_22825_, _22480_, _22461_);
  nor (_22826_, _22825_, _22672_);
  nand (_22827_, _22466_, _22326_);
  nor (_22828_, _22684_, _22325_);
  not (_22829_, _22828_);
  nand (_22830_, _22829_, _22827_);
  nor (_22831_, _22830_, _22826_);
  nand (_22832_, _22831_, _22824_);
  nand (_22833_, _22832_, _22823_);
  nor (_22834_, _22674_, _22416_);
  nor (_22835_, _22834_, _22372_);
  nand (_22837_, _22835_, _22833_);
  not (_22838_, _22824_);
  not (_22839_, _22675_);
  not (_22840_, _22684_);
  nand (_22841_, _22840_, _22417_);
  nand (_22842_, _22841_, _22839_);
  nor (_22843_, _22842_, _22838_);
  nor (_22844_, _22684_, _22417_);
  not (_22845_, _22493_);
  not (_22846_, _22466_);
  nor (_22848_, _22478_, _22846_);
  nor (_22849_, _22848_, _22151_);
  nand (_22850_, _22849_, _22845_);
  nor (_22851_, _22850_, _22844_);
  nor (_22852_, _22851_, _22843_);
  nand (_22853_, _22828_, _22417_);
  nand (_22854_, _22853_, _22372_);
  nor (_22855_, _22854_, _22852_);
  nor (_22856_, _22525_, _05142_);
  nor (_22857_, _22856_, _05069_);
  nor (_22858_, _22857_, _22532_);
  nor (_22859_, _22858_, _22527_);
  nor (_22860_, _22524_, _05139_);
  nor (_22861_, _22523_, _18733_);
  nor (_22862_, _22861_, _22860_);
  nor (_22863_, _22862_, _05066_);
  nand (_22864_, _22862_, _05066_);
  not (_22865_, _22532_);
  nand (_22866_, _22865_, _22527_);
  nand (_22867_, _22866_, _22864_);
  nor (_22868_, _22867_, _22863_);
  nor (_22869_, _22856_, _22527_);
  nor (_22870_, _22869_, _18674_);
  nor (_22871_, _22520_, _05136_);
  nor (_22872_, _22871_, _22523_);
  nor (_22873_, _22872_, _18665_);
  not (_22874_, _22872_);
  nor (_22875_, _22874_, _05063_);
  nor (_22876_, _22875_, _22873_);
  nor (_22877_, _22513_, _18713_);
  nor (_22879_, _22512_, _05124_);
  nor (_22880_, _22879_, _22877_);
  nand (_22881_, _22880_, _05051_);
  not (_22882_, _22880_);
  nand (_22883_, _22882_, _18649_);
  nand (_22884_, _22883_, _22881_);
  nor (_22885_, _22571_, _18704_);
  not (_22886_, _22885_);
  nand (_22887_, _22572_, _22886_);
  nor (_22888_, _22887_, _18640_);
  not (_22890_, _22887_);
  nor (_22891_, _22890_, _05046_);
  nor (_22892_, _22891_, _22888_);
  nor (_22893_, _22877_, _05127_);
  nor (_22894_, _22893_, _22564_);
  nor (_22895_, _22894_, _18653_);
  nor (_22896_, _22895_, _22892_);
  nand (_22897_, _22896_, _22884_);
  nor (_22898_, _22517_, _22513_);
  nor (_22899_, _22565_, _22898_);
  not (_22900_, _22899_);
  nor (_22901_, _22900_, _05057_);
  nor (_22902_, _22899_, _18657_);
  nor (_22903_, _22902_, _22901_);
  not (_22904_, _22898_);
  nor (_22905_, _05133_, _18661_);
  nor (_22906_, _18725_, _05060_);
  nor (_22907_, _22906_, _22905_);
  not (_22908_, _22907_);
  nand (_22909_, _22908_, _22904_);
  nor (_22910_, _22511_, _18695_);
  nand (_22911_, _18699_, _18636_);
  nand (_22912_, _05115_, _05043_);
  nand (_22913_, _22912_, _22911_);
  nor (_22914_, _22913_, _22910_);
  nor (_22915_, _18687_, _18683_);
  not (_22916_, _22915_);
  nor (_22917_, _22916_, _05110_);
  nor (_22918_, _22915_, _18691_);
  nor (_22919_, _22918_, _22917_);
  not (_22921_, _22919_);
  nand (_22922_, _22921_, _18627_);
  nand (_22923_, _22913_, _22910_);
  nand (_22924_, _22923_, _22922_);
  nor (_22925_, _22924_, _22914_);
  nand (_22926_, _22628_, _22059_);
  nand (_22927_, _22926_, _18623_);
  nor (_22928_, _22926_, _18623_);
  nand (_22929_, _18683_, _05031_);
  nand (_22930_, _05104_, _18619_);
  nand (_22932_, _22930_, _22929_);
  nand (_22933_, _22649_, _22932_);
  nor (_22934_, _22933_, _22928_);
  nand (_22935_, _22934_, _22927_);
  nand (_22936_, _22645_, _22511_);
  nand (_22937_, _22644_, _22509_);
  nand (_22938_, _22937_, _22936_);
  nand (_22939_, _22919_, _05036_);
  nand (_22940_, _22939_, _22938_);
  nor (_22941_, _22940_, _22935_);
  nand (_22943_, _22941_, _22925_);
  nor (_22944_, _05121_, _05048_);
  nor (_22945_, _18708_, _18645_);
  nor (_22946_, _22945_, _22944_);
  nand (_22947_, _22946_, _22886_);
  not (_22948_, _22946_);
  nand (_22949_, _22948_, _22885_);
  nand (_22950_, _22949_, _22947_);
  nor (_22951_, _22950_, _22943_);
  nand (_22952_, _22951_, _22909_);
  nand (_22953_, _22907_, _22898_);
  nand (_22954_, _22894_, _18653_);
  nand (_22955_, _22954_, _22953_);
  nor (_22956_, _22955_, _22952_);
  nand (_22957_, _22956_, _22903_);
  nor (_22958_, _22957_, _22897_);
  nand (_22959_, _22958_, _22876_);
  nor (_22960_, _22959_, _22870_);
  nand (_22961_, _22960_, _22868_);
  nor (_22962_, _22961_, _22859_);
  nor (_22964_, _22962_, _22855_);
  nand (_22965_, _22964_, _22837_);
  nand (_22966_, _22965_, _22821_);
  nor (_22967_, _22966_, _22670_);
  nor (_22968_, _18623_, _18619_);
  not (_22969_, _22968_);
  nor (_22970_, _22969_, _18615_);
  nor (_22971_, _22970_, _05036_);
  not (_22972_, _22970_);
  nor (_22973_, _22972_, _18627_);
  nor (_22975_, _22973_, _22971_);
  nor (_22976_, _22975_, _07915_);
  nor (_22977_, _18619_, _18615_);
  nor (_22978_, _22977_, _05034_);
  nor (_22979_, _22978_, _22970_);
  nand (_22980_, _18920_, _05036_);
  nand (_22981_, _22980_, _22979_);
  nor (_22982_, _22981_, _22976_);
  nor (_22983_, _22975_, _07743_);
  not (_22984_, _22979_);
  nand (_22985_, _22975_, _18914_);
  nand (_22986_, _22985_, _22984_);
  nor (_22987_, _22986_, _22983_);
  nor (_22988_, _22987_, _22982_);
  nand (_22989_, _22988_, _05031_);
  nand (_22990_, _18765_, _18627_);
  nor (_22991_, _07679_, _18627_);
  nor (_22992_, _22991_, _22969_);
  nand (_22993_, _22992_, _22990_);
  nand (_22994_, _07817_, _18627_);
  not (_22995_, _22994_);
  nor (_22996_, _18948_, _18627_);
  nor (_22997_, _22996_, _22995_);
  not (_22998_, _22997_);
  nor (_22999_, _05034_, _18619_);
  nand (_23000_, _22999_, _22998_);
  nand (_23001_, _23000_, _22993_);
  nor (_23002_, _05031_, _05028_);
  nor (_23003_, _23002_, _18623_);
  nor (_23004_, _23003_, _05036_);
  not (_23006_, _23003_);
  nor (_23007_, _23006_, _18627_);
  nor (_23008_, _23007_, _23004_);
  nand (_23009_, _23008_, _07902_);
  nand (_23010_, _23002_, _18623_);
  nand (_23011_, _23010_, _23006_);
  nor (_23012_, _18918_, _05036_);
  nor (_23013_, _23012_, _23011_);
  nand (_23014_, _23013_, _23009_);
  nand (_23015_, _23014_, _18619_);
  not (_23017_, _23008_);
  nor (_23018_, _23017_, _07546_);
  nor (_23019_, _23008_, _07743_);
  nor (_23020_, _23019_, _23018_);
  not (_23021_, _23011_);
  nor (_23022_, _23021_, _23020_);
  nor (_23023_, _23022_, _23015_);
  nor (_23024_, _23023_, _23001_);
  nand (_23025_, _07638_, _05036_);
  nand (_23026_, _07658_, _18627_);
  nand (_23027_, _23026_, _23025_);
  nand (_23028_, _23027_, _18623_);
  nor (_23029_, _18931_, _05036_);
  not (_23030_, _23029_);
  nand (_23031_, _07726_, _05036_);
  nand (_23032_, _23031_, _23030_);
  nand (_23033_, _23032_, _05034_);
  nand (_23034_, _23033_, _23028_);
  nand (_23035_, _23034_, _18619_);
  nor (_23036_, _18902_, _18627_);
  nor (_23037_, _18899_, _05036_);
  nor (_23038_, _23037_, _18623_);
  not (_23039_, _23038_);
  nor (_23040_, _23039_, _23036_);
  nor (_23041_, _07708_, _05036_);
  nor (_23042_, _07835_, _18627_);
  nor (_23043_, _23042_, _23041_);
  nor (_23044_, _23043_, _05034_);
  nor (_23045_, _23044_, _23040_);
  nand (_23046_, _23045_, _05031_);
  nand (_23048_, _23046_, _23035_);
  nand (_23049_, _23048_, _18615_);
  nor (_23050_, _07638_, _05036_);
  nand (_23051_, _18800_, _05036_);
  nand (_23052_, _23051_, _22968_);
  nor (_23053_, _23052_, _23050_);
  nand (_23054_, _23032_, _22999_);
  nand (_23055_, _23045_, _18619_);
  nand (_23056_, _23055_, _23054_);
  nor (_23057_, _23056_, _23053_);
  nor (_23059_, _23057_, _23049_);
  nor (_23060_, _22975_, _07817_);
  nand (_23061_, _18948_, _05036_);
  nand (_23062_, _22979_, _23061_);
  nor (_23063_, _23062_, _23060_);
  nor (_23064_, _22975_, _07679_);
  nand (_23065_, _22975_, _18765_);
  nand (_23066_, _23065_, _22984_);
  nor (_23067_, _23066_, _23064_);
  nor (_23068_, _23067_, _23063_);
  nand (_23069_, _23068_, _18619_);
  nand (_23070_, _23069_, _23059_);
  nor (_23071_, _23070_, _23024_);
  nand (_23072_, _23071_, _22989_);
  nor (_23073_, _23008_, _18800_);
  nor (_23074_, _23017_, _18802_);
  nor (_23075_, _23074_, _23073_);
  nand (_23076_, _23075_, _23011_);
  nand (_23077_, _23008_, _07726_);
  nand (_23078_, _23077_, _23021_);
  nor (_23079_, _23078_, _23029_);
  nor (_23080_, _23079_, _05031_);
  nand (_23081_, _23080_, _23076_);
  nand (_23082_, _23008_, _07690_);
  nor (_23083_, _23037_, _23011_);
  nand (_23084_, _23083_, _23082_);
  nand (_23085_, _23017_, _07708_);
  nand (_23086_, _23008_, _07835_);
  nand (_23087_, _23086_, _23085_);
  nor (_23088_, _23087_, _23021_);
  nor (_23090_, _23088_, _18619_);
  nand (_23091_, _23090_, _23084_);
  nand (_23092_, _23091_, _23081_);
  nor (_23093_, _22975_, _07863_);
  nor (_23094_, _07690_, _18627_);
  nor (_23095_, _23094_, _23093_);
  nor (_23096_, _23095_, _22984_);
  not (_23097_, _22975_);
  nor (_23098_, _23097_, _07835_);
  nor (_23099_, _22975_, _07708_);
  nor (_23101_, _23099_, _23098_);
  nor (_23102_, _23101_, _22979_);
  nor (_23103_, _23102_, _23096_);
  nor (_23104_, _23103_, _05031_);
  nand (_23105_, _22975_, _18802_);
  nor (_23106_, _22975_, _07658_);
  nor (_23107_, _23106_, _22979_);
  nand (_23108_, _23107_, _23105_);
  nor (_23109_, _22975_, _07780_);
  nand (_23110_, _18933_, _05036_);
  nand (_23111_, _23110_, _22979_);
  nor (_23112_, _23111_, _23109_);
  nor (_23113_, _23112_, _18619_);
  nand (_23114_, _23113_, _23108_);
  not (_23115_, _22977_);
  nand (_23116_, _18918_, _18627_);
  nand (_23117_, _23116_, _22980_);
  nand (_23118_, _23117_, _05034_);
  nand (_23119_, _18910_, _18627_);
  nand (_23120_, _18914_, _05036_);
  nand (_23121_, _23120_, _23119_);
  nand (_23122_, _23121_, _18623_);
  nand (_23123_, _23122_, _23118_);
  nor (_23124_, _23123_, _23115_);
  nand (_23125_, _18619_, _05028_);
  nand (_23126_, _22997_, _05034_);
  nand (_23127_, _18761_, _18627_);
  nand (_23128_, _18765_, _05036_);
  nand (_23129_, _23128_, _23127_);
  nand (_23130_, _23129_, _18623_);
  nand (_23131_, _23130_, _23126_);
  nor (_23132_, _23131_, _23125_);
  nor (_23133_, _23132_, _23124_);
  nor (_23134_, _23123_, _05031_);
  nor (_23135_, _23134_, _23001_);
  nor (_23136_, _23135_, _23133_);
  nand (_23137_, _23136_, _23114_);
  nor (_23138_, _23137_, _23104_);
  nand (_23139_, _23138_, _23092_);
  nand (_23140_, _23139_, _23072_);
  nand (_23142_, _22617_, _07880_);
  nand (_23143_, _22619_, _07817_);
  nand (_23144_, _23143_, _23142_);
  nand (_23145_, _23144_, _22633_);
  nand (_23146_, _22617_, _07731_);
  nand (_23147_, _22619_, _07679_);
  nand (_23148_, _23147_, _23146_);
  nand (_23149_, _23148_, _22631_);
  nand (_23150_, _23149_, _23145_);
  nand (_23151_, _23150_, _22107_);
  nand (_23153_, _22619_, _07915_);
  nand (_23154_, _22617_, _07902_);
  nand (_23155_, _23154_, _23153_);
  nand (_23156_, _23155_, _22633_);
  nand (_23157_, _22617_, _07546_);
  nand (_23158_, _22619_, _07743_);
  nand (_23159_, _23158_, _23157_);
  nand (_23160_, _23159_, _22631_);
  nand (_23161_, _23160_, _23156_);
  nand (_23162_, _23161_, _22095_);
  nand (_23163_, _23162_, _23151_);
  nand (_23164_, _22617_, _07726_);
  nand (_23165_, _22619_, _07780_);
  nand (_23166_, _23165_, _23164_);
  nand (_23167_, _23166_, _22633_);
  nand (_23168_, _22617_, _18802_);
  nor (_23169_, _22617_, _07658_);
  nor (_23170_, _23169_, _22633_);
  nand (_23171_, _23170_, _23168_);
  nand (_23172_, _23171_, _23167_);
  nand (_23173_, _23172_, _22098_);
  nand (_23174_, _22619_, _07863_);
  nand (_23175_, _22617_, _07690_);
  nand (_23176_, _23175_, _23174_);
  nand (_23177_, _23176_, _22633_);
  nand (_23178_, _22617_, _07835_);
  nand (_23179_, _22619_, _07708_);
  nand (_23180_, _23179_, _23178_);
  nand (_23181_, _23180_, _22631_);
  nand (_23182_, _23181_, _23177_);
  nand (_23184_, _23182_, _22105_);
  nand (_23185_, _23184_, _23173_);
  nor (_23186_, _23185_, _23163_);
  nor (_23187_, _22724_, _22694_);
  not (_23188_, _23187_);
  nor (_23189_, _23188_, _18802_);
  nor (_23190_, _23187_, _18800_);
  nor (_23191_, _23190_, _23189_);
  nor (_23192_, _23191_, _22130_);
  nor (_23193_, _23192_, _22804_);
  nor (_23195_, _23188_, _18893_);
  nor (_23196_, _23187_, _18887_);
  nor (_23197_, _23196_, _23195_);
  nor (_23198_, _23197_, _22099_);
  nand (_23199_, _23187_, _07546_);
  nand (_23200_, _23188_, _07743_);
  nand (_23201_, _23200_, _23199_);
  nand (_23202_, _23201_, _22107_);
  nand (_23203_, _23187_, _07731_);
  nand (_23204_, _23188_, _07679_);
  nand (_23205_, _23204_, _23203_);
  nand (_23206_, _23205_, _22095_);
  nand (_23207_, _23206_, _23202_);
  nor (_23208_, _23207_, _23198_);
  nand (_23209_, _23208_, _23193_);
  nand (_23210_, _23188_, _18931_);
  nor (_23211_, _22130_, _22053_);
  nand (_23212_, _23211_, _23210_);
  nand (_23213_, _23212_, _22804_);
  nand (_23214_, _23187_, _18902_);
  nor (_23215_, _22099_, _22041_);
  nand (_23216_, _23215_, _23214_);
  nor (_23217_, _23187_, _07915_);
  not (_23218_, _22070_);
  nand (_23219_, _22107_, _23218_);
  nor (_23220_, _23219_, _23217_);
  nor (_23221_, _23187_, _07817_);
  not (_23222_, _22085_);
  nand (_23223_, _22095_, _23222_);
  nor (_23224_, _23223_, _23221_);
  nor (_23226_, _23224_, _23220_);
  nand (_23227_, _23226_, _23216_);
  nor (_23228_, _23227_, _23213_);
  not (_23229_, _22051_);
  nand (_23230_, _23229_, _18683_);
  not (_23231_, _22917_);
  nor (_23232_, _23231_, _18802_);
  nand (_23233_, _22627_, _22055_);
  nand (_23234_, _22509_, _07658_);
  nand (_23235_, _23234_, _23233_);
  nor (_23237_, _23235_, _23232_);
  nand (_23238_, _23237_, _23230_);
  nand (_23239_, _23238_, _18679_);
  nor (_23240_, _22130_, _22079_);
  nor (_23241_, _07679_, _18691_);
  nor (_23242_, _07731_, _05110_);
  nor (_23243_, _23242_, _23241_);
  nand (_23244_, _23243_, _22615_);
  nand (_23245_, _22629_, _22087_);
  nand (_23246_, _23245_, _23244_);
  nor (_23247_, _23246_, _23240_);
  nand (_23248_, _23247_, _23239_);
  not (_23249_, _10219_);
  nand (_23250_, _18604_, _23249_);
  nor (_23251_, _23250_, _22094_);
  nand (_23252_, _23251_, _23248_);
  nor (_23253_, _23252_, _23228_);
  nand (_23254_, _23253_, _23209_);
  nor (_23255_, _23254_, _23186_);
  nand (_23256_, _23255_, _23140_);
  nor (_10258_, _23256_, _22967_);
  nand (_23257_, _18601_, _10219_);
  nand (_10272_, _23257_, _29344_);
  nand (_25588_, _03362_, _03332_);
  not (_25590_, _25588_);
  not (_25592_, _03332_);
  nor (_25595_, _03783_, _03330_);
  not (_25597_, _25595_);
  nand (_25599_, _25597_, _25592_);
  not (_25601_, _25599_);
  not (_25603_, _04344_);
  nor (_25605_, _04342_, _04340_);
  nand (_25607_, _25605_, _25603_);
  nor (_25609_, _25597_, _03332_);
  not (_25611_, _25609_);
  nor (_25613_, _25611_, _25607_);
  not (_25615_, _04637_);
  not (_25617_, _05446_);
  nor (_25619_, _04414_, _04412_);
  nand (_25621_, _25619_, _04417_);
  nor (_25623_, _25621_, _25617_);
  not (_25625_, _05420_);
  nand (_25627_, _04414_, _04412_);
  nor (_25629_, _25627_, _04417_);
  not (_25631_, _25629_);
  nor (_25633_, _25631_, _25625_);
  nor (_25635_, _25633_, _25623_);
  not (_25637_, _05459_);
  not (_25639_, _04417_);
  nor (_25641_, _25619_, _25639_);
  not (_25643_, _25641_);
  nor (_25645_, _25643_, _25637_);
  not (_25647_, _25645_);
  nand (_25649_, _25647_, _25635_);
  not (_25651_, _05375_);
  not (_25653_, _04414_);
  nor (_25655_, _25653_, _04412_);
  nand (_25657_, _25655_, _25639_);
  nor (_25659_, _25657_, _25651_);
  not (_25661_, _05921_);
  nand (_25663_, _25619_, _25639_);
  nor (_25665_, _25663_, _25661_);
  nor (_25667_, _25665_, _25659_);
  not (_25669_, _05398_);
  not (_25671_, _04412_);
  nor (_25673_, _04414_, _25671_);
  nand (_25676_, _25673_, _25639_);
  nor (_25678_, _25676_, _25669_);
  not (_25680_, _30658_);
  not (_25682_, _04376_);
  nor (_25684_, _25682_, _25680_);
  nor (_25686_, _25684_, _25678_);
  nand (_25688_, _25686_, _25667_);
  nor (_25690_, _25688_, _25649_);
  nand (_25692_, _25690_, _25615_);
  nor (_25694_, _06047_, _25615_);
  nor (_25696_, _25694_, _00291_);
  nand (_25698_, _25696_, _25692_);
  nand (_25700_, _25698_, _25613_);
  nor (_25702_, _25609_, _03796_);
  nor (_25704_, _25702_, _25607_);
  nand (_25706_, _25704_, _25700_);
  not (_25708_, _25706_);
  not (_25710_, _25613_);
  not (_25712_, _25684_);
  not (_25714_, _06067_);
  nor (_25716_, _25643_, _25714_);
  not (_25718_, _06061_);
  nor (_25720_, _25657_, _25718_);
  nor (_25722_, _25720_, _25716_);
  nand (_25724_, _25629_, _04660_);
  not (_25726_, _25676_);
  nand (_25728_, _25726_, _06063_);
  nand (_25730_, _25728_, _25724_);
  not (_25732_, _06059_);
  nor (_25734_, _25663_, _25732_);
  not (_25736_, _06065_);
  nor (_25738_, _25621_, _25736_);
  nor (_25740_, _25738_, _25734_);
  not (_25742_, _25740_);
  nor (_25744_, _25742_, _25730_);
  nand (_25746_, _25744_, _25722_);
  nand (_25748_, _25746_, _25712_);
  nand (_25750_, _25748_, _25615_);
  nor (_25752_, _25615_, _04636_);
  nor (_25754_, _25752_, _00291_);
  nand (_25757_, _25754_, _25750_);
  not (_25759_, _25757_);
  nor (_25761_, _25759_, _25710_);
  nor (_25763_, _25609_, _03341_);
  nor (_25765_, _25763_, _25607_);
  not (_25767_, _25765_);
  nor (_25769_, _25767_, _25761_);
  not (_25771_, _04349_);
  nor (_25773_, _25643_, _25771_);
  not (_25775_, _25773_);
  not (_25777_, _05450_);
  nor (_25779_, _25621_, _25777_);
  not (_25781_, _05382_);
  nor (_25783_, _25657_, _25781_);
  nor (_25785_, _25783_, _25779_);
  nand (_25787_, _25629_, _05427_);
  not (_25789_, _25787_);
  not (_25791_, _05405_);
  nor (_25793_, _25676_, _25791_);
  nor (_25795_, _25793_, _25789_);
  nand (_25797_, _25795_, _25785_);
  not (_25799_, _05946_);
  nor (_25801_, _25663_, _25799_);
  nor (_25803_, _25801_, _25797_);
  nand (_25805_, _25803_, _25775_);
  nand (_25807_, _25805_, _25712_);
  nand (_25809_, _25807_, _25615_);
  nor (_25811_, _06051_, _25615_);
  nor (_25813_, _25811_, _00291_);
  nand (_25815_, _25813_, _25809_);
  not (_25817_, _25815_);
  nor (_25819_, _25817_, _25710_);
  nor (_25821_, _25609_, _03802_);
  nor (_25823_, _25821_, _25607_);
  not (_25825_, _25823_);
  nor (_25827_, _25825_, _25819_);
  nand (_25829_, _25641_, _05461_);
  not (_25831_, _05924_);
  nor (_25833_, _25663_, _25831_);
  not (_25835_, _05448_);
  nor (_25838_, _25621_, _25835_);
  nand (_25840_, _25629_, _05422_);
  not (_25842_, _25840_);
  nor (_25844_, _25842_, _25838_);
  not (_25846_, _05403_);
  nor (_25848_, _25676_, _25846_);
  not (_25850_, _05379_);
  nor (_25852_, _25657_, _25850_);
  nor (_25854_, _25852_, _25848_);
  nand (_25856_, _25854_, _25844_);
  nor (_25858_, _25856_, _25833_);
  nand (_25860_, _25858_, _25829_);
  nand (_25862_, _25860_, _25712_);
  nand (_25864_, _25862_, _25615_);
  nor (_25866_, _06049_, _25615_);
  nor (_25868_, _25866_, _00291_);
  nand (_25870_, _25868_, _25864_);
  not (_25872_, _25870_);
  nor (_25874_, _25872_, _25710_);
  nor (_25876_, _25609_, _03799_);
  nor (_25878_, _25876_, _25607_);
  not (_25880_, _25878_);
  nor (_25882_, _25880_, _25874_);
  not (_25884_, _25882_);
  nor (_25886_, _25884_, _25827_);
  nand (_25888_, _25886_, _25769_);
  nor (_25890_, _25888_, _25708_);
  not (_25892_, _25890_);
  nand (_25894_, _25641_, _05452_);
  not (_25896_, _05897_);
  nor (_25898_, _25663_, _25896_);
  not (_25900_, _05407_);
  nor (_25902_, _25631_, _25900_);
  not (_25904_, _05429_);
  nor (_25906_, _25621_, _25904_);
  nor (_25908_, _25906_, _25902_);
  not (_25910_, _05355_);
  nor (_25912_, _25657_, _25910_);
  not (_25914_, _05388_);
  nor (_25916_, _25676_, _25914_);
  nor (_25920_, _25916_, _25912_);
  nand (_25922_, _25920_, _25908_);
  nor (_25924_, _25922_, _25898_);
  nand (_25926_, _25924_, _25894_);
  nand (_25928_, _25926_, _25712_);
  nand (_25930_, _25928_, _25615_);
  nor (_25932_, _06040_, _25615_);
  nor (_25934_, _25932_, _00291_);
  nand (_25936_, _25934_, _25930_);
  not (_25938_, _25936_);
  nor (_25940_, _25938_, _25710_);
  nor (_25942_, _25609_, _03785_);
  nor (_25944_, _25942_, _25607_);
  not (_25946_, _25944_);
  nor (_25948_, _25946_, _25940_);
  not (_25950_, _25948_);
  not (_25952_, _00291_);
  not (_25954_, _05915_);
  nor (_25956_, _25663_, _25954_);
  not (_25958_, _05413_);
  nor (_25960_, _25631_, _25958_);
  nor (_25962_, _25960_, _25956_);
  not (_25964_, _25962_);
  not (_25966_, _05392_);
  nor (_25968_, _25676_, _25966_);
  not (_25970_, _05362_);
  nor (_25972_, _25657_, _25970_);
  nor (_25974_, _25972_, _25968_);
  nand (_25976_, _25641_, _05455_);
  not (_25978_, _25976_);
  not (_25980_, _05439_);
  nor (_25982_, _25621_, _25980_);
  nor (_25984_, _25982_, _25978_);
  nand (_25986_, _25984_, _25974_);
  nor (_25988_, _25986_, _25964_);
  nor (_25990_, _25988_, _25684_);
  nand (_25992_, _25990_, _25615_);
  nand (_25994_, _06043_, _04637_);
  nand (_25996_, _25994_, _25992_);
  nand (_25998_, _25996_, _25952_);
  not (_26001_, _25998_);
  nor (_26003_, _26001_, _25710_);
  nor (_26005_, _25609_, _03791_);
  nor (_26007_, _26005_, _25607_);
  not (_26009_, _26007_);
  nor (_26011_, _26009_, _26003_);
  not (_26013_, _05918_);
  nor (_26015_, _25663_, _26013_);
  not (_26017_, _05415_);
  nor (_26019_, _25631_, _26017_);
  nor (_26021_, _26019_, _26015_);
  not (_26023_, _26021_);
  not (_26025_, _05394_);
  nor (_26027_, _25676_, _26025_);
  not (_26029_, _05367_);
  nor (_26031_, _25657_, _26029_);
  nor (_26033_, _26031_, _26027_);
  nand (_26035_, _25641_, _05457_);
  not (_26037_, _26035_);
  not (_26039_, _05443_);
  nor (_26041_, _25621_, _26039_);
  nor (_26043_, _26041_, _26037_);
  nand (_26045_, _26043_, _26033_);
  nor (_26047_, _26045_, _26023_);
  nor (_26049_, _26047_, _25684_);
  nand (_26051_, _26049_, _25615_);
  nand (_26053_, _06045_, _04637_);
  nand (_26055_, _26053_, _26051_);
  nand (_26057_, _26055_, _25952_);
  not (_26059_, _26057_);
  nor (_26061_, _26059_, _25710_);
  nor (_26063_, _25609_, _03793_);
  nor (_26065_, _26063_, _25607_);
  not (_26067_, _26065_);
  nor (_26069_, _26067_, _26061_);
  nor (_26071_, _26069_, _26011_);
  not (_26073_, _05433_);
  nor (_26075_, _25621_, _26073_);
  not (_26077_, _05409_);
  nor (_26079_, _25631_, _26077_);
  nor (_26082_, _26079_, _26075_);
  not (_26084_, _05390_);
  nor (_26086_, _25676_, _26084_);
  not (_26088_, _26086_);
  nand (_26090_, _26088_, _26082_);
  not (_26092_, _05359_);
  nor (_26094_, _25657_, _26092_);
  nor (_26096_, _26094_, _25684_);
  not (_26098_, _05453_);
  nor (_26100_, _25643_, _26098_);
  not (_26102_, _05900_);
  nor (_26104_, _25663_, _26102_);
  nor (_26106_, _26104_, _26100_);
  nand (_26108_, _26106_, _26096_);
  nor (_26110_, _26108_, _26090_);
  nand (_26112_, _26110_, _25615_);
  nor (_26114_, _06042_, _25615_);
  nor (_26116_, _26114_, _00291_);
  nand (_26118_, _26116_, _26112_);
  nand (_26120_, _26118_, _25613_);
  nor (_26122_, _25609_, _03788_);
  nor (_26124_, _26122_, _25607_);
  nand (_26126_, _26124_, _26120_);
  not (_26128_, _26126_);
  nand (_26130_, _26128_, _26071_);
  nor (_26132_, _26130_, _25950_);
  not (_26134_, _26132_);
  nor (_26136_, _26134_, _25892_);
  not (_26138_, _25769_);
  not (_26140_, _25827_);
  nor (_26142_, _25884_, _26140_);
  nand (_26144_, _26142_, _26138_);
  nor (_26146_, _26144_, _25706_);
  nor (_26148_, _25827_, _26138_);
  nor (_26150_, _25882_, _25706_);
  nand (_26152_, _26150_, _26148_);
  not (_26154_, _26152_);
  nor (_26156_, _26154_, _26146_);
  nor (_26158_, _26156_, _26134_);
  nor (_26160_, _26158_, _26136_);
  nor (_26163_, _26160_, _25601_);
  not (_26165_, _03783_);
  not (_26167_, _03330_);
  nor (_26169_, _03332_, _26167_);
  nand (_26171_, _26169_, _26165_);
  not (_26173_, _26071_);
  nor (_26175_, _26128_, _25948_);
  not (_26177_, _26175_);
  nor (_26179_, _26177_, _26173_);
  not (_26181_, _26179_);
  nor (_26183_, _26181_, _26144_);
  nor (_26185_, _25882_, _26140_);
  nand (_26187_, _26185_, _26138_);
  nor (_26189_, _26187_, _26181_);
  nor (_26191_, _26189_, _26183_);
  nor (_26193_, _26191_, _26171_);
  nand (_26195_, _26148_, _25884_);
  nor (_26197_, _26195_, _25708_);
  not (_26199_, _26197_);
  not (_26201_, _26011_);
  nor (_26203_, _26069_, _26201_);
  nand (_26205_, _26203_, _26175_);
  nor (_26207_, _26205_, _26199_);
  nor (_26209_, _26205_, _25892_);
  nor (_26211_, _26209_, _26207_);
  not (_26213_, _26211_);
  nor (_26215_, _26213_, _26193_);
  not (_26217_, _26215_);
  nor (_26219_, _26217_, _26163_);
  nor (_26221_, _26219_, _03332_);
  nor (_26223_, _26221_, _25590_);
  not (_26225_, _26223_);
  nand (_26227_, _03819_, _03332_);
  not (_26229_, _26227_);
  nor (_26231_, _26130_, _25948_);
  nand (_26233_, _26231_, _26146_);
  not (_26235_, _26233_);
  nor (_26237_, _25892_, _26181_);
  nor (_26239_, _26237_, _26235_);
  not (_26241_, _26239_);
  not (_26244_, _26231_);
  nor (_26246_, _26187_, _25708_);
  not (_26248_, _26246_);
  nor (_26250_, _26248_, _26244_);
  nor (_26252_, _26134_, _26248_);
  nor (_26254_, _26252_, _26250_);
  not (_26256_, _26254_);
  nor (_26258_, _26256_, _26241_);
  nor (_26260_, _26199_, _26244_);
  nand (_26262_, _26140_, _25769_);
  nor (_26264_, _26262_, _25884_);
  nand (_26266_, _26264_, _25708_);
  nor (_26268_, _26266_, _26181_);
  nor (_26270_, _26268_, _26260_);
  nor (_26272_, _26187_, _25706_);
  not (_26274_, _26272_);
  nor (_26276_, _26274_, _26244_);
  nor (_26278_, _26274_, _26134_);
  nor (_26280_, _26278_, _26276_);
  nand (_26282_, _26280_, _26270_);
  nor (_26284_, _25827_, _25769_);
  nand (_26286_, _26284_, _25882_);
  nor (_26288_, _26286_, _25708_);
  nand (_26290_, _26288_, _26179_);
  nand (_26292_, _26284_, _25884_);
  nor (_26294_, _26292_, _25706_);
  nand (_26296_, _26294_, _26179_);
  not (_26298_, _26296_);
  nor (_26300_, _26286_, _25706_);
  not (_26302_, _26300_);
  nor (_26304_, _26302_, _26181_);
  nor (_26306_, _26304_, _26298_);
  nand (_26308_, _26306_, _26290_);
  nor (_26310_, _26308_, _26282_);
  nand (_26312_, _26310_, _26258_);
  nand (_26314_, _26128_, _26011_);
  nor (_26316_, _26314_, _26069_);
  nand (_26318_, _26316_, _25706_);
  nor (_26320_, _26318_, _25888_);
  not (_26322_, _26320_);
  nor (_26325_, _26128_, _25950_);
  nand (_26327_, _26325_, _26203_);
  not (_26329_, _26327_);
  nand (_26331_, _26142_, _25769_);
  nor (_26333_, _26331_, _25708_);
  nand (_26335_, _26333_, _26329_);
  nand (_26337_, _26335_, _26322_);
  nand (_26339_, _26154_, _26329_);
  nand (_26341_, _25890_, _26069_);
  nand (_26343_, _26341_, _26339_);
  nor (_26345_, _26343_, _26337_);
  nor (_26347_, _26144_, _25708_);
  nand (_26349_, _26347_, _26231_);
  nand (_26351_, _26347_, _26132_);
  nand (_26353_, _26351_, _26349_);
  nand (_26355_, _26264_, _26231_);
  nor (_26357_, _26355_, _25708_);
  nor (_26359_, _26357_, _26353_);
  nand (_26361_, _26359_, _26345_);
  nand (_26363_, _26329_, _26288_);
  nand (_26365_, _26154_, _26231_);
  nand (_26367_, _26365_, _26363_);
  nand (_26369_, _26347_, _26329_);
  nand (_26371_, _26329_, _26197_);
  nand (_26373_, _26371_, _26369_);
  nor (_26375_, _26373_, _26367_);
  nor (_26377_, _26140_, _26138_);
  nand (_26379_, _26377_, _25884_);
  nor (_26381_, _26379_, _25708_);
  nand (_26383_, _26381_, _26231_);
  nor (_26385_, _26327_, _25706_);
  nand (_26387_, _26385_, _26264_);
  nand (_26389_, _26387_, _26383_);
  nand (_26391_, _26381_, _26329_);
  nand (_26393_, _26329_, _26246_);
  nand (_26395_, _26393_, _26391_);
  nor (_26397_, _26395_, _26389_);
  nand (_26399_, _26397_, _26375_);
  nor (_26401_, _26399_, _26361_);
  nor (_26403_, _25882_, _25708_);
  nand (_26406_, _26284_, _26403_);
  nor (_26408_, _26406_, _26327_);
  not (_26410_, _26408_);
  nor (_26412_, _26355_, _25706_);
  not (_26414_, _26385_);
  not (_26416_, _26292_);
  not (_26418_, _26377_);
  nor (_26420_, _26418_, _25882_);
  nor (_26422_, _26420_, _26416_);
  nor (_26424_, _26422_, _26414_);
  nor (_26426_, _26424_, _26412_);
  nand (_26428_, _26426_, _26410_);
  not (_26430_, _26286_);
  nand (_26432_, _26430_, _26231_);
  nor (_26434_, _26379_, _25706_);
  nand (_26436_, _26434_, _26179_);
  nand (_26438_, _26436_, _26432_);
  not (_26440_, _26438_);
  nor (_26442_, _26300_, _26272_);
  nor (_26444_, _26442_, _26327_);
  nand (_26446_, _26381_, _26179_);
  nand (_26448_, _26434_, _26231_);
  nand (_26450_, _26448_, _26446_);
  nor (_26452_, _26450_, _26444_);
  nand (_26454_, _26452_, _26440_);
  nor (_26456_, _26454_, _26428_);
  nand (_26458_, _26456_, _26401_);
  nor (_26460_, _26458_, _26312_);
  nor (_26462_, _26460_, _25601_);
  nor (_26464_, _26165_, _03332_);
  not (_26466_, _26464_);
  nor (_26468_, _26466_, _26167_);
  not (_26470_, _26468_);
  nor (_26472_, _26470_, _26432_);
  nor (_26474_, _26472_, _26193_);
  not (_26476_, _26474_);
  nor (_26478_, _26476_, _26462_);
  nor (_26480_, _26478_, _03332_);
  nor (_26482_, _26480_, _26229_);
  nand (_26484_, _03817_, _03332_);
  not (_26487_, _26472_);
  not (_26489_, _26183_);
  nor (_26491_, _26489_, _26171_);
  not (_26493_, _26316_);
  nor (_26495_, _26493_, _26266_);
  not (_26497_, _26495_);
  nor (_26499_, _26379_, _26493_);
  nand (_26501_, _26316_, _26416_);
  not (_26503_, _26501_);
  nor (_26505_, _26503_, _26499_);
  nand (_26507_, _26505_, _26497_);
  nor (_26509_, _26318_, _26195_);
  not (_26511_, _26288_);
  nor (_26513_, _26493_, _26511_);
  nor (_26515_, _26513_, _26509_);
  not (_26517_, _26515_);
  nor (_26519_, _26517_, _26507_);
  nor (_26521_, _26318_, _26144_);
  nor (_26523_, _26152_, _26493_);
  nor (_26525_, _26523_, _26521_);
  not (_26527_, _26525_);
  nor (_26529_, _26527_, _26438_);
  nand (_26531_, _26529_, _26519_);
  not (_26533_, _26187_);
  nor (_26535_, _26333_, _26533_);
  nand (_26537_, _26535_, _26302_);
  nand (_26539_, _26537_, _26316_);
  nand (_26541_, _26539_, _26160_);
  nor (_26543_, _26541_, _26531_);
  nor (_26545_, _26543_, _25601_);
  nor (_26547_, _26545_, _26491_);
  nand (_26549_, _26547_, _26487_);
  nand (_26551_, _26549_, _25592_);
  nand (_26553_, _26551_, _26484_);
  nand (_26555_, _26553_, _26482_);
  nor (_26557_, _26555_, _26225_);
  not (_26559_, _26557_);
  not (_26561_, _30870_);
  not (_26563_, _30855_);
  not (_26565_, _30857_);
  nor (_26568_, _26565_, _26563_);
  nand (_26570_, _26568_, _30868_);
  nor (_26572_, _26570_, _26561_);
  nor (_26574_, _26572_, _30873_);
  not (_26576_, _03821_);
  not (_26578_, _03364_);
  not (_26580_, _03823_);
  nor (_26582_, _26580_, _03332_);
  nand (_26584_, _26582_, _26578_);
  nor (_26586_, _26584_, _26576_);
  nand (_26588_, _26572_, _30873_);
  nand (_26590_, _26588_, _26586_);
  nor (_26592_, _26590_, _26574_);
  not (_26594_, _03291_);
  nor (_26596_, _26576_, _03332_);
  not (_26598_, _26596_);
  nor (_26600_, _26598_, _03823_);
  nand (_26602_, _26600_, _03364_);
  nor (_26604_, _26602_, _26594_);
  nor (_26606_, _26604_, _26592_);
  nor (_26608_, _03821_, _03364_);
  nand (_26610_, _26608_, _26580_);
  nand (_26612_, _26610_, _25592_);
  nand (_26614_, _26612_, _05942_);
  not (_26616_, _26614_);
  not (_26618_, _03185_);
  nand (_26620_, _26600_, _26578_);
  nor (_26622_, _26620_, _26618_);
  nor (_26624_, _26622_, _26616_);
  not (_26626_, _26624_);
  nor (_26628_, _26598_, _26580_);
  nand (_26630_, _26628_, _03364_);
  nor (_26632_, _26584_, _03821_);
  nand (_26634_, _26632_, _05963_);
  nand (_26636_, _26634_, _26630_);
  nor (_26638_, _26636_, _26626_);
  nand (_26640_, _26638_, _26606_);
  not (_26642_, _26640_);
  not (_26644_, _30655_);
  not (_26646_, _30875_);
  nor (_26649_, _26588_, _26646_);
  nand (_26651_, _26588_, _26646_);
  nand (_26653_, _26651_, _26586_);
  nor (_26655_, _26653_, _26649_);
  not (_26657_, _26630_);
  not (_26659_, _03194_);
  nor (_26661_, _26620_, _26659_);
  nor (_26663_, _26661_, _26657_);
  nand (_26665_, _26632_, _05964_);
  not (_26667_, _26665_);
  not (_26669_, _03293_);
  nor (_26671_, _26602_, _26669_);
  nor (_26673_, _26671_, _26667_);
  nand (_26675_, _26673_, _26663_);
  nor (_26677_, _26675_, _26655_);
  not (_26679_, _26677_);
  nor (_26681_, _26679_, _26642_);
  not (_26683_, _26681_);
  nand (_26685_, _26649_, _30878_);
  not (_26687_, _26685_);
  nor (_26689_, _26687_, _30822_);
  not (_26691_, _26586_);
  not (_26693_, _30822_);
  nor (_26695_, _26685_, _26693_);
  nor (_26697_, _26695_, _26691_);
  not (_26699_, _26697_);
  nor (_26701_, _26699_, _26689_);
  not (_26703_, _03116_);
  nor (_26705_, _26620_, _26703_);
  nor (_26707_, _26705_, _26657_);
  nand (_26709_, _26632_, _06101_);
  not (_26711_, _26709_);
  not (_26713_, _03135_);
  nor (_26715_, _26602_, _26713_);
  nor (_26717_, _26715_, _26711_);
  nand (_26719_, _26717_, _26707_);
  nor (_26721_, _26719_, _26701_);
  nor (_26723_, _26649_, _30878_);
  nand (_26725_, _26685_, _26586_);
  nor (_26727_, _26725_, _26723_);
  not (_26731_, _03113_);
  nor (_26733_, _26620_, _26731_);
  nor (_26735_, _26733_, _26657_);
  nand (_26737_, _26632_, _05967_);
  not (_26739_, _26737_);
  not (_26741_, _03295_);
  nor (_26743_, _26602_, _26741_);
  nor (_26745_, _26743_, _26739_);
  nand (_26747_, _26745_, _26735_);
  nor (_26749_, _26747_, _26727_);
  nor (_26751_, _26749_, _26721_);
  not (_26753_, _03287_);
  nor (_26755_, _26602_, _26753_);
  not (_26757_, _03183_);
  nor (_26759_, _26620_, _26757_);
  nor (_26761_, _26759_, _26755_);
  nand (_26763_, _26570_, _26561_);
  nand (_26765_, _26763_, _26586_);
  nor (_26767_, _26765_, _26572_);
  nand (_26769_, _26612_, _05937_);
  nand (_26771_, _26632_, _05959_);
  nand (_26773_, _26771_, _26769_);
  nor (_26775_, _26773_, _26767_);
  nand (_26777_, _26775_, _26761_);
  not (_26779_, _26584_);
  nand (_26781_, _03366_, _25592_);
  nor (_26783_, _26781_, _30308_);
  not (_26785_, _26783_);
  nor (_26787_, _26785_, _26779_);
  not (_26789_, _26787_);
  nor (_26791_, _26789_, _26777_);
  not (_26793_, _26791_);
  not (_26795_, _26570_);
  nor (_26797_, _26568_, _30868_);
  nor (_26799_, _26797_, _26795_);
  nand (_26801_, _26799_, _26586_);
  nand (_26803_, _26632_, _05957_);
  nand (_26805_, _26803_, _26801_);
  not (_26807_, _26805_);
  not (_26809_, _03285_);
  nor (_26812_, _26602_, _26809_);
  not (_26814_, _03177_);
  nor (_26816_, _26620_, _26814_);
  not (_26818_, _26816_);
  nand (_26820_, _26612_, _05935_);
  nand (_26822_, _26820_, _26818_);
  nor (_26824_, _26822_, _26812_);
  nand (_26826_, _26824_, _26807_);
  nor (_26828_, _30857_, _30855_);
  nor (_26830_, _26828_, _26568_);
  nand (_26832_, _26830_, _26586_);
  nand (_26834_, _26632_, _05954_);
  nand (_26836_, _26834_, _26832_);
  not (_26838_, _03169_);
  nor (_26840_, _26620_, _26838_);
  not (_26842_, _26840_);
  not (_26844_, _03284_);
  nor (_26846_, _26602_, _26844_);
  nand (_26848_, _26612_, _05931_);
  not (_26850_, _26848_);
  nor (_26852_, _26850_, _26846_);
  nand (_26854_, _26852_, _26842_);
  nor (_26856_, _26854_, _26836_);
  not (_26858_, _26856_);
  not (_26860_, _03282_);
  nor (_26862_, _26602_, _26860_);
  not (_26864_, _03167_);
  nor (_26866_, _26620_, _26864_);
  nor (_26868_, _26866_, _26862_);
  not (_26870_, _26868_);
  nand (_26872_, _26632_, _05949_);
  nor (_26874_, _26691_, _30857_);
  nand (_26876_, _26612_, _05927_);
  not (_26878_, _26876_);
  nor (_26880_, _26878_, _26874_);
  nand (_26882_, _26880_, _26872_);
  nor (_26884_, _26882_, _26870_);
  not (_26886_, _26884_);
  nor (_26888_, _26886_, _26858_);
  not (_26890_, _26888_);
  nor (_26893_, _26890_, _26826_);
  not (_26895_, _26893_);
  nor (_26897_, _26895_, _26793_);
  nand (_26899_, _26897_, _26751_);
  nor (_26901_, _26899_, _26683_);
  nor (_26903_, _26901_, _26644_);
  not (_26905_, _03358_);
  nor (_26907_, _26905_, _03332_);
  not (_26909_, _26907_);
  nor (_26911_, _26909_, _03813_);
  not (_26913_, _26911_);
  not (_26915_, _03809_);
  nor (_26917_, _26915_, _03332_);
  not (_26919_, _26917_);
  nor (_26921_, _26919_, _03811_);
  not (_26923_, _26921_);
  nor (_26925_, _26923_, _26913_);
  not (_26927_, _26925_);
  not (_26929_, _03188_);
  not (_26931_, _03174_);
  nor (_26933_, _03181_, _26931_);
  nand (_26935_, _26933_, _03172_);
  nor (_26937_, _26935_, _26929_);
  not (_26939_, _03082_);
  nor (_26941_, _03181_, _03174_);
  nand (_26943_, _26941_, _03172_);
  nor (_26945_, _26943_, _26939_);
  nor (_26947_, _26945_, _26937_);
  not (_26949_, _03172_);
  nand (_26951_, _26933_, _26949_);
  nor (_26953_, _26951_, _26618_);
  nor (_26955_, _03174_, _03172_);
  nand (_26957_, _26955_, _03181_);
  nor (_26959_, _26957_, _26594_);
  nor (_26961_, _26959_, _26953_);
  nand (_26963_, _26961_, _26947_);
  not (_26965_, _26955_);
  nor (_26967_, _26965_, _03181_);
  not (_26969_, _04361_);
  nor (_26971_, _26969_, _04358_);
  nor (_26974_, _06135_, _23689_);
  not (_26976_, _06135_);
  nor (_26978_, _06172_, _26976_);
  nor (_26980_, _26978_, _26974_);
  nor (_26982_, _26980_, _26971_);
  not (_26984_, _04358_);
  nand (_26986_, _04361_, _26984_);
  nor (_26988_, _26986_, _06125_);
  nor (_26990_, _26988_, _26982_);
  nand (_26992_, _26990_, _26967_);
  nand (_26994_, _03181_, _03174_);
  nor (_26996_, _26994_, _26949_);
  nand (_26998_, _26996_, _03276_);
  not (_27000_, _03181_);
  nor (_27002_, _27000_, _26931_);
  nand (_27004_, _27002_, _26949_);
  not (_27006_, _27004_);
  nand (_27008_, _27006_, _01710_);
  nand (_27010_, _27008_, _26998_);
  not (_27012_, _27010_);
  nand (_27014_, _27012_, _26992_);
  nor (_27016_, _27014_, _26963_);
  not (_27018_, _27016_);
  nor (_27020_, _03090_, _03089_);
  nand (_27022_, _27020_, _26990_);
  nand (_27024_, _03090_, _03089_);
  nor (_27026_, _27024_, _26618_);
  not (_27028_, _27026_);
  not (_27030_, _03089_);
  nor (_27032_, _03090_, _27030_);
  nand (_27034_, _27032_, _01710_);
  nand (_27036_, _27034_, _27028_);
  not (_27038_, _27036_);
  nand (_27040_, _27038_, _27022_);
  nor (_27042_, _27040_, _27018_);
  nor (_27044_, _27042_, _26927_);
  not (_27046_, _03811_);
  nor (_27048_, _27046_, _03332_);
  nor (_27050_, _26917_, _27048_);
  not (_27052_, _27050_);
  nor (_27055_, _27052_, _26913_);
  not (_27057_, _27055_);
  not (_27059_, _23689_);
  nand (_27061_, _26976_, _27059_);
  not (_27063_, _06172_);
  nand (_27065_, _27063_, _06135_);
  nand (_27067_, _27065_, _27061_);
  nand (_27069_, _27067_, _26986_);
  not (_27071_, _06125_);
  nand (_27073_, _26971_, _27071_);
  nand (_27075_, _27073_, _27069_);
  not (_27077_, _27020_);
  nor (_27079_, _27077_, _27075_);
  nor (_27081_, _27036_, _27079_);
  nor (_27083_, _27081_, _27016_);
  nor (_27085_, _27083_, _27042_);
  not (_27087_, _27085_);
  nor (_27089_, _27087_, _27057_);
  nor (_27091_, _27089_, _27044_);
  not (_27093_, _27091_);
  not (_27095_, _30702_);
  not (_27097_, _03313_);
  nor (_27099_, _27097_, _27095_);
  nor (_27101_, _27099_, _03308_);
  not (_27103_, _06243_);
  not (_27105_, _23684_);
  nand (_27107_, _26976_, _27105_);
  not (_27109_, _06165_);
  nand (_27111_, _27109_, _06135_);
  nand (_27113_, _27111_, _27107_);
  nand (_27115_, _27113_, _27103_);
  nor (_27117_, _06269_, _06264_);
  not (_27119_, _27117_);
  nor (_27121_, _26980_, _27103_);
  nor (_27123_, _27121_, _27119_);
  nand (_27125_, _27123_, _27115_);
  nor (_27127_, _06135_, _23686_);
  nor (_27129_, _06167_, _26976_);
  nor (_27131_, _27129_, _27127_);
  nor (_27133_, _27131_, _06243_);
  not (_27136_, _06269_);
  nor (_27138_, _27136_, _06264_);
  not (_27140_, _23690_);
  nand (_27142_, _26976_, _27140_);
  not (_27144_, _06174_);
  nand (_27146_, _27144_, _06135_);
  nand (_27148_, _27146_, _27142_);
  nand (_27150_, _27148_, _06243_);
  nand (_27152_, _27150_, _27138_);
  nor (_27154_, _27152_, _27133_);
  nor (_27156_, _06135_, _23687_);
  nor (_27158_, _06169_, _26976_);
  nor (_27160_, _27158_, _27156_);
  nor (_27162_, _27160_, _06243_);
  not (_27164_, _06264_);
  nor (_27166_, _06269_, _27164_);
  nor (_27168_, _06135_, _23691_);
  not (_27170_, _27168_);
  not (_27172_, _06176_);
  nand (_27174_, _27172_, _06135_);
  nand (_27176_, _27174_, _27170_);
  nand (_27178_, _27176_, _06243_);
  nand (_27180_, _27178_, _27166_);
  nor (_27182_, _27180_, _27162_);
  nor (_27184_, _27182_, _27154_);
  nand (_27186_, _27184_, _27125_);
  nor (_27188_, _06135_, _04666_);
  not (_27190_, _27188_);
  not (_27192_, _06133_);
  nand (_27194_, _06135_, _27192_);
  nand (_27196_, _27194_, _27190_);
  nand (_27198_, _27196_, _06243_);
  nand (_27200_, _06269_, _06264_);
  nor (_27202_, _06135_, _23688_);
  nor (_27204_, _06170_, _26976_);
  nor (_27206_, _27204_, _27202_);
  nor (_27208_, _27206_, _06243_);
  nor (_27210_, _27208_, _27200_);
  nand (_27212_, _27210_, _27198_);
  nand (_27214_, _27212_, _26986_);
  nor (_27217_, _27214_, _27186_);
  nor (_27219_, _26986_, _04371_);
  nor (_27221_, _27219_, _27217_);
  nor (_27223_, _27221_, _03313_);
  nor (_27225_, _27223_, _27101_);
  not (_27227_, _03074_);
  nor (_27229_, _26943_, _27227_);
  not (_27231_, _03297_);
  nor (_27233_, _26935_, _27231_);
  nor (_27235_, _27233_, _27229_);
  nand (_27237_, _27006_, _01728_);
  not (_27239_, _27237_);
  nor (_27241_, _26957_, _26860_);
  nor (_27243_, _27241_, _27239_);
  nand (_27245_, _27243_, _27235_);
  nor (_27247_, _06135_, _23684_);
  nor (_27249_, _06165_, _26976_);
  nor (_27251_, _27249_, _27247_);
  nor (_27253_, _27251_, _26971_);
  nor (_27255_, _26986_, _06114_);
  nor (_27257_, _27255_, _27253_);
  nand (_27259_, _27257_, _26967_);
  nor (_27261_, _26951_, _26864_);
  nand (_27263_, _26996_, _03268_);
  not (_27265_, _27263_);
  nor (_27267_, _27265_, _27261_);
  nand (_27269_, _27267_, _27259_);
  nor (_27271_, _27269_, _27245_);
  nor (_27273_, _27131_, _26971_);
  nor (_27275_, _26986_, _06117_);
  nor (_27277_, _27275_, _27273_);
  nand (_27279_, _27277_, _26967_);
  not (_27281_, _03299_);
  nor (_27283_, _26935_, _27281_);
  not (_27285_, _27283_);
  nor (_27287_, _26957_, _26844_);
  not (_27289_, _27287_);
  nand (_27291_, _27289_, _27285_);
  not (_27293_, _03270_);
  not (_27295_, _26996_);
  nor (_27298_, _27295_, _27293_);
  not (_27300_, _01722_);
  nor (_27302_, _27004_, _27300_);
  nor (_27304_, _27302_, _27298_);
  not (_27306_, _03076_);
  nor (_27308_, _26943_, _27306_);
  nor (_27310_, _26951_, _26838_);
  nor (_27312_, _27310_, _27308_);
  nand (_27314_, _27312_, _27304_);
  nor (_27316_, _27314_, _27291_);
  nand (_27318_, _27316_, _27279_);
  nor (_27320_, _27160_, _26971_);
  nor (_27322_, _26986_, _06119_);
  nor (_27324_, _27322_, _27320_);
  nand (_27326_, _27324_, _26967_);
  nand (_27328_, _27000_, _03174_);
  nor (_27330_, _27328_, _26949_);
  nand (_27332_, _27330_, _03301_);
  nand (_27334_, _26996_, _03272_);
  nand (_27336_, _27334_, _27332_);
  nor (_27338_, _26957_, _26809_);
  not (_27340_, _01718_);
  nor (_27342_, _27004_, _27340_);
  nor (_27344_, _27342_, _27338_);
  not (_27346_, _03078_);
  nor (_27348_, _26943_, _27346_);
  nor (_27350_, _26951_, _26814_);
  nor (_27352_, _27350_, _27348_);
  nand (_27354_, _27352_, _27344_);
  nor (_27356_, _27354_, _27336_);
  nand (_27358_, _27356_, _27326_);
  nor (_27360_, _27358_, _27318_);
  nand (_27362_, _27360_, _27271_);
  not (_27364_, _03128_);
  nor (_27366_, _26935_, _27364_);
  not (_27368_, _03080_);
  nor (_27370_, _26943_, _27368_);
  nor (_27372_, _27370_, _27366_);
  nor (_27374_, _26957_, _26753_);
  nor (_27376_, _26951_, _26757_);
  nor (_27379_, _27376_, _27374_);
  nand (_27381_, _27379_, _27372_);
  nor (_27383_, _27206_, _26971_);
  nor (_27385_, _26986_, _06122_);
  nor (_27387_, _27385_, _27383_);
  nand (_27389_, _27387_, _26967_);
  not (_27391_, _01714_);
  nor (_27393_, _27004_, _27391_);
  not (_27395_, _03274_);
  nor (_27397_, _27295_, _27395_);
  nor (_27399_, _27397_, _27393_);
  nand (_27401_, _27399_, _27389_);
  nor (_27403_, _27401_, _27381_);
  not (_27405_, _27403_);
  nor (_27407_, _27405_, _27362_);
  nand (_27409_, _27407_, _27225_);
  not (_27411_, _27101_);
  nor (_27413_, _06176_, _26976_);
  nor (_27415_, _27413_, _27168_);
  nand (_27417_, _27415_, _06243_);
  nand (_27419_, _27160_, _27103_);
  nand (_27421_, _27419_, _27417_);
  nand (_27423_, _27421_, _27166_);
  nor (_27425_, _27200_, _06243_);
  nand (_27427_, _27425_, _27206_);
  nor (_27429_, _27119_, _27103_);
  nand (_27431_, _27429_, _26980_);
  nand (_27433_, _27431_, _27427_);
  nor (_27435_, _27119_, _06243_);
  nand (_27437_, _27435_, _27251_);
  nor (_27439_, _26976_, _06133_);
  nor (_27441_, _27439_, _27188_);
  nor (_27443_, _27200_, _27103_);
  nand (_27445_, _27443_, _27441_);
  nand (_27447_, _27445_, _27437_);
  nor (_27449_, _27447_, _27433_);
  nand (_27451_, _27449_, _27423_);
  nor (_27453_, _27451_, _27154_);
  nor (_27455_, _27453_, _26971_);
  not (_27457_, _04371_);
  nor (_27460_, _26986_, _27457_);
  nor (_27462_, _27460_, _27455_);
  nand (_27464_, _27462_, _27097_);
  nand (_27466_, _27464_, _27411_);
  nor (_27468_, _27308_, _27283_);
  nor (_27470_, _27310_, _27287_);
  nand (_27472_, _27470_, _27468_);
  nand (_27474_, _27304_, _27279_);
  nor (_27476_, _27474_, _27472_);
  nor (_27478_, _27476_, _27271_);
  nand (_27480_, _27478_, _27358_);
  nor (_27482_, _27480_, _27403_);
  nand (_27484_, _27482_, _27466_);
  nand (_27486_, _27484_, _27409_);
  nand (_27488_, _27486_, _27018_);
  not (_27490_, _27048_);
  nor (_27492_, _27490_, _03809_);
  not (_27494_, _27492_);
  not (_27496_, _03813_);
  nor (_27498_, _27496_, _03332_);
  not (_27500_, _27498_);
  nor (_27502_, _27500_, _26905_);
  not (_27504_, _27502_);
  nor (_27506_, _27504_, _27494_);
  not (_27508_, _27506_);
  nor (_27510_, _27486_, _27018_);
  nor (_27512_, _27510_, _27508_);
  nand (_27514_, _27512_, _27488_);
  nor (_27516_, _27040_, _27466_);
  not (_27518_, _27516_);
  nor (_27520_, _27490_, _26915_);
  not (_27522_, _27520_);
  nor (_27524_, _27522_, _27504_);
  not (_27526_, _27524_);
  nor (_27528_, _27018_, _27225_);
  nor (_27530_, _27528_, _27526_);
  nand (_27532_, _27530_, _27518_);
  nand (_27534_, _27532_, _27514_);
  nor (_27536_, _27534_, _27093_);
  not (_27538_, _27536_);
  nor (_27542_, _27500_, _03358_);
  not (_27544_, _27542_);
  nor (_27546_, _27544_, _27522_);
  not (_27548_, _27546_);
  not (_27550_, _27083_);
  nor (_27552_, _27550_, _27548_);
  not (_27554_, _27552_);
  nor (_27556_, _26913_, _03811_);
  not (_27558_, _27556_);
  nor (_27560_, _26907_, _27498_);
  not (_27562_, _27560_);
  nor (_27564_, _27562_, _27494_);
  nor (_27566_, _27500_, _27046_);
  nor (_27568_, _27566_, _27564_);
  nand (_27570_, _27568_, _27558_);
  nor (_27572_, _27570_, _27016_);
  nor (_27574_, _27544_, _27494_);
  not (_27576_, _27574_);
  nor (_27578_, _27576_, _27018_);
  nor (_27580_, _27578_, _27572_);
  nand (_27582_, _27580_, _27554_);
  nor (_27584_, _27582_, _27538_);
  not (_27586_, _26901_);
  nor (_27588_, _27586_, _27584_);
  nor (_27590_, _27588_, _26903_);
  not (_27592_, _27590_);
  nor (_27594_, _27592_, _26642_);
  nor (_27596_, _27590_, _26640_);
  nor (_27598_, _27596_, _27594_);
  not (_27600_, _27598_);
  nor (_27602_, _26886_, _25950_);
  nor (_27604_, _26884_, _25948_);
  nor (_27606_, _27604_, _27602_);
  not (_27608_, _26721_);
  not (_27610_, _26749_);
  nor (_27612_, _27610_, _27608_);
  not (_27614_, _27612_);
  nor (_27616_, _26826_, _26858_);
  nand (_27618_, _27616_, _26783_);
  nor (_27620_, _27618_, _27614_);
  nand (_27623_, _27620_, _27606_);
  nor (_27625_, _27623_, _26679_);
  not (_27627_, _30691_);
  nor (_27629_, _26901_, _27627_);
  nor (_27631_, _27570_, _27403_);
  nand (_27633_, _27020_, _27387_);
  nor (_27635_, _27024_, _26757_);
  not (_27637_, _27635_);
  nand (_27639_, _27032_, _01714_);
  nand (_27641_, _27639_, _27637_);
  not (_27643_, _27641_);
  nand (_27645_, _27643_, _27633_);
  nor (_27647_, _27645_, _27405_);
  nor (_27649_, _27647_, _26927_);
  not (_27651_, _23688_);
  nand (_27653_, _26976_, _27651_);
  not (_27655_, _06170_);
  nand (_27657_, _27655_, _06135_);
  nand (_27659_, _27657_, _27653_);
  nand (_27661_, _27659_, _26986_);
  not (_27663_, _06122_);
  nand (_27665_, _26971_, _27663_);
  nand (_27667_, _27665_, _27661_);
  nor (_27669_, _27077_, _27667_);
  nor (_27671_, _27641_, _27669_);
  nor (_27673_, _27671_, _27403_);
  nor (_27675_, _27673_, _27647_);
  not (_27677_, _27675_);
  nor (_27679_, _27677_, _27057_);
  nor (_27681_, _27679_, _27649_);
  not (_27683_, _27681_);
  nand (_27685_, _27362_, _27225_);
  nand (_27687_, _27480_, _27466_);
  nand (_27689_, _27687_, _27685_);
  nand (_27691_, _27689_, _27403_);
  nor (_27693_, _27689_, _27403_);
  nor (_27695_, _27693_, _27508_);
  nand (_27697_, _27695_, _27691_);
  nor (_27699_, _27671_, _27526_);
  not (_27701_, _27699_);
  nand (_27704_, _27701_, _27697_);
  nor (_27706_, _27704_, _27683_);
  nor (_27708_, _27576_, _27405_);
  not (_27710_, _27673_);
  nor (_27712_, _27710_, _27548_);
  nor (_27714_, _27712_, _27708_);
  nand (_27716_, _27714_, _27706_);
  nor (_27718_, _27716_, _27631_);
  nor (_27720_, _27586_, _27718_);
  nor (_27722_, _27720_, _27629_);
  nor (_27724_, _27722_, _26777_);
  not (_27726_, _26777_);
  not (_27728_, _27629_);
  nand (_27730_, _27691_, _27506_);
  nor (_27732_, _27730_, _27693_);
  nor (_27734_, _27699_, _27732_);
  nand (_27736_, _27734_, _27681_);
  nor (_27738_, _27736_, _27708_);
  nor (_27740_, _27712_, _27631_);
  nand (_27742_, _27740_, _27738_);
  nand (_27744_, _26901_, _27742_);
  nand (_27746_, _27744_, _27728_);
  nor (_27748_, _27746_, _27726_);
  nor (_27750_, _27748_, _27724_);
  nand (_27752_, _27750_, _27625_);
  nor (_27754_, _27752_, _27600_);
  not (_27756_, _06438_);
  nor (_27758_, _27722_, _25948_);
  nand (_27760_, _27758_, _27592_);
  nor (_27762_, _27760_, _27756_);
  not (_27764_, _06482_);
  nor (_27766_, _27722_, _25950_);
  nand (_27768_, _27766_, _27592_);
  nor (_27770_, _27768_, _27764_);
  nor (_27772_, _27770_, _27762_);
  not (_27774_, _06610_);
  nor (_27776_, _27746_, _25950_);
  nand (_27778_, _27776_, _27592_);
  nor (_27780_, _27778_, _27774_);
  not (_27782_, _06567_);
  nand (_27785_, _27766_, _27590_);
  nor (_27787_, _27785_, _27782_);
  nor (_27789_, _27787_, _27780_);
  nand (_27791_, _27789_, _27772_);
  not (_27793_, _06525_);
  nand (_27795_, _27776_, _27590_);
  nor (_27797_, _27795_, _27793_);
  not (_27799_, _06503_);
  nor (_27801_, _27746_, _25948_);
  nand (_27803_, _27801_, _27590_);
  nor (_27805_, _27803_, _27799_);
  nor (_27807_, _27805_, _27797_);
  not (_27809_, _06546_);
  nand (_27811_, _27758_, _27590_);
  nor (_27813_, _27811_, _27809_);
  not (_27815_, _06589_);
  nand (_27817_, _27801_, _27592_);
  nor (_27819_, _27817_, _27815_);
  nor (_27821_, _27819_, _27813_);
  nand (_27823_, _27821_, _27807_);
  nor (_27825_, _27823_, _27791_);
  nor (_27827_, _27825_, _27754_);
  nor (_27829_, _27570_, _27271_);
  nand (_27831_, _27113_, _26986_);
  not (_27833_, _06114_);
  nand (_27835_, _26971_, _27833_);
  nand (_27837_, _27835_, _27831_);
  nor (_27839_, _27077_, _27837_);
  nor (_27841_, _27024_, _26864_);
  not (_27843_, _27841_);
  nand (_27845_, _27032_, _01728_);
  nand (_27847_, _27845_, _27843_);
  nor (_27849_, _27847_, _27839_);
  nor (_27851_, _27849_, _27271_);
  not (_27853_, _27851_);
  nor (_27855_, _27853_, _27548_);
  nor (_27857_, _27855_, _27829_);
  nor (_27859_, _27849_, _27526_);
  not (_27861_, _27271_);
  nor (_27863_, _27508_, _27861_);
  nor (_27866_, _27863_, _27859_);
  nand (_27868_, _27849_, _27271_);
  nand (_27870_, _27868_, _27853_);
  nor (_27872_, _27870_, _27057_);
  not (_27874_, _27868_);
  nor (_27876_, _27874_, _26927_);
  nor (_27878_, _27876_, _27872_);
  nand (_27880_, _27878_, _27866_);
  nor (_27882_, _27576_, _27861_);
  nor (_27884_, _27882_, _27880_);
  nand (_27886_, _27884_, _27857_);
  not (_27888_, _27886_);
  not (_27890_, _27754_);
  nor (_27892_, _27890_, _27888_);
  nor (_27894_, _27892_, _27827_);
  nor (_27896_, _27894_, _26559_);
  not (_27898_, _27896_);
  nor (_27900_, _26553_, _26482_);
  nand (_27902_, _27900_, _26223_);
  nor (_27904_, _25609_, _26864_);
  nor (_27906_, _25684_, _25611_);
  not (_27908_, _27906_);
  not (_27910_, _05464_);
  nor (_27912_, _25643_, _27910_);
  not (_27914_, _05452_);
  nor (_27916_, _25621_, _27914_);
  nor (_27918_, _27916_, _27912_);
  not (_27920_, _27918_);
  nor (_27922_, _25663_, _25910_);
  nor (_27924_, _25676_, _25900_);
  nor (_27926_, _27924_, _27922_);
  nor (_27928_, _25631_, _25904_);
  nor (_27930_, _25657_, _25914_);
  nor (_27932_, _27930_, _27928_);
  nand (_27934_, _27932_, _27926_);
  nor (_27936_, _27934_, _27920_);
  nor (_27938_, _27936_, _27908_);
  nor (_27940_, _27938_, _27904_);
  nor (_27942_, _27940_, _27902_);
  nand (_27944_, _26553_, _26223_);
  nor (_27947_, _27944_, _26482_);
  nor (_27949_, _26781_, _26779_);
  nor (_27951_, _26679_, _26640_);
  nor (_27953_, _27610_, _26721_);
  nand (_27955_, _27953_, _27951_);
  nor (_27957_, _26884_, _26858_);
  not (_27959_, _27957_);
  nor (_27961_, _26826_, _27959_);
  nand (_27963_, _27961_, _27726_);
  nor (_27965_, _27963_, _27955_);
  nand (_27967_, _27965_, _27949_);
  nor (_27969_, _27967_, _30308_);
  nand (_27971_, _27886_, _27969_);
  not (_27973_, _27971_);
  not (_27975_, _30951_);
  not (_27977_, _27955_);
  nor (_27979_, _26793_, _26826_);
  not (_27981_, _27979_);
  nor (_27983_, _27981_, _27959_);
  nand (_27985_, _27983_, _27977_);
  not (_27987_, _27985_);
  nor (_27989_, _27987_, _26565_);
  not (_27991_, _27989_);
  nand (_27993_, _27971_, _27991_);
  nor (_27995_, _27993_, _27975_);
  nor (_27997_, _27973_, _27989_);
  nor (_27999_, _27997_, _30951_);
  nor (_28001_, _27999_, _27995_);
  nor (_28003_, _28001_, _26586_);
  nor (_28005_, _28003_, _26874_);
  nor (_28007_, _28005_, _27969_);
  nor (_28009_, _28007_, _27973_);
  not (_28011_, _28009_);
  nand (_28013_, _28011_, _27947_);
  nor (_28015_, _26553_, _26225_);
  nand (_28017_, _28015_, _26482_);
  not (_28019_, _28017_);
  nand (_28021_, _28019_, _25948_);
  nand (_28023_, _28021_, _28013_);
  nor (_28025_, _28023_, _27942_);
  nand (_28028_, _28025_, _27898_);
  nor (_28030_, _25609_, _26838_);
  not (_28032_, _05468_);
  nor (_28034_, _25643_, _28032_);
  nor (_28036_, _25621_, _26098_);
  nor (_28038_, _28036_, _28034_);
  not (_28040_, _28038_);
  nor (_28042_, _25657_, _26084_);
  nor (_28044_, _25676_, _26077_);
  nor (_28046_, _28044_, _28042_);
  nor (_28048_, _25663_, _26092_);
  nor (_28050_, _25631_, _26073_);
  nor (_28052_, _28050_, _28048_);
  nand (_28054_, _28052_, _28046_);
  nor (_28056_, _28054_, _28040_);
  nor (_28058_, _28056_, _27908_);
  nor (_28060_, _28058_, _28030_);
  nor (_28062_, _28060_, _27902_);
  nor (_28064_, _26555_, _26223_);
  not (_28066_, _27969_);
  nor (_28068_, _27318_, _27861_);
  not (_28070_, _28068_);
  not (_28072_, _27478_);
  nand (_28074_, _28072_, _28070_);
  nand (_28076_, _28074_, _27466_);
  nor (_28078_, _28074_, _27466_);
  nor (_28080_, _28078_, _27508_);
  nand (_28082_, _28080_, _28076_);
  nand (_28084_, _27020_, _27277_);
  nor (_28086_, _27024_, _26838_);
  not (_28088_, _28086_);
  nand (_28090_, _27032_, _01722_);
  nand (_28092_, _28090_, _28088_);
  not (_28094_, _28092_);
  nand (_28096_, _28094_, _28084_);
  nor (_28098_, _28096_, _27318_);
  nor (_28100_, _28098_, _26927_);
  not (_28102_, _23686_);
  nand (_28104_, _26976_, _28102_);
  not (_28106_, _06167_);
  nand (_28109_, _28106_, _06135_);
  nand (_28111_, _28109_, _28104_);
  nand (_28113_, _28111_, _26986_);
  not (_28115_, _06117_);
  nand (_28117_, _26971_, _28115_);
  nand (_28119_, _28117_, _28113_);
  nor (_28121_, _27077_, _28119_);
  nor (_28123_, _28092_, _28121_);
  nor (_28125_, _28123_, _27476_);
  nor (_28127_, _28125_, _28098_);
  not (_28129_, _28127_);
  nor (_28131_, _28129_, _27057_);
  nor (_28133_, _28131_, _28100_);
  not (_28135_, _28133_);
  nor (_28137_, _28123_, _27526_);
  nor (_28139_, _28137_, _28135_);
  nand (_28141_, _28139_, _28082_);
  not (_28143_, _28125_);
  nor (_28145_, _28143_, _27548_);
  not (_28147_, _28145_);
  nor (_28149_, _27570_, _27476_);
  nor (_28151_, _27576_, _27318_);
  nor (_28153_, _28151_, _28149_);
  nand (_28155_, _28153_, _28147_);
  nor (_28157_, _28155_, _28141_);
  nor (_28159_, _28157_, _28066_);
  not (_28161_, _26832_);
  nand (_28163_, _27997_, _30951_);
  nand (_28165_, _27985_, _30855_);
  not (_28167_, _28165_);
  nor (_28169_, _28159_, _28167_);
  not (_28171_, _28169_);
  nor (_28173_, _28171_, _28163_);
  nor (_28175_, _28169_, _27995_);
  nor (_28177_, _28175_, _28173_);
  nor (_28179_, _28177_, _26586_);
  nor (_28181_, _28179_, _28161_);
  nor (_28183_, _28181_, _27969_);
  nor (_28185_, _28183_, _28159_);
  not (_28187_, _28185_);
  nand (_28190_, _28187_, _27947_);
  not (_28192_, _28190_);
  nor (_28194_, _28192_, _28064_);
  not (_28196_, _06441_);
  nor (_28198_, _27768_, _28196_);
  not (_28200_, _06506_);
  nor (_28202_, _27803_, _28200_);
  nor (_28204_, _28202_, _28198_);
  not (_28206_, _06549_);
  nor (_28208_, _27811_, _28206_);
  not (_28210_, _06613_);
  nor (_28212_, _27778_, _28210_);
  nor (_28214_, _28212_, _28208_);
  nand (_28216_, _28214_, _28204_);
  not (_28218_, _06592_);
  nor (_28220_, _27817_, _28218_);
  not (_28222_, _06528_);
  nor (_28224_, _27795_, _28222_);
  nor (_28226_, _28224_, _28220_);
  not (_28228_, _06444_);
  nor (_28230_, _27760_, _28228_);
  not (_28232_, _06570_);
  nor (_28234_, _27785_, _28232_);
  nor (_28236_, _28234_, _28230_);
  nand (_28238_, _28236_, _28226_);
  nor (_28240_, _28238_, _28216_);
  nor (_28242_, _28240_, _27754_);
  not (_28244_, _28157_);
  nand (_28246_, _27754_, _28244_);
  not (_28248_, _28246_);
  nor (_28250_, _28248_, _28242_);
  nor (_28252_, _28250_, _26559_);
  nor (_28254_, _28017_, _26126_);
  nor (_28256_, _28254_, _28252_);
  nand (_28258_, _28256_, _28194_);
  nor (_28260_, _28258_, _28062_);
  nor (_28262_, _28260_, _28028_);
  not (_28264_, _28262_);
  not (_28266_, _03131_);
  nor (_28268_, _26935_, _28266_);
  not (_28271_, _03047_);
  nor (_28273_, _26943_, _28271_);
  nor (_28275_, _28273_, _28268_);
  nor (_28277_, _26957_, _26713_);
  nor (_28279_, _26951_, _26703_);
  nor (_28281_, _28279_, _28277_);
  nand (_28283_, _28281_, _28275_);
  not (_28285_, _26967_);
  nand (_28287_, _27196_, _26986_);
  not (_28289_, _04368_);
  nand (_28291_, _26971_, _28289_);
  nand (_28293_, _28291_, _28287_);
  nor (_28295_, _28293_, _28285_);
  nand (_28297_, _26996_, _03138_);
  not (_28299_, _28297_);
  not (_28301_, _01678_);
  nor (_28303_, _27004_, _28301_);
  nor (_28305_, _28303_, _28299_);
  not (_28307_, _28305_);
  nor (_28309_, _28307_, _28295_);
  not (_28311_, _28309_);
  nor (_28313_, _28311_, _28283_);
  not (_28315_, _28313_);
  nor (_28317_, _27077_, _28293_);
  nor (_28319_, _27024_, _26703_);
  not (_28321_, _28319_);
  nand (_28323_, _27032_, _01678_);
  nand (_28325_, _28323_, _28321_);
  nor (_28327_, _28325_, _28317_);
  not (_28329_, _28327_);
  nor (_28331_, _28329_, _28315_);
  not (_28333_, _28331_);
  nor (_28335_, _28327_, _28313_);
  not (_28337_, _28335_);
  nand (_28339_, _28337_, _27055_);
  nand (_28341_, _28339_, _26927_);
  nand (_28343_, _28341_, _28333_);
  nand (_28345_, _27016_, _27407_);
  not (_28347_, _03119_);
  nor (_28349_, _26935_, _28347_);
  not (_28353_, _03083_);
  nor (_28355_, _26943_, _28353_);
  nor (_28357_, _28355_, _28349_);
  nor (_28359_, _26951_, _26659_);
  nor (_28361_, _26957_, _26669_);
  nor (_28363_, _28361_, _28359_);
  nand (_28365_, _28363_, _28357_);
  nor (_28367_, _06135_, _23690_);
  nor (_28369_, _06174_, _26976_);
  nor (_28371_, _28369_, _28367_);
  nor (_28373_, _28371_, _26971_);
  nor (_28375_, _26986_, _06128_);
  nor (_28377_, _28375_, _28373_);
  nand (_28379_, _28377_, _26967_);
  nand (_28381_, _27006_, _01703_);
  nand (_28383_, _26996_, _03278_);
  nand (_28385_, _28383_, _28381_);
  not (_28387_, _28385_);
  nand (_28389_, _28387_, _28379_);
  nor (_28391_, _28389_, _28365_);
  not (_28393_, _28391_);
  nor (_28395_, _28393_, _28345_);
  nor (_28397_, _28395_, _27466_);
  nand (_28399_, _27482_, _27018_);
  nor (_28401_, _28399_, _28391_);
  nor (_28403_, _28401_, _27225_);
  nor (_28405_, _28403_, _28397_);
  not (_28407_, _03122_);
  nor (_28409_, _26935_, _28407_);
  not (_28411_, _03085_);
  nor (_28413_, _26943_, _28411_);
  nor (_28415_, _28413_, _28409_);
  nor (_28417_, _26951_, _26731_);
  nor (_28419_, _26957_, _26741_);
  nor (_28421_, _28419_, _28417_);
  nand (_28423_, _28421_, _28415_);
  nand (_28425_, _27176_, _26986_);
  nor (_28427_, _26986_, _06131_);
  not (_28429_, _28427_);
  nand (_28431_, _28429_, _28425_);
  nor (_28434_, _28431_, _28285_);
  not (_28436_, _01740_);
  nor (_28438_, _27004_, _28436_);
  nand (_28440_, _26996_, _03280_);
  not (_28442_, _28440_);
  nor (_28444_, _28442_, _28438_);
  not (_28446_, _28444_);
  nor (_28448_, _28446_, _28434_);
  not (_28450_, _28448_);
  nor (_28452_, _28450_, _28423_);
  not (_28454_, _28452_);
  nor (_28456_, _28454_, _27225_);
  nor (_28458_, _28452_, _27466_);
  nor (_28460_, _28458_, _28456_);
  nand (_28461_, _28460_, _28405_);
  not (_28462_, _28461_);
  nor (_28463_, _28462_, _28315_);
  nor (_28464_, _28461_, _28313_);
  nor (_28465_, _28464_, _27508_);
  not (_28466_, _28465_);
  nor (_28467_, _28466_, _28463_);
  nor (_28468_, _28329_, _27466_);
  nor (_28469_, _27225_, _28315_);
  nor (_28470_, _28469_, _27526_);
  not (_28471_, _28470_);
  nor (_28472_, _28471_, _28468_);
  nor (_28473_, _28472_, _28467_);
  nand (_28474_, _28473_, _28343_);
  nor (_28475_, _27548_, _28337_);
  not (_28476_, _28475_);
  nor (_28477_, _27570_, _28313_);
  nor (_28478_, _27576_, _28315_);
  nor (_28479_, _28478_, _28477_);
  nand (_28480_, _28479_, _28476_);
  nor (_28481_, _28480_, _28474_);
  not (_28482_, _28481_);
  nor (_28483_, _28482_, _27985_);
  nand (_28484_, _27985_, _30868_);
  not (_28485_, _28484_);
  nor (_28486_, _27478_, _27225_);
  nor (_28488_, _28068_, _27466_);
  nor (_28489_, _28488_, _28486_);
  nand (_28490_, _28489_, _27358_);
  nor (_28491_, _28489_, _27358_);
  nor (_28492_, _28491_, _27508_);
  nand (_28493_, _28492_, _28490_);
  nand (_28494_, _27020_, _27324_);
  nor (_28495_, _27024_, _26814_);
  not (_28496_, _28495_);
  nand (_28497_, _27032_, _01718_);
  nand (_28498_, _28497_, _28496_);
  not (_28499_, _28498_);
  nand (_28500_, _28499_, _28494_);
  nor (_28501_, _28500_, _27358_);
  nor (_28502_, _28501_, _26927_);
  not (_28503_, _03301_);
  nor (_28504_, _26935_, _28503_);
  nor (_28505_, _27348_, _28504_);
  nand (_28506_, _28505_, _27344_);
  not (_28507_, _27334_);
  nor (_28508_, _27350_, _28507_);
  nand (_28509_, _28508_, _27326_);
  nor (_28510_, _28509_, _28506_);
  not (_28511_, _23687_);
  nand (_28512_, _26976_, _28511_);
  not (_28513_, _06169_);
  nand (_28514_, _28513_, _06135_);
  nand (_28515_, _28514_, _28512_);
  nand (_28516_, _28515_, _26986_);
  not (_28517_, _06119_);
  nand (_28518_, _26971_, _28517_);
  nand (_28519_, _28518_, _28516_);
  nor (_28520_, _27077_, _28519_);
  nor (_28521_, _28498_, _28520_);
  nor (_28522_, _28521_, _28510_);
  nor (_28523_, _28522_, _28501_);
  not (_28524_, _28523_);
  nor (_28525_, _28524_, _27057_);
  nor (_28526_, _28525_, _28502_);
  not (_28527_, _28526_);
  nor (_28529_, _28521_, _27526_);
  nor (_28530_, _28529_, _28527_);
  nand (_28531_, _28530_, _28493_);
  nor (_28532_, _27570_, _28510_);
  not (_28533_, _28522_);
  nor (_28534_, _28533_, _27548_);
  nor (_28535_, _27576_, _27358_);
  nor (_28536_, _28535_, _28534_);
  not (_28537_, _28536_);
  nor (_28538_, _28537_, _28532_);
  not (_28539_, _28538_);
  nor (_28540_, _28539_, _28531_);
  nor (_28541_, _28540_, _28066_);
  nor (_28542_, _28541_, _28485_);
  nand (_28543_, _28542_, _28173_);
  nor (_28544_, _27987_, _26561_);
  not (_28545_, _28544_);
  nand (_28546_, _27742_, _27969_);
  nand (_28547_, _28546_, _28545_);
  nor (_28548_, _28547_, _28543_);
  not (_28549_, _30873_);
  nor (_28550_, _27987_, _28549_);
  nor (_28551_, _27584_, _28066_);
  nor (_28552_, _28551_, _28550_);
  nand (_28553_, _28552_, _28548_);
  nor (_28554_, _27987_, _26646_);
  not (_28555_, _27528_);
  nand (_28556_, _27484_, _28345_);
  nand (_28557_, _28556_, _28555_);
  not (_28558_, _28557_);
  nand (_28559_, _28558_, _28391_);
  nand (_28560_, _28557_, _28393_);
  nand (_28561_, _28560_, _28559_);
  nand (_28562_, _28561_, _27506_);
  nand (_28563_, _27020_, _28377_);
  nor (_28564_, _27024_, _26659_);
  not (_28565_, _28564_);
  nand (_28566_, _27032_, _01703_);
  nand (_28567_, _28566_, _28565_);
  not (_28568_, _28567_);
  nand (_28570_, _28568_, _28563_);
  nor (_28571_, _28570_, _28393_);
  nor (_28572_, _28571_, _26927_);
  nand (_28573_, _27148_, _26986_);
  not (_28574_, _06128_);
  nand (_28575_, _26971_, _28574_);
  nand (_28576_, _28575_, _28573_);
  nor (_28577_, _27077_, _28576_);
  nor (_28578_, _28567_, _28577_);
  nor (_28579_, _28578_, _28391_);
  nor (_28580_, _28579_, _28571_);
  not (_28581_, _28580_);
  nor (_28582_, _28581_, _27057_);
  nor (_28583_, _28582_, _28572_);
  not (_28584_, _28583_);
  nor (_28585_, _28578_, _27466_);
  nor (_28586_, _28391_, _27225_);
  nor (_28587_, _28586_, _28585_);
  nor (_28588_, _28587_, _27526_);
  nor (_28589_, _28588_, _28584_);
  nand (_28590_, _28589_, _28562_);
  not (_28591_, _28579_);
  nor (_28592_, _28591_, _27548_);
  not (_28593_, _28592_);
  nor (_28594_, _27570_, _28391_);
  nor (_28595_, _27576_, _28393_);
  nor (_28596_, _28595_, _28594_);
  nand (_28597_, _28596_, _28593_);
  nor (_28598_, _28597_, _28590_);
  nor (_28599_, _28598_, _28066_);
  nor (_28600_, _28599_, _28554_);
  not (_28601_, _28600_);
  nor (_28602_, _28601_, _28553_);
  not (_28603_, _30878_);
  nor (_28604_, _27987_, _28603_);
  nor (_28605_, _27077_, _28431_);
  nor (_28606_, _27024_, _26731_);
  not (_28607_, _28606_);
  nand (_28608_, _27032_, _01740_);
  nand (_28609_, _28608_, _28607_);
  nor (_28611_, _28609_, _28605_);
  not (_28612_, _28611_);
  nor (_28613_, _28612_, _28454_);
  nor (_28614_, _28611_, _28452_);
  nor (_28615_, _28614_, _28613_);
  not (_28616_, _28615_);
  nor (_28617_, _28616_, _27057_);
  nor (_28618_, _28613_, _26927_);
  nor (_28619_, _28618_, _28617_);
  nor (_28620_, _28452_, _28405_);
  not (_28621_, _28405_);
  nor (_28622_, _28454_, _28621_);
  nor (_28623_, _28622_, _28620_);
  nor (_28624_, _28623_, _27508_);
  nor (_28625_, _28612_, _27466_);
  not (_28626_, _28625_);
  nor (_28627_, _27526_, _28456_);
  nand (_28628_, _28627_, _28626_);
  not (_28629_, _28628_);
  nor (_28630_, _28629_, _28624_);
  nand (_28631_, _28630_, _28619_);
  not (_28632_, _28614_);
  nor (_28633_, _28632_, _27548_);
  not (_28634_, _28633_);
  nor (_28635_, _27570_, _28452_);
  nor (_28636_, _27576_, _28454_);
  nor (_28637_, _28636_, _28635_);
  nand (_28638_, _28637_, _28634_);
  nor (_28639_, _28638_, _28631_);
  nor (_28640_, _28639_, _28066_);
  nor (_28641_, _28640_, _28604_);
  nand (_28642_, _28641_, _28602_);
  nor (_28643_, _27987_, _26693_);
  nor (_28644_, _28643_, _28642_);
  nand (_28645_, _28169_, _27995_);
  not (_28646_, _28542_);
  nor (_28647_, _28646_, _28645_);
  nor (_28648_, _27718_, _28066_);
  nor (_28649_, _28648_, _28544_);
  nand (_28650_, _28649_, _28647_);
  not (_28652_, _28552_);
  nor (_28653_, _28652_, _28650_);
  nand (_28654_, _28600_, _28653_);
  not (_28655_, _28641_);
  nor (_28656_, _28655_, _28654_);
  not (_28657_, _28643_);
  nor (_28658_, _28657_, _28656_);
  nor (_28659_, _28658_, _28644_);
  nor (_28660_, _28659_, _26586_);
  nor (_28661_, _27987_, _26701_);
  not (_28662_, _28661_);
  nor (_28663_, _28662_, _28660_);
  nor (_28664_, _28663_, _28483_);
  nand (_28665_, _28664_, _27947_);
  nor (_28666_, _25609_, _26703_);
  not (_28667_, _06072_);
  nor (_28668_, _25643_, _28667_);
  nor (_28669_, _25621_, _25714_);
  nor (_28670_, _28669_, _28668_);
  not (_28671_, _28670_);
  nor (_28672_, _25663_, _25718_);
  not (_28673_, _04660_);
  nor (_28674_, _25676_, _28673_);
  nor (_28675_, _28674_, _28672_);
  nor (_28676_, _25631_, _25736_);
  not (_28677_, _06063_);
  nor (_28678_, _25657_, _28677_);
  nor (_28679_, _28678_, _28676_);
  nand (_28680_, _28679_, _28675_);
  nor (_28681_, _28680_, _28671_);
  nor (_28682_, _27908_, _28681_);
  nor (_28683_, _28682_, _28666_);
  not (_28684_, _28683_);
  nand (_28685_, _28684_, _27900_);
  nand (_28686_, _28685_, _26223_);
  not (_28687_, _06384_);
  nor (_28688_, _27795_, _28687_);
  not (_28689_, _06376_);
  nor (_28690_, _27803_, _28689_);
  nor (_28691_, _28690_, _28688_);
  not (_28693_, _06392_);
  nor (_28694_, _27785_, _28693_);
  not (_28695_, _06388_);
  nor (_28696_, _27811_, _28695_);
  nor (_28697_, _28696_, _28694_);
  nand (_28698_, _28697_, _28691_);
  not (_28699_, _06380_);
  nor (_28700_, _27760_, _28699_);
  not (_28701_, _06359_);
  nor (_28702_, _27768_, _28701_);
  nor (_28703_, _28702_, _28700_);
  not (_28704_, _06398_);
  nor (_28705_, _27817_, _28704_);
  not (_28706_, _06402_);
  nor (_28707_, _27778_, _28706_);
  nor (_28708_, _28707_, _28705_);
  nand (_28709_, _28708_, _28703_);
  nor (_28710_, _28709_, _28698_);
  nor (_28711_, _28710_, _27754_);
  nand (_28712_, _27754_, _28482_);
  not (_28713_, _28712_);
  nor (_28714_, _28713_, _28711_);
  nor (_28715_, _28714_, _26555_);
  nor (_28716_, _28715_, _28686_);
  nand (_28717_, _28716_, _28665_);
  not (_28718_, _28717_);
  nor (_28719_, _28017_, _27590_);
  nor (_28720_, _25609_, _26618_);
  not (_28721_, _05491_);
  nor (_28722_, _25643_, _28721_);
  nor (_28723_, _25621_, _25637_);
  nor (_28724_, _28723_, _28722_);
  not (_28725_, _28724_);
  nor (_28726_, _25657_, _25669_);
  nor (_28727_, _25676_, _25625_);
  nor (_28728_, _28727_, _28726_);
  nor (_28729_, _25663_, _25651_);
  nor (_28730_, _25631_, _25617_);
  nor (_28731_, _28730_, _28729_);
  nand (_28732_, _28731_, _28728_);
  nor (_28734_, _28732_, _28725_);
  nor (_28735_, _28734_, _27908_);
  nor (_28736_, _28735_, _28720_);
  nor (_28737_, _28736_, _27902_);
  nor (_28738_, _28737_, _28719_);
  not (_28739_, _28738_);
  not (_28740_, _06580_);
  nor (_28741_, _27785_, _28740_);
  not (_28742_, _06537_);
  nor (_28743_, _27795_, _28742_);
  nor (_28744_, _28743_, _28741_);
  not (_28745_, _06422_);
  nor (_28746_, _27768_, _28745_);
  not (_28747_, _06622_);
  nor (_28748_, _27778_, _28747_);
  nor (_28749_, _28748_, _28746_);
  nand (_28750_, _28749_, _28744_);
  not (_28751_, _06516_);
  nor (_28752_, _27803_, _28751_);
  not (_28753_, _06489_);
  nor (_28754_, _27760_, _28753_);
  nor (_28755_, _28754_, _28752_);
  not (_28756_, _06558_);
  nor (_28757_, _27811_, _28756_);
  not (_28758_, _06601_);
  nor (_28759_, _27817_, _28758_);
  nor (_28760_, _28759_, _28757_);
  nand (_28761_, _28760_, _28755_);
  nor (_28762_, _28761_, _28750_);
  nor (_28763_, _28762_, _27754_);
  nor (_28764_, _27890_, _27584_);
  nor (_28765_, _28764_, _28763_);
  not (_28766_, _28765_);
  nand (_28767_, _28766_, _26557_);
  not (_28768_, _27947_);
  nor (_28769_, _28552_, _28548_);
  nor (_28770_, _28769_, _28653_);
  nor (_28771_, _28770_, _26586_);
  nor (_28772_, _28771_, _26592_);
  nor (_28773_, _28772_, _27969_);
  nor (_28775_, _28773_, _28551_);
  nor (_28776_, _28775_, _28768_);
  nor (_28777_, _26553_, _26223_);
  nor (_28778_, _28777_, _28776_);
  nand (_28779_, _28778_, _28767_);
  nor (_28780_, _28779_, _28739_);
  not (_28781_, _28780_);
  nor (_28782_, _28781_, _28718_);
  nor (_28783_, _28641_, _28602_);
  nor (_28784_, _28783_, _28656_);
  nor (_28785_, _28784_, _26586_);
  nor (_28786_, _28785_, _26727_);
  nor (_28787_, _28786_, _27969_);
  nor (_28788_, _28787_, _28640_);
  nor (_28789_, _28788_, _28768_);
  not (_28790_, _06411_);
  nor (_28791_, _27768_, _28790_);
  not (_28792_, _06628_);
  nor (_28793_, _27778_, _28792_);
  nor (_28794_, _28793_, _28791_);
  not (_28795_, _06564_);
  nor (_28796_, _27811_, _28795_);
  not (_28797_, _06522_);
  nor (_28798_, _27803_, _28797_);
  nor (_28799_, _28798_, _28796_);
  nand (_28800_, _28799_, _28794_);
  not (_28801_, _06607_);
  nor (_28802_, _27817_, _28801_);
  not (_28803_, _06543_);
  nor (_28804_, _27795_, _28803_);
  nor (_28805_, _28804_, _28802_);
  not (_28806_, _06495_);
  nor (_28807_, _27760_, _28806_);
  not (_28808_, _06586_);
  nor (_28809_, _27785_, _28808_);
  nor (_28810_, _28809_, _28807_);
  nand (_28811_, _28810_, _28805_);
  nor (_28812_, _28811_, _28800_);
  nor (_28813_, _28812_, _27754_);
  nor (_28814_, _27890_, _28639_);
  nor (_28817_, _28814_, _28813_);
  nor (_28818_, _28817_, _26559_);
  not (_28819_, _26555_);
  nor (_28820_, _28819_, _26223_);
  not (_28821_, _27900_);
  nor (_28822_, _25609_, _26731_);
  not (_28823_, _05497_);
  nor (_28824_, _25643_, _28823_);
  nor (_28825_, _25621_, _25771_);
  nor (_28826_, _28825_, _28824_);
  not (_28827_, _28826_);
  nor (_28828_, _25663_, _25781_);
  not (_28829_, _05427_);
  nor (_28830_, _25676_, _28829_);
  nor (_28831_, _28830_, _28828_);
  nor (_28832_, _25631_, _25777_);
  nor (_28833_, _25657_, _25791_);
  nor (_28834_, _28833_, _28832_);
  nand (_28835_, _28834_, _28831_);
  nor (_28836_, _28835_, _28827_);
  nor (_28837_, _28836_, _27908_);
  nor (_28838_, _28837_, _28822_);
  nor (_28839_, _28838_, _28821_);
  nor (_28840_, _28839_, _28820_);
  not (_28841_, _28840_);
  nor (_28842_, _28841_, _28818_);
  not (_28843_, _28842_);
  nor (_28844_, _28843_, _28789_);
  not (_28845_, _28844_);
  not (_28846_, _06604_);
  nor (_28847_, _27817_, _28846_);
  not (_28848_, _06415_);
  nor (_28849_, _27768_, _28848_);
  nor (_28850_, _28849_, _28847_);
  not (_28851_, _06492_);
  nor (_28852_, _27760_, _28851_);
  not (_28853_, _06540_);
  nor (_28854_, _27795_, _28853_);
  nor (_28855_, _28854_, _28852_);
  nand (_28856_, _28855_, _28850_);
  not (_28858_, _06519_);
  nor (_28859_, _27803_, _28858_);
  not (_28860_, _06583_);
  nor (_28861_, _27785_, _28860_);
  nor (_28862_, _28861_, _28859_);
  not (_28863_, _06561_);
  nor (_28864_, _27811_, _28863_);
  not (_28865_, _06625_);
  nor (_28866_, _27778_, _28865_);
  nor (_28867_, _28866_, _28864_);
  nand (_28868_, _28867_, _28862_);
  nor (_28869_, _28868_, _28856_);
  nor (_28870_, _28869_, _27754_);
  nor (_28871_, _27890_, _28598_);
  nor (_28872_, _28871_, _28870_);
  nor (_28873_, _28872_, _26559_);
  nor (_28874_, _25609_, _26659_);
  not (_28875_, _05493_);
  nor (_28876_, _25643_, _28875_);
  not (_28877_, _05461_);
  nor (_28878_, _25621_, _28877_);
  nor (_28879_, _28878_, _28876_);
  not (_28880_, _28879_);
  nor (_28881_, _25657_, _25846_);
  not (_28882_, _05422_);
  nor (_28883_, _25676_, _28882_);
  nor (_28884_, _28883_, _28881_);
  nor (_28885_, _25663_, _25850_);
  nor (_28886_, _25631_, _25835_);
  nor (_28887_, _28886_, _28885_);
  nand (_28888_, _28887_, _28884_);
  nor (_28889_, _28888_, _28880_);
  nor (_28890_, _28889_, _27908_);
  nor (_28891_, _28890_, _28874_);
  nor (_28892_, _28891_, _27902_);
  nor (_28893_, _28892_, _28873_);
  nor (_28894_, _28600_, _28653_);
  nor (_28895_, _28894_, _28602_);
  nor (_28896_, _28895_, _26586_);
  nor (_28897_, _28896_, _26655_);
  nor (_28899_, _28897_, _27969_);
  nor (_28900_, _28899_, _28599_);
  nor (_28901_, _28900_, _28768_);
  nand (_28902_, _28820_, _28821_);
  not (_28903_, _28902_);
  nor (_28904_, _28903_, _28901_);
  nand (_28905_, _28904_, _28893_);
  nor (_28906_, _28905_, _28845_);
  nand (_28907_, _28906_, _28782_);
  nor (_28908_, _28649_, _28647_);
  nor (_28909_, _28908_, _28548_);
  nor (_28910_, _28909_, _26586_);
  nor (_28911_, _28910_, _26767_);
  nor (_28912_, _28911_, _27969_);
  nor (_28913_, _28912_, _28648_);
  not (_28914_, _28913_);
  nand (_28915_, _28914_, _27947_);
  nor (_28916_, _28017_, _27722_);
  not (_28917_, _28916_);
  nand (_28918_, _28917_, _28915_);
  not (_28919_, _06577_);
  nor (_28920_, _27785_, _28919_);
  not (_28921_, _06534_);
  nor (_28922_, _27795_, _28921_);
  nor (_28923_, _28922_, _28920_);
  not (_28924_, _06426_);
  nor (_28925_, _27768_, _28924_);
  not (_28926_, _06598_);
  nor (_28927_, _27817_, _28926_);
  nor (_28928_, _28927_, _28925_);
  nand (_28929_, _28928_, _28923_);
  not (_28930_, _06512_);
  nor (_28931_, _27803_, _28930_);
  not (_28932_, _06479_);
  nor (_28933_, _27760_, _28932_);
  nor (_28934_, _28933_, _28931_);
  not (_28935_, _06555_);
  nor (_28936_, _27811_, _28935_);
  not (_28937_, _06619_);
  nor (_28938_, _27778_, _28937_);
  nor (_28940_, _28938_, _28936_);
  nand (_28941_, _28940_, _28934_);
  nor (_28942_, _28941_, _28929_);
  nor (_28943_, _28942_, _27754_);
  nand (_28944_, _27754_, _27742_);
  not (_28945_, _28944_);
  nor (_28946_, _28945_, _28943_);
  not (_28947_, _28946_);
  nand (_28948_, _28947_, _26557_);
  not (_28949_, _27902_);
  nor (_28950_, _25609_, _26757_);
  not (_28951_, _05478_);
  nor (_28952_, _25643_, _28951_);
  not (_28953_, _05457_);
  nor (_28954_, _25621_, _28953_);
  nor (_28955_, _28954_, _28952_);
  not (_28956_, _28955_);
  nor (_28957_, _25657_, _26025_);
  nor (_28958_, _25676_, _26017_);
  nor (_28959_, _28958_, _28957_);
  nor (_28960_, _25663_, _26029_);
  nor (_28961_, _25631_, _26039_);
  nor (_28962_, _28961_, _28960_);
  nand (_28963_, _28962_, _28959_);
  nor (_28964_, _28963_, _28956_);
  nor (_28965_, _28964_, _27908_);
  nor (_28966_, _28965_, _28950_);
  not (_28967_, _28966_);
  nand (_28968_, _28967_, _28949_);
  nand (_28969_, _28968_, _28948_);
  nor (_28970_, _28969_, _28918_);
  not (_28971_, _28970_);
  not (_28972_, _26801_);
  nor (_28973_, _28542_, _28173_);
  nor (_28974_, _28973_, _28647_);
  nor (_28975_, _28974_, _26586_);
  nor (_28976_, _28975_, _28972_);
  nor (_28977_, _28976_, _27969_);
  nor (_28978_, _28977_, _28541_);
  nor (_28979_, _28978_, _28768_);
  nor (_28981_, _28017_, _26201_);
  nor (_28982_, _28981_, _28979_);
  not (_28983_, _06616_);
  nor (_28984_, _27778_, _28983_);
  not (_28985_, _06595_);
  nor (_28986_, _27817_, _28985_);
  nor (_28987_, _28986_, _28984_);
  not (_28988_, _06406_);
  nor (_28989_, _27768_, _28988_);
  not (_28990_, _06573_);
  nor (_28991_, _27785_, _28990_);
  nor (_28992_, _28991_, _28989_);
  nand (_28993_, _28992_, _28987_);
  not (_28994_, _06531_);
  nor (_28995_, _27795_, _28994_);
  not (_28996_, _06509_);
  nor (_28997_, _27803_, _28996_);
  nor (_28998_, _28997_, _28995_);
  not (_28999_, _06476_);
  nor (_29000_, _27760_, _28999_);
  not (_29001_, _06552_);
  nor (_29002_, _27811_, _29001_);
  nor (_29003_, _29002_, _29000_);
  nand (_29004_, _29003_, _28998_);
  nor (_29005_, _29004_, _28993_);
  nor (_29006_, _29005_, _27754_);
  nor (_29007_, _27890_, _28540_);
  nor (_29008_, _29007_, _29006_);
  nor (_29009_, _29008_, _26559_);
  nor (_29010_, _25609_, _26814_);
  not (_29011_, _05472_);
  nor (_29012_, _25643_, _29011_);
  not (_29013_, _05455_);
  nor (_29014_, _25621_, _29013_);
  nor (_29015_, _29014_, _29012_);
  not (_29016_, _29015_);
  nor (_29017_, _25663_, _25970_);
  nor (_29018_, _25676_, _25958_);
  nor (_29019_, _29018_, _29017_);
  nor (_29020_, _25631_, _25980_);
  nor (_29022_, _25657_, _25966_);
  nor (_29023_, _29022_, _29020_);
  nand (_29024_, _29023_, _29019_);
  nor (_29025_, _29024_, _29016_);
  nor (_29026_, _29025_, _27908_);
  nor (_29027_, _29026_, _29010_);
  nor (_29028_, _29027_, _27902_);
  nor (_29029_, _29028_, _29009_);
  nand (_29030_, _29029_, _28982_);
  nor (_29031_, _29030_, _28971_);
  not (_29032_, _29031_);
  nor (_29033_, _29032_, _28907_);
  not (_29034_, _29033_);
  nor (_29035_, _29034_, _28264_);
  not (_29036_, _29035_);
  not (_29037_, _03815_);
  nand (_29038_, _03360_, _25592_);
  nor (_29039_, _29038_, _29037_);
  not (_29040_, _29039_);
  nor (_29041_, _29040_, _29036_);
  nor (_29042_, _29030_, _28970_);
  not (_29043_, _29042_);
  nor (_29044_, _29043_, _28264_);
  not (_29045_, _29044_);
  nor (_29046_, _28905_, _28844_);
  nand (_29047_, _29046_, _28782_);
  nor (_29048_, _29047_, _29045_);
  nand (_29049_, _29048_, _01459_);
  not (_29050_, _28013_);
  nor (_29051_, _29050_, _27942_);
  nand (_29052_, _29051_, _28021_);
  nor (_29053_, _29052_, _27896_);
  not (_29054_, _28260_);
  nor (_29055_, _29054_, _29053_);
  not (_29056_, _29055_);
  not (_29057_, _29030_);
  nor (_29058_, _29057_, _28970_);
  not (_29059_, _29058_);
  nor (_29060_, _29059_, _29056_);
  not (_29061_, _29060_);
  nor (_29063_, _29047_, _29061_);
  nand (_29064_, _29063_, _01265_);
  nand (_29065_, _29064_, _29049_);
  nor (_29066_, _29054_, _28028_);
  not (_29067_, _29066_);
  nor (_29068_, _29067_, _29043_);
  not (_29069_, _29068_);
  nor (_29070_, _29069_, _29047_);
  nand (_29071_, _29070_, _01249_);
  nor (_29072_, _29067_, _29059_);
  not (_29073_, _29072_);
  nor (_29074_, _29073_, _29047_);
  nand (_29075_, _29074_, _01369_);
  nand (_29076_, _29075_, _29071_);
  nor (_29077_, _29076_, _29065_);
  nor (_29078_, _28260_, _29053_);
  not (_29079_, _29078_);
  nor (_29080_, _29079_, _29043_);
  not (_29081_, _29080_);
  nor (_29082_, _29081_, _29047_);
  nand (_29083_, _29082_, _01488_);
  nor (_29084_, _29069_, _28907_);
  nand (_29085_, _29084_, _30981_);
  nand (_29086_, _29085_, _29083_);
  nor (_29087_, _28845_, _28718_);
  not (_29088_, _29087_);
  not (_29089_, _28905_);
  nor (_29090_, _29089_, _28781_);
  not (_29091_, _29090_);
  nor (_29092_, _29091_, _29088_);
  nand (_29093_, _29092_, _29068_);
  not (_29094_, _29093_);
  nand (_29095_, _29094_, _00390_);
  nor (_29096_, _29079_, _29057_);
  not (_29097_, _29096_);
  nor (_29098_, _29097_, _28971_);
  nor (_29099_, _29089_, _28780_);
  not (_29100_, _29099_);
  nor (_29101_, _29100_, _29088_);
  nand (_29102_, _29101_, _29098_);
  not (_29104_, _29102_);
  nand (_29105_, _29104_, _00402_);
  nand (_29106_, _29105_, _29095_);
  nor (_29107_, _29106_, _29086_);
  nand (_29108_, _29107_, _29077_);
  nor (_29109_, _29045_, _28907_);
  nand (_29110_, _29109_, _31254_);
  nor (_29111_, _29061_, _28907_);
  nand (_29112_, _29111_, _31268_);
  nand (_29113_, _29112_, _29110_);
  nor (_29114_, _29081_, _28907_);
  nand (_29115_, _29114_, _31290_);
  nor (_29116_, _29056_, _29043_);
  not (_29117_, _29116_);
  nor (_29118_, _29117_, _28907_);
  nand (_29119_, _29118_, _30984_);
  nand (_29120_, _29119_, _29115_);
  nor (_29121_, _29120_, _29113_);
  nor (_29122_, _28905_, _28780_);
  not (_29123_, _29122_);
  nor (_29124_, _29123_, _29088_);
  not (_29125_, _29124_);
  nor (_29126_, _29125_, _29117_);
  nand (_29127_, _29126_, _01036_);
  nor (_29128_, _29069_, _29125_);
  nand (_29129_, _29128_, _00801_);
  nand (_29130_, _29129_, _29127_);
  not (_29131_, _29098_);
  nor (_29132_, _29131_, _28907_);
  nand (_29133_, _29132_, _01197_);
  nor (_29134_, _29073_, _28907_);
  nand (_29135_, _29134_, _31018_);
  nand (_29136_, _29135_, _29133_);
  nor (_29137_, _29136_, _29130_);
  nand (_29138_, _29137_, _29121_);
  nor (_29139_, _29138_, _29108_);
  nor (_29140_, _28844_, _28718_);
  nor (_29141_, _29032_, _29067_);
  nand (_29142_, _29141_, _29140_);
  nor (_29143_, _29142_, _29123_);
  nand (_29145_, _29143_, _30666_);
  nor (_29146_, _29142_, _29091_);
  nand (_29147_, _29146_, _01740_);
  nand (_29148_, _29147_, _29145_);
  nor (_29149_, _29100_, _29142_);
  nand (_29150_, _29149_, _01609_);
  not (_29151_, _28788_);
  nand (_29152_, _29031_, _29055_);
  nor (_29153_, _29152_, _28907_);
  nand (_29154_, _29153_, _29151_);
  nand (_29155_, _29154_, _29150_);
  nor (_29156_, _29034_, _29079_);
  nand (_29157_, _29156_, _30783_);
  nand (_29158_, _29035_, _30812_);
  nand (_29159_, _29158_, _29157_);
  nor (_29160_, _29159_, _29155_);
  not (_29161_, _29092_);
  not (_29162_, _29141_);
  nor (_29163_, _29162_, _29161_);
  not (_29164_, _26347_);
  nor (_29165_, _29164_, _26327_);
  not (_29166_, _26203_);
  nor (_29167_, _29166_, _26128_);
  not (_29168_, _29167_);
  nor (_29169_, _29168_, _26274_);
  nor (_29170_, _29169_, _29165_);
  not (_29171_, _26069_);
  nor (_29172_, _29171_, _25706_);
  not (_29173_, _29172_);
  nor (_29174_, _29173_, _26422_);
  nand (_29175_, _26533_, _26069_);
  nor (_29176_, _29175_, _25706_);
  nor (_29177_, _29176_, _29174_);
  nand (_29178_, _29177_, _29170_);
  nor (_29179_, _29178_, _26282_);
  nand (_29180_, _29179_, _26258_);
  not (_29181_, _26383_);
  not (_29182_, _26355_);
  nand (_29183_, _29182_, _25708_);
  not (_29184_, _26424_);
  nand (_29186_, _29184_, _29183_);
  nor (_29187_, _29186_, _29181_);
  not (_29188_, _26393_);
  not (_29189_, _26448_);
  nor (_29190_, _29189_, _29188_);
  nor (_29191_, _29171_, _25708_);
  not (_29192_, _29191_);
  nor (_29193_, _29192_, _25769_);
  not (_29194_, _29193_);
  nor (_29195_, _29194_, _25886_);
  not (_29196_, _29195_);
  nand (_29197_, _29196_, _26501_);
  nor (_29198_, _29197_, _26408_);
  nand (_29199_, _29198_, _29190_);
  not (_29200_, _26353_);
  nor (_29201_, _26347_, _26533_);
  not (_29202_, _29201_);
  nand (_29203_, _29202_, _26316_);
  nand (_29204_, _29203_, _29200_);
  nor (_29205_, _29204_, _29199_);
  nand (_29206_, _29205_, _29187_);
  nor (_29207_, _29206_, _29180_);
  nor (_29208_, _29207_, _25601_);
  nor (_29209_, _29208_, _30591_);
  not (_29210_, _29208_);
  nor (_29211_, _29210_, _30321_);
  nor (_29212_, _29211_, _29209_);
  nand (_29213_, _29212_, _29163_);
  nor (_29214_, _29208_, _30613_);
  nor (_29215_, _29210_, _30346_);
  nor (_29216_, _29215_, _29214_);
  not (_29217_, _29101_);
  nor (_29218_, _29217_, _29162_);
  nand (_29219_, _29218_, _29216_);
  nand (_29220_, _29219_, _29213_);
  nor (_29221_, _29208_, _30570_);
  nor (_29222_, _29210_, _30313_);
  nor (_29223_, _29222_, _29221_);
  nor (_29224_, _29162_, _29125_);
  nand (_29225_, _29224_, _29223_);
  nor (_29229_, _29208_, _30549_);
  nor (_29230_, _29210_, _30409_);
  nor (_29231_, _29230_, _29229_);
  nor (_29232_, _29162_, _28907_);
  nand (_29233_, _29232_, _29231_);
  nand (_29234_, _29233_, _29225_);
  nor (_29235_, _29234_, _29220_);
  nand (_29236_, _29235_, _29160_);
  nor (_29237_, _29236_, _29148_);
  nand (_29238_, _29237_, _29139_);
  not (_29239_, _29156_);
  nor (_29240_, _29040_, _29239_);
  not (_29241_, _29143_);
  nor (_29242_, _30689_, _30685_);
  nor (_29243_, _29242_, _29241_);
  nor (_29244_, _29243_, _29240_);
  nor (_29245_, _29244_, _03332_);
  nor (_29246_, _28970_, _26777_);
  nor (_29247_, _28971_, _27726_);
  nor (_29248_, _29247_, _29246_);
  nor (_29249_, _28780_, _26640_);
  nor (_29250_, _28781_, _26642_);
  nor (_29251_, _29250_, _29249_);
  nand (_29252_, _29251_, _29248_);
  nor (_29253_, _28718_, _26721_);
  nor (_29254_, _28717_, _27608_);
  nor (_29255_, _29254_, _29253_);
  nor (_29256_, _29089_, _26679_);
  nor (_29257_, _28905_, _26677_);
  nor (_29258_, _29257_, _29256_);
  nor (_29259_, _28845_, _26749_);
  nor (_29260_, _28844_, _27610_);
  nor (_29261_, _29260_, _29259_);
  nand (_29262_, _29261_, _29258_);
  nor (_29263_, _29262_, _29255_);
  not (_29264_, _29263_);
  nor (_29265_, _29264_, _29252_);
  nor (_29266_, _29054_, _26856_);
  not (_29267_, _26826_);
  nor (_29268_, _29057_, _29267_);
  nor (_29270_, _29030_, _26826_);
  nor (_29271_, _29270_, _29268_);
  nor (_29272_, _29271_, _29266_);
  nor (_29273_, _29053_, _26884_);
  nor (_29274_, _28028_, _26886_);
  nor (_29275_, _29274_, _29273_);
  nor (_29276_, _28260_, _26858_);
  not (_29277_, _29276_);
  nand (_29278_, _29277_, _27949_);
  nor (_29279_, _29278_, _29275_);
  nand (_29280_, _29279_, _29272_);
  not (_29281_, _29280_);
  nand (_29282_, _29281_, _29265_);
  not (_29283_, _29282_);
  nor (_29284_, _26721_, _30308_);
  nand (_29285_, _29284_, _29283_);
  not (_29286_, _29146_);
  nor (_29287_, _29038_, _03815_);
  nor (_29288_, _29037_, _03332_);
  nand (_29289_, _29288_, _29038_);
  not (_29290_, _29289_);
  nor (_29291_, _29290_, _29287_);
  nor (_29292_, _29291_, _29286_);
  not (_29293_, _30308_);
  not (_29294_, _27949_);
  nor (_29295_, _29294_, _29293_);
  not (_29297_, _29295_);
  nor (_29298_, _29297_, _26721_);
  not (_29299_, _29298_);
  nor (_29300_, _29299_, _29096_);
  nand (_29301_, _29300_, _29265_);
  not (_29302_, _29301_);
  nor (_29303_, _29302_, _29292_);
  nand (_29304_, _29303_, _29285_);
  nor (_29305_, _29304_, _29245_);
  nand (_29306_, _29305_, _29238_);
  nor (_29307_, _29162_, _29088_);
  not (_29308_, _29307_);
  nor (_29309_, _29074_, _29070_);
  nand (_29310_, _29309_, _29308_);
  not (_29312_, _29048_);
  not (_29313_, _29082_);
  nand (_29314_, _29313_, _29312_);
  not (_29315_, _29063_);
  not (_29316_, _29084_);
  nand (_29317_, _29316_, _29315_);
  nor (_29318_, _29317_, _29314_);
  nand (_29319_, _29318_, _29036_);
  nor (_29320_, _29319_, _29310_);
  not (_29321_, _28907_);
  nand (_29322_, _29080_, _29321_);
  nor (_29323_, _29134_, _29111_);
  nor (_29324_, _29132_, _29109_);
  nand (_29325_, _29324_, _29323_);
  nor (_29326_, _29104_, _29118_);
  nand (_29327_, _29326_, _29093_);
  nor (_29328_, _29327_, _29325_);
  nand (_29329_, _29328_, _29322_);
  nand (_29330_, _29033_, _29055_);
  nor (_29331_, _29146_, _29143_);
  nand (_29332_, _29331_, _29330_);
  not (_29333_, _29149_);
  nor (_29334_, _29128_, _29126_);
  nand (_29335_, _29334_, _29333_);
  nor (_29336_, _29335_, _29332_);
  nand (_29337_, _29336_, _29239_);
  nor (_29338_, _29337_, _29329_);
  nand (_29339_, _29338_, _29320_);
  nand (_29340_, _29339_, _29305_);
  nand (_29341_, _29340_, _06131_);
  nand (_29342_, _29341_, _29306_);
  nor (_29343_, _29342_, _29041_);
  not (_29344_, _23698_);
  nor (_29345_, _27544_, _27052_);
  not (_29346_, _29345_);
  nor (_29347_, _28612_, _28329_);
  nor (_29348_, _29347_, _02091_);
  not (_29349_, _02093_);
  nor (_29350_, _27040_, _02091_);
  not (_29351_, _02091_);
  nor (_29353_, _28612_, _29351_);
  nor (_29354_, _29353_, _29350_);
  nor (_29355_, _28570_, _02091_);
  nor (_29356_, _28329_, _29351_);
  nor (_29357_, _29356_, _29355_);
  nor (_29358_, _29357_, _29354_);
  nor (_29359_, _27645_, _02091_);
  nor (_29360_, _28570_, _29351_);
  nor (_29361_, _29360_, _29359_);
  nor (_29362_, _28500_, _02091_);
  nor (_29363_, _27040_, _29351_);
  nor (_29364_, _29363_, _29362_);
  nor (_29365_, _29364_, _29361_);
  nand (_29366_, _29365_, _29358_);
  nand (_29367_, _29366_, _29349_);
  not (_29368_, _29367_);
  nor (_29369_, _29368_, _29348_);
  not (_29370_, _29369_);
  nor (_29371_, _28096_, _02091_);
  nor (_29372_, _27645_, _29351_);
  nor (_29373_, _29372_, _29371_);
  nor (_29374_, _29373_, _02093_);
  nor (_29375_, _29357_, _29349_);
  nor (_29376_, _29375_, _29374_);
  nor (_29377_, _02093_, _02091_);
  not (_29378_, _29377_);
  nor (_29379_, _29378_, _28315_);
  nor (_29380_, _29377_, _02096_);
  nor (_29381_, _29380_, _29379_);
  not (_29382_, _29381_);
  nand (_29383_, _27020_, _27257_);
  not (_29384_, _27847_);
  nand (_29385_, _29384_, _29383_);
  nor (_29386_, _29385_, _02091_);
  nor (_29387_, _28500_, _29351_);
  nor (_29388_, _29387_, _29386_);
  nor (_29389_, _29388_, _02093_);
  nor (_29390_, _29354_, _29349_);
  nor (_29391_, _29390_, _29389_);
  nor (_29392_, _29391_, _29382_);
  not (_29394_, _29391_);
  nor (_29395_, _29394_, _29381_);
  nor (_29396_, _29377_, _02224_);
  nor (_29397_, _29378_, _28454_);
  nor (_29398_, _29397_, _29396_);
  not (_29399_, _29398_);
  nor (_29400_, _28123_, _29351_);
  nor (_29401_, _29400_, _02093_);
  nor (_29402_, _29361_, _29349_);
  nor (_29403_, _29402_, _29401_);
  nor (_29404_, _29403_, _29399_);
  not (_29405_, _29404_);
  nor (_29406_, _29405_, _29395_);
  nor (_29407_, _29406_, _29392_);
  not (_29408_, _29407_);
  nor (_29409_, _29395_, _29392_);
  not (_29410_, _29409_);
  not (_29411_, _29403_);
  nor (_29412_, _29411_, _29398_);
  nor (_29413_, _29412_, _29404_);
  not (_29414_, _29413_);
  nor (_29415_, _29414_, _29410_);
  not (_29416_, _29415_);
  nor (_29417_, _29377_, _02222_);
  nor (_29418_, _29378_, _28393_);
  nor (_29419_, _29418_, _29417_);
  not (_29420_, _29419_);
  nor (_29421_, _27849_, _29351_);
  nor (_29422_, _29421_, _02093_);
  nor (_29423_, _29364_, _29349_);
  nor (_29424_, _29423_, _29422_);
  nor (_29425_, _29424_, _29420_);
  not (_29426_, _29424_);
  nor (_29427_, _29426_, _29419_);
  nand (_29428_, _29373_, _02093_);
  nor (_29429_, _29378_, _27018_);
  nor (_29430_, _29377_, _02220_);
  nor (_29431_, _29430_, _29429_);
  nand (_29432_, _29431_, _29428_);
  not (_29433_, _29432_);
  nand (_29435_, _29388_, _02093_);
  not (_29436_, _29435_);
  nand (_29437_, _29377_, _27403_);
  nor (_29438_, _29377_, _02218_);
  not (_29439_, _29438_);
  nand (_29440_, _29439_, _29437_);
  nor (_29441_, _29440_, _29436_);
  not (_29442_, _29440_);
  nand (_29443_, _29442_, _29435_);
  nand (_29444_, _29440_, _29436_);
  nand (_29445_, _29444_, _29443_);
  nand (_29446_, _28096_, _02091_);
  nor (_29447_, _29446_, _29349_);
  nand (_29448_, _29377_, _28510_);
  nor (_29449_, _29377_, _02216_);
  not (_29450_, _29449_);
  nand (_29451_, _29450_, _29448_);
  nor (_29452_, _29451_, _29447_);
  nand (_29453_, _29421_, _02093_);
  nor (_29454_, _29377_, _02214_);
  nor (_29455_, _29378_, _27318_);
  nor (_29456_, _29455_, _29454_);
  nor (_29457_, _29456_, _29453_);
  nand (_29458_, _29400_, _02093_);
  nor (_29459_, _29378_, _27358_);
  nor (_29460_, _29449_, _29459_);
  nand (_29461_, _29460_, _29458_);
  nand (_29462_, _29451_, _29447_);
  nand (_29463_, _29462_, _29461_);
  nor (_29464_, _29463_, _29457_);
  nor (_29465_, _29464_, _29452_);
  nor (_29466_, _29465_, _29445_);
  nor (_29467_, _29466_, _29441_);
  nor (_29468_, _29431_, _29428_);
  not (_29469_, _29468_);
  nand (_29470_, _29469_, _29432_);
  nor (_29471_, _29470_, _29467_);
  nor (_29472_, _29471_, _29433_);
  nor (_29473_, _29472_, _29427_);
  nor (_29474_, _29473_, _29425_);
  nor (_29476_, _29474_, _29416_);
  nor (_29477_, _29476_, _29408_);
  nor (_29478_, _29376_, _29370_);
  not (_29479_, _29478_);
  nor (_29480_, _29479_, _29477_);
  nor (_29481_, _29480_, _29381_);
  nor (_29482_, _29442_, _29435_);
  nor (_29483_, _29482_, _29441_);
  not (_29484_, _29453_);
  not (_29485_, _29454_);
  nand (_29486_, _29377_, _27476_);
  nand (_29487_, _29486_, _29485_);
  nand (_29488_, _29487_, _29484_);
  nor (_29489_, _29460_, _29458_);
  nor (_29490_, _29489_, _29452_);
  nand (_29491_, _29490_, _29488_);
  nand (_29492_, _29491_, _29461_);
  nand (_29493_, _29492_, _29483_);
  nand (_29494_, _29493_, _29443_);
  nor (_29495_, _29468_, _29433_);
  nand (_29496_, _29495_, _29494_);
  nand (_29497_, _29496_, _29432_);
  nor (_29498_, _29497_, _29425_);
  nor (_29499_, _29498_, _29427_);
  nand (_29500_, _29499_, _29415_);
  nand (_29501_, _29500_, _29407_);
  nand (_29502_, _29478_, _29501_);
  nor (_29503_, _29474_, _29414_);
  nor (_29504_, _29503_, _29404_);
  nor (_29505_, _29504_, _29409_);
  nor (_29506_, _29505_, _29502_);
  nor (_29507_, _29506_, _29481_);
  not (_29508_, _29507_);
  nor (_29509_, _29508_, _29376_);
  nand (_29510_, _29508_, _29376_);
  not (_29511_, _29510_);
  nor (_29512_, _29499_, _29413_);
  nor (_29513_, _29512_, _29503_);
  nor (_29514_, _29513_, _29502_);
  nor (_29515_, _29480_, _29398_);
  nor (_29517_, _29515_, _29514_);
  not (_29518_, _29517_);
  nor (_29519_, _29518_, _29391_);
  not (_29520_, _29519_);
  nor (_29521_, _29520_, _29511_);
  nor (_29522_, _29521_, _29509_);
  not (_29523_, _29509_);
  nand (_29524_, _29510_, _29523_);
  nor (_29525_, _29517_, _29394_);
  nor (_29526_, _29525_, _29519_);
  not (_29527_, _29526_);
  nor (_29528_, _29527_, _29524_);
  nor (_29529_, _29427_, _29425_);
  nor (_29530_, _29529_, _29497_);
  nand (_29531_, _29529_, _29497_);
  not (_29532_, _29531_);
  nor (_29533_, _29532_, _29530_);
  nor (_29534_, _29533_, _29502_);
  nor (_29535_, _29480_, _29419_);
  nor (_29536_, _29535_, _29534_);
  not (_29537_, _29536_);
  nor (_29538_, _29537_, _29403_);
  not (_29539_, _29538_);
  nor (_29540_, _29536_, _29411_);
  not (_29541_, _29540_);
  nor (_29542_, _29495_, _29494_);
  nor (_29543_, _29542_, _29471_);
  nor (_29544_, _29543_, _29502_);
  nor (_29545_, _29480_, _29431_);
  nor (_29546_, _29545_, _29544_);
  not (_29547_, _29546_);
  nor (_29548_, _29547_, _29424_);
  nand (_29549_, _29548_, _29541_);
  nand (_29550_, _29549_, _29539_);
  nand (_29551_, _29550_, _29528_);
  nand (_29552_, _29551_, _29522_);
  nor (_29553_, _29492_, _29483_);
  nor (_29554_, _29553_, _29466_);
  nor (_29555_, _29554_, _29502_);
  nor (_29556_, _29480_, _29442_);
  nor (_29558_, _29556_, _29555_);
  nand (_29559_, _29558_, _29428_);
  nor (_29560_, _29490_, _29488_);
  nor (_29561_, _29560_, _29464_);
  not (_29562_, _29561_);
  nand (_29563_, _29562_, _29480_);
  nand (_29564_, _29502_, _29451_);
  nand (_29565_, _29564_, _29563_);
  nor (_29566_, _29565_, _29436_);
  nor (_29567_, _29558_, _29428_);
  not (_29568_, _29428_);
  not (_29569_, _29554_);
  nand (_29570_, _29569_, _29480_);
  nand (_29571_, _29502_, _29440_);
  nand (_29572_, _29571_, _29570_);
  nor (_29573_, _29572_, _29568_);
  nor (_29574_, _29573_, _29567_);
  nand (_29575_, _29574_, _29566_);
  nand (_29576_, _29575_, _29559_);
  nor (_29577_, _29480_, _29487_);
  nor (_29578_, _29456_, _29484_);
  nor (_29579_, _29487_, _29453_);
  nor (_29580_, _29579_, _29578_);
  not (_29581_, _29580_);
  nor (_29582_, _29502_, _29581_);
  nor (_29583_, _29582_, _29577_);
  nor (_29584_, _29583_, _29447_);
  nand (_29585_, _29502_, _29456_);
  nand (_29586_, _29480_, _29580_);
  nand (_29587_, _29586_, _29585_);
  nand (_29588_, _29587_, _29458_);
  nand (_29589_, _29583_, _29447_);
  nand (_29590_, _29589_, _29588_);
  nor (_29591_, _29378_, _27861_);
  nor (_29592_, _29377_, _02212_);
  nor (_29593_, _29592_, _29591_);
  nor (_29594_, _29593_, _29453_);
  nor (_29595_, _29594_, _29590_);
  nor (_29596_, _29595_, _29584_);
  nor (_29597_, _29561_, _29502_);
  nor (_29599_, _29480_, _29460_);
  nor (_29600_, _29599_, _29597_);
  nor (_29601_, _29600_, _29435_);
  nor (_29602_, _29601_, _29566_);
  nand (_29603_, _29574_, _29602_);
  nor (_29604_, _29603_, _29596_);
  nor (_29605_, _29604_, _29576_);
  nor (_29606_, _29540_, _29538_);
  nor (_29607_, _29546_, _29426_);
  nor (_29608_, _29607_, _29548_);
  nand (_29609_, _29608_, _29606_);
  not (_29610_, _29609_);
  nand (_29611_, _29610_, _29528_);
  nor (_29612_, _29611_, _29605_);
  nor (_29613_, _29612_, _29552_);
  nor (_29614_, _29613_, _29370_);
  not (_29615_, _29550_);
  nand (_29616_, _29600_, _29435_);
  nand (_29617_, _29572_, _29568_);
  nand (_29618_, _29559_, _29617_);
  nor (_29619_, _29618_, _29616_);
  nor (_29620_, _29619_, _29573_);
  nor (_29621_, _29587_, _29458_);
  nor (_29622_, _29621_, _29584_);
  not (_29623_, _29594_);
  nand (_29624_, _29623_, _29622_);
  nand (_29625_, _29624_, _29588_);
  nand (_29626_, _29565_, _29436_);
  nand (_29627_, _29626_, _29616_);
  nor (_29628_, _29618_, _29627_);
  nand (_29629_, _29628_, _29625_);
  nand (_29630_, _29629_, _29620_);
  nand (_29631_, _29610_, _29630_);
  nand (_29632_, _29631_, _29615_);
  nand (_29633_, _29632_, _29526_);
  nor (_29634_, _29609_, _29605_);
  nor (_29635_, _29634_, _29550_);
  nand (_29636_, _29635_, _29527_);
  nand (_29637_, _29636_, _29633_);
  nand (_29638_, _29637_, _29614_);
  not (_29641_, _29522_);
  nor (_29642_, _29511_, _29509_);
  nand (_29643_, _29526_, _29642_);
  nor (_29644_, _29615_, _29643_);
  nor (_29645_, _29644_, _29641_);
  nor (_29646_, _29609_, _29643_);
  nand (_29647_, _29646_, _29630_);
  nand (_29648_, _29647_, _29645_);
  nand (_29649_, _29648_, _29369_);
  nand (_29650_, _29649_, _29518_);
  nand (_29651_, _29650_, _29638_);
  nor (_29652_, _29651_, _29346_);
  nor (_29653_, _27562_, _27522_);
  nor (_29654_, _01904_, _01866_);
  not (_29655_, _29654_);
  nand (_29656_, _29655_, _02008_);
  nand (_29657_, _29655_, _01995_);
  not (_29658_, _29657_);
  nand (_29659_, _29654_, _28611_);
  not (_29660_, _29659_);
  not (_29661_, _01904_);
  nor (_29662_, _29661_, _01866_);
  nand (_29663_, _29662_, _27040_);
  not (_29664_, _01866_);
  nor (_29665_, _01904_, _29664_);
  nand (_29666_, _29665_, _28500_);
  nand (_29667_, _29666_, _29663_);
  nor (_29668_, _29665_, _29662_);
  not (_29669_, _29668_);
  nor (_29670_, _29385_, _29664_);
  nor (_29671_, _29670_, _29669_);
  nor (_29672_, _29671_, _29667_);
  nor (_29673_, _29672_, _29660_);
  nand (_29674_, _29673_, _28454_);
  not (_29675_, _29674_);
  nand (_29676_, _29654_, _28327_);
  not (_29677_, _29662_);
  nor (_29678_, _29677_, _28578_);
  not (_29679_, _29665_);
  nor (_29680_, _29679_, _27671_);
  nor (_29682_, _29680_, _29678_);
  nand (_29683_, _28123_, _01866_);
  nand (_29684_, _29683_, _29668_);
  nand (_29685_, _29684_, _29682_);
  nand (_29686_, _29685_, _29676_);
  nor (_29687_, _29686_, _28313_);
  not (_29688_, _29687_);
  nor (_29689_, _29688_, _29675_);
  not (_29690_, _29689_);
  nor (_29691_, _29677_, _27081_);
  nor (_29692_, _29679_, _28521_);
  nor (_29693_, _29692_, _29691_);
  nand (_29694_, _27849_, _01866_);
  nand (_29695_, _29694_, _29668_);
  nand (_29696_, _29695_, _29693_);
  nand (_29697_, _29696_, _29659_);
  nor (_29698_, _29697_, _27016_);
  nor (_29699_, _29686_, _28391_);
  nand (_29700_, _29699_, _29698_);
  nand (_29701_, _29700_, _29674_);
  not (_29702_, _29676_);
  nand (_29703_, _29662_, _28570_);
  nand (_29704_, _29665_, _27645_);
  nand (_29705_, _29704_, _29703_);
  nor (_29706_, _28096_, _29664_);
  nor (_29707_, _29706_, _29669_);
  nor (_29708_, _29707_, _29705_);
  nor (_29709_, _29708_, _29702_);
  nand (_29710_, _29709_, _28393_);
  nor (_29711_, _29700_, _28452_);
  nor (_29712_, _29711_, _29710_);
  nand (_29713_, _29712_, _29701_);
  nor (_29714_, _29688_, _29674_);
  nor (_29715_, _29697_, _28313_);
  nor (_29716_, _29686_, _28452_);
  nor (_29717_, _29716_, _29715_);
  nor (_29718_, _29717_, _29714_);
  not (_29719_, _29718_);
  nor (_29720_, _29719_, _29713_);
  nand (_29721_, _29673_, _27018_);
  nor (_29723_, _29710_, _29721_);
  nand (_29724_, _29723_, _28454_);
  nor (_29725_, _29719_, _29724_);
  nor (_29726_, _29725_, _29720_);
  nor (_29727_, _29726_, _29690_);
  nand (_29728_, _29726_, _29690_);
  not (_29729_, _29728_);
  nor (_29730_, _29729_, _29727_);
  nor (_29731_, _29686_, _27016_);
  not (_29732_, _29731_);
  nor (_29733_, _29697_, _27403_);
  not (_29734_, _29733_);
  nor (_29735_, _29734_, _29732_);
  nor (_29736_, _29697_, _28391_);
  nor (_29737_, _29736_, _29731_);
  nor (_29738_, _29737_, _29723_);
  nand (_29739_, _29738_, _29735_);
  nor (_29740_, _29699_, _29675_);
  not (_29741_, _29740_);
  nand (_29742_, _29741_, _29713_);
  nor (_29743_, _29742_, _29739_);
  nand (_29744_, _29724_, _29701_);
  nor (_29745_, _29744_, _29710_);
  nor (_29746_, _29718_, _29745_);
  nor (_29747_, _29746_, _29720_);
  nor (_29748_, _29747_, _29711_);
  nor (_29749_, _29748_, _29725_);
  nand (_29750_, _29749_, _29743_);
  not (_29751_, _29739_);
  nor (_29752_, _29740_, _29745_);
  nand (_29753_, _29752_, _29751_);
  not (_29754_, _29725_);
  nand (_29755_, _29718_, _29745_);
  nand (_29756_, _29719_, _29713_);
  nand (_29757_, _29756_, _29755_);
  nand (_29758_, _29757_, _29724_);
  nand (_29759_, _29758_, _29754_);
  nor (_29760_, _29759_, _29753_);
  nor (_29761_, _29749_, _29743_);
  nor (_29762_, _29761_, _29760_);
  nor (_29764_, _29686_, _27476_);
  nor (_29765_, _29697_, _28510_);
  nand (_29766_, _29765_, _29764_);
  nor (_29767_, _29697_, _27476_);
  nor (_29768_, _29686_, _28510_);
  not (_29769_, _29768_);
  nor (_29770_, _29769_, _29767_);
  nand (_29771_, _29770_, _29733_);
  nand (_29772_, _29771_, _29766_);
  nor (_29773_, _29686_, _27403_);
  nor (_29774_, _29773_, _29698_);
  nor (_29775_, _29774_, _29735_);
  nand (_29776_, _29775_, _29772_);
  nor (_29777_, _29738_, _29735_);
  not (_29778_, _29777_);
  nand (_29779_, _29778_, _29739_);
  nor (_29780_, _29779_, _29776_);
  nor (_29781_, _29752_, _29751_);
  nor (_29782_, _29781_, _29743_);
  nand (_29783_, _29782_, _29780_);
  not (_29784_, _29764_);
  nor (_29785_, _29697_, _27271_);
  not (_29786_, _29785_);
  nor (_29787_, _29786_, _29784_);
  not (_29788_, _29766_);
  nor (_29789_, _29765_, _29764_);
  nor (_29790_, _29789_, _29788_);
  nand (_29791_, _29790_, _29787_);
  not (_29792_, _29767_);
  nand (_29793_, _29768_, _29792_);
  nand (_29794_, _29793_, _29734_);
  nand (_29795_, _29794_, _29771_);
  nor (_29796_, _29795_, _29791_);
  nor (_29797_, _29793_, _29734_);
  nor (_29798_, _29797_, _29788_);
  not (_29799_, _29775_);
  nor (_29800_, _29799_, _29798_);
  nor (_29801_, _29775_, _29772_);
  nor (_29802_, _29801_, _29800_);
  nand (_29803_, _29802_, _29796_);
  nor (_29805_, _29777_, _29751_);
  nand (_29806_, _29805_, _29800_);
  nand (_29807_, _29779_, _29776_);
  nand (_29808_, _29807_, _29806_);
  nor (_29809_, _29808_, _29803_);
  nand (_29810_, _29742_, _29739_);
  nand (_29811_, _29810_, _29753_);
  nor (_29812_, _29811_, _29806_);
  nor (_29813_, _29782_, _29780_);
  nor (_29814_, _29813_, _29812_);
  nand (_29815_, _29814_, _29809_);
  nand (_29816_, _29815_, _29783_);
  nand (_29817_, _29816_, _29762_);
  nand (_29818_, _29817_, _29750_);
  nand (_29819_, _29818_, _29730_);
  nor (_29820_, _29727_, _29714_);
  nand (_29821_, _29820_, _29819_);
  nand (_29822_, _29821_, _29658_);
  not (_29823_, _29730_);
  nand (_29824_, _29759_, _29753_);
  nand (_29825_, _29824_, _29750_);
  not (_29826_, _29787_);
  not (_29827_, _29789_);
  nand (_29828_, _29827_, _29766_);
  nor (_29829_, _29828_, _29826_);
  nor (_29830_, _29770_, _29733_);
  nor (_29831_, _29830_, _29797_);
  nand (_29832_, _29831_, _29829_);
  nand (_29833_, _29799_, _29798_);
  nand (_29834_, _29833_, _29776_);
  nor (_29835_, _29834_, _29832_);
  nor (_29836_, _29805_, _29800_);
  nor (_29837_, _29836_, _29780_);
  nand (_29838_, _29837_, _29835_);
  nand (_29839_, _29811_, _29806_);
  nand (_29840_, _29839_, _29783_);
  nor (_29841_, _29840_, _29838_);
  nor (_29842_, _29841_, _29812_);
  nor (_29843_, _29842_, _29825_);
  nor (_29844_, _29843_, _29760_);
  nor (_29846_, _29844_, _29823_);
  not (_29847_, _29820_);
  nor (_29848_, _29847_, _29846_);
  nand (_29849_, _29848_, _29657_);
  nand (_29850_, _29655_, _01993_);
  nand (_29851_, _29844_, _29823_);
  nand (_29852_, _29851_, _29819_);
  nor (_29853_, _29852_, _29850_);
  nand (_29854_, _29853_, _29849_);
  nand (_29855_, _29854_, _29822_);
  nand (_29856_, _29655_, _01998_);
  nand (_29857_, _29655_, _02000_);
  nor (_29858_, _29857_, _29856_);
  nand (_29859_, _29858_, _29855_);
  nand (_29860_, _29655_, _01991_);
  not (_29861_, _29860_);
  nor (_29862_, _29816_, _29762_);
  nor (_29863_, _29862_, _29843_);
  nand (_29864_, _29863_, _29861_);
  not (_29865_, _29864_);
  nor (_29866_, _29863_, _29861_);
  nor (_29867_, _29866_, _29865_);
  nand (_29868_, _29655_, _01988_);
  not (_29869_, _29868_);
  nor (_29870_, _29814_, _29809_);
  nor (_29871_, _29870_, _29841_);
  nand (_29872_, _29871_, _29869_);
  not (_29873_, _29872_);
  nor (_29874_, _29871_, _29869_);
  nor (_29875_, _29874_, _29873_);
  nand (_29876_, _29655_, _01985_);
  not (_29877_, _29876_);
  nor (_29878_, _29837_, _29835_);
  nor (_29879_, _29878_, _29809_);
  nand (_29880_, _29879_, _29877_);
  not (_29881_, _29880_);
  nor (_29882_, _29879_, _29877_);
  nor (_29883_, _29882_, _29881_);
  nand (_29884_, _29655_, _01983_);
  not (_29885_, _29884_);
  nor (_29887_, _29802_, _29796_);
  nor (_29888_, _29887_, _29835_);
  nand (_29889_, _29888_, _29885_);
  nand (_29890_, _29655_, _01981_);
  not (_29891_, _29890_);
  nor (_29892_, _29831_, _29829_);
  nor (_29893_, _29892_, _29796_);
  nand (_29894_, _29893_, _29891_);
  nand (_29895_, _29655_, _01977_);
  not (_29896_, _29895_);
  nor (_29897_, _29790_, _29787_);
  nor (_29898_, _29897_, _29829_);
  nand (_29899_, _29898_, _29896_);
  not (_29900_, _29899_);
  nand (_29901_, _29795_, _29791_);
  nand (_29902_, _29901_, _29832_);
  nor (_29903_, _29902_, _29890_);
  nor (_29904_, _29893_, _29891_);
  nor (_29905_, _29904_, _29903_);
  nand (_29906_, _29905_, _29900_);
  nand (_29907_, _29906_, _29894_);
  nand (_29908_, _29834_, _29832_);
  nand (_29909_, _29908_, _29803_);
  nor (_29910_, _29909_, _29884_);
  nor (_29911_, _29888_, _29885_);
  nor (_29912_, _29911_, _29910_);
  nand (_29913_, _29912_, _29907_);
  nand (_29914_, _29913_, _29889_);
  nand (_29915_, _29914_, _29883_);
  nand (_29916_, _29915_, _29880_);
  nand (_29917_, _29916_, _29875_);
  nand (_29918_, _29917_, _29872_);
  nand (_29919_, _29918_, _29867_);
  nand (_29920_, _29919_, _29864_);
  not (_29921_, _29850_);
  nor (_29922_, _29818_, _29730_);
  nor (_29923_, _29922_, _29846_);
  nor (_29924_, _29923_, _29921_);
  nor (_29925_, _29924_, _29853_);
  nor (_29926_, _29821_, _29658_);
  nor (_29928_, _29848_, _29657_);
  nor (_29929_, _29928_, _29926_);
  nand (_29930_, _29929_, _29925_);
  not (_29931_, _29858_);
  nor (_29932_, _29931_, _29930_);
  nand (_29933_, _29932_, _29920_);
  nand (_29934_, _29933_, _29859_);
  nand (_29935_, _29655_, _02002_);
  nand (_29936_, _29655_, _02005_);
  nor (_29937_, _29936_, _29935_);
  nand (_29938_, _29937_, _29934_);
  nor (_29939_, _29938_, _29656_);
  not (_29940_, _29656_);
  nand (_29941_, _29923_, _29921_);
  nor (_29942_, _29941_, _29926_);
  nor (_29943_, _29942_, _29928_);
  nor (_29944_, _29931_, _29943_);
  not (_29945_, _29866_);
  nand (_29946_, _29945_, _29864_);
  not (_29947_, _29874_);
  nand (_29948_, _29947_, _29872_);
  not (_29949_, _29882_);
  nand (_29950_, _29949_, _29880_);
  nand (_29951_, _29902_, _29890_);
  nand (_29952_, _29951_, _29894_);
  nor (_29953_, _29952_, _29899_);
  nor (_29954_, _29953_, _29903_);
  nand (_29955_, _29909_, _29884_);
  nand (_29956_, _29955_, _29889_);
  nor (_29957_, _29956_, _29954_);
  nor (_29958_, _29957_, _29910_);
  nor (_29959_, _29958_, _29950_);
  nor (_29960_, _29959_, _29881_);
  nor (_29961_, _29960_, _29948_);
  nor (_29962_, _29961_, _29873_);
  nor (_29963_, _29962_, _29946_);
  nor (_29964_, _29963_, _29865_);
  nand (_29965_, _29852_, _29850_);
  nand (_29966_, _29965_, _29941_);
  nand (_29967_, _29822_, _29849_);
  nor (_29969_, _29967_, _29966_);
  nand (_29970_, _29858_, _29969_);
  nor (_29971_, _29970_, _29964_);
  nor (_29972_, _29971_, _29944_);
  not (_29973_, _29937_);
  nor (_29974_, _29973_, _29972_);
  nor (_29975_, _29974_, _29940_);
  nor (_29976_, _29975_, _29939_);
  nand (_29977_, _29976_, _29653_);
  nor (_29978_, _28129_, _27853_);
  nor (_29979_, _29978_, _28125_);
  nor (_29980_, _29979_, _28524_);
  nor (_29981_, _29980_, _28522_);
  nor (_29982_, _29981_, _27675_);
  nand (_29983_, _29981_, _27675_);
  not (_29984_, _29983_);
  nor (_29985_, _29984_, _29982_);
  nor (_29986_, _27870_, _27466_);
  not (_29987_, _29986_);
  nor (_29988_, _29987_, _28129_);
  nand (_29989_, _29979_, _28524_);
  not (_29990_, _29989_);
  nor (_29991_, _29990_, _29980_);
  nand (_29992_, _29991_, _29988_);
  nor (_29993_, _29992_, _29985_);
  nor (_29994_, _29981_, _27647_);
  nor (_29995_, _29994_, _27673_);
  not (_29996_, _29995_);
  nor (_29997_, _29996_, _29993_);
  nor (_29998_, _29997_, _27087_);
  nand (_29999_, _29998_, _28580_);
  not (_30000_, _29999_);
  nor (_30001_, _28581_, _27550_);
  nor (_30002_, _30001_, _28579_);
  nor (_30003_, _30002_, _28616_);
  not (_30004_, _30003_);
  nand (_30005_, _30002_, _28616_);
  nand (_30006_, _30005_, _30004_);
  not (_30007_, _30006_);
  nor (_30008_, _30007_, _30000_);
  nor (_30010_, _27562_, _26923_);
  not (_30011_, _30010_);
  nor (_30012_, _30006_, _29999_);
  nor (_30013_, _30012_, _30011_);
  not (_30014_, _30013_);
  nor (_30015_, _30014_, _30008_);
  not (_30016_, _27564_);
  nor (_30017_, _27081_, _27018_);
  nor (_30018_, _28580_, _30017_);
  not (_30019_, _30018_);
  nand (_30020_, _28580_, _30017_);
  nand (_30021_, _30020_, _30019_);
  not (_30022_, _30021_);
  nor (_30023_, _28500_, _28510_);
  nor (_30024_, _28096_, _27476_);
  nor (_30025_, _27849_, _27861_);
  nor (_30026_, _28127_, _30025_);
  nor (_30027_, _30026_, _30024_);
  nor (_30028_, _30027_, _28523_);
  nor (_30029_, _30028_, _30023_);
  nor (_30030_, _30029_, _27675_);
  not (_30031_, _30029_);
  nor (_30032_, _30031_, _27677_);
  nor (_30033_, _30032_, _30030_);
  nand (_30034_, _30027_, _28523_);
  not (_30035_, _30034_);
  nor (_30036_, _30035_, _30028_);
  nand (_30037_, _28127_, _30025_);
  not (_30038_, _30037_);
  nor (_30039_, _30038_, _30026_);
  not (_30040_, _27870_);
  nor (_30041_, _30040_, _27466_);
  not (_30042_, _30041_);
  nor (_30043_, _30042_, _30039_);
  not (_30044_, _30043_);
  nor (_30045_, _30044_, _30036_);
  not (_30046_, _30045_);
  nor (_30047_, _30046_, _30033_);
  nor (_30048_, _27645_, _27403_);
  nor (_30049_, _27671_, _27405_);
  nor (_30052_, _30029_, _30049_);
  nor (_30053_, _30052_, _30048_);
  nor (_30054_, _30053_, _30047_);
  nor (_30055_, _30054_, _27085_);
  not (_30056_, _30055_);
  nor (_30057_, _30056_, _30022_);
  nor (_30058_, _28570_, _28391_);
  nor (_30059_, _30018_, _30058_);
  nor (_30060_, _30059_, _28615_);
  not (_30061_, _30060_);
  nand (_30062_, _30059_, _28615_);
  nand (_30063_, _30062_, _30061_);
  nor (_30064_, _30063_, _30057_);
  nand (_30065_, _30063_, _30057_);
  not (_30066_, _30065_);
  nor (_30067_, _30066_, _30064_);
  nor (_30068_, _30067_, _30016_);
  nor (_30069_, _27544_, _26923_);
  nor (_30070_, _28454_, _28393_);
  nor (_30071_, _30070_, _28313_);
  not (_30072_, _30069_);
  nor (_30073_, _27403_, _27360_);
  not (_30074_, _30073_);
  nor (_30075_, _30074_, _30072_);
  nor (_30076_, _30075_, _30071_);
  nand (_30077_, _30076_, _27466_);
  not (_30078_, _30077_);
  not (_30079_, _30075_);
  nor (_30080_, _30079_, _27016_);
  nor (_30081_, _30080_, _28393_);
  nor (_30082_, _30081_, _30078_);
  nand (_30083_, _30082_, _28454_);
  not (_30084_, _30070_);
  nor (_30085_, _30080_, _30084_);
  not (_30086_, _30085_);
  nor (_30087_, _30086_, _30078_);
  not (_30088_, _30080_);
  nor (_30089_, _30088_, _28391_);
  nor (_30090_, _30089_, _28454_);
  nor (_30091_, _30090_, _30077_);
  nor (_30093_, _30091_, _30087_);
  nand (_30094_, _30093_, _30083_);
  nand (_30095_, _30094_, _30069_);
  nor (_30096_, _30010_, _27564_);
  not (_30097_, _30096_);
  nor (_30098_, _27546_, _26907_);
  nor (_30099_, _27544_, _27520_);
  nor (_30100_, _30099_, _29653_);
  nand (_30101_, _30100_, _30098_);
  nor (_30102_, _30101_, _30097_);
  not (_30103_, _30102_);
  nor (_30104_, _30103_, _28452_);
  nor (_30105_, _27504_, _03811_);
  not (_30106_, _30105_);
  nor (_30107_, _30106_, _28313_);
  nor (_30108_, _30107_, _30104_);
  nor (_30109_, _26913_, _27046_);
  not (_30110_, _30109_);
  nor (_30111_, _30110_, _28391_);
  nor (_30112_, _30111_, _28636_);
  nand (_30113_, _30112_, _30108_);
  nor (_30114_, _30113_, _28633_);
  nand (_30115_, _30114_, _30095_);
  nor (_30116_, _30115_, _28631_);
  not (_30117_, _30116_);
  nor (_30118_, _30117_, _30068_);
  not (_30119_, _30118_);
  nor (_30120_, _30119_, _30015_);
  nand (_30121_, _30120_, _29977_);
  nor (_30122_, _30121_, _29652_);
  nand (_30123_, _30122_, _29041_);
  nand (_30124_, _30123_, _29344_);
  nor (_29226_, _30124_, _29343_);
  nand (_30125_, _29063_, _01432_);
  nand (_30126_, _29048_, _01456_);
  nand (_30127_, _30126_, _30125_);
  nand (_30128_, _29070_, _00841_);
  nand (_30129_, _29074_, _01389_);
  nand (_30130_, _30129_, _30128_);
  nor (_30131_, _30130_, _30127_);
  nand (_30133_, _29082_, _01485_);
  nand (_30134_, _29084_, _00343_);
  nand (_30135_, _30134_, _30133_);
  nand (_30136_, _29094_, _00207_);
  nand (_30137_, _29104_, _00204_);
  nand (_30138_, _30137_, _30136_);
  nor (_30139_, _30138_, _30135_);
  nand (_30140_, _30139_, _30131_);
  nand (_30141_, _29111_, _31271_);
  nand (_30142_, _29109_, _31251_);
  nand (_30143_, _30142_, _30141_);
  nand (_30144_, _29114_, _31029_);
  nand (_30145_, _29118_, _00018_);
  nand (_30146_, _30145_, _30144_);
  nor (_30147_, _30146_, _30143_);
  nand (_30148_, _29126_, _01032_);
  nand (_30149_, _29128_, _00762_);
  nand (_30150_, _30149_, _30148_);
  nand (_30151_, _29134_, _31064_);
  nand (_30152_, _29132_, _01195_);
  nand (_30153_, _30152_, _30151_);
  nor (_30154_, _30153_, _30150_);
  nand (_30155_, _30154_, _30147_);
  nor (_30156_, _30155_, _30140_);
  nand (_30157_, _29156_, _30780_);
  nand (_30158_, _29035_, _30809_);
  nand (_30159_, _30158_, _30157_);
  nand (_30160_, _29149_, _01585_);
  not (_30161_, _28900_);
  nand (_30162_, _29153_, _30161_);
  nand (_30163_, _30162_, _30160_);
  nor (_30164_, _30163_, _30159_);
  nor (_30165_, _29208_, _30588_);
  nor (_30166_, _29210_, _30517_);
  nor (_30167_, _30166_, _30165_);
  nand (_30168_, _30167_, _29163_);
  nor (_30169_, _29208_, _30610_);
  nor (_30170_, _29210_, _30297_);
  nor (_30171_, _30170_, _30169_);
  nand (_30172_, _30171_, _29218_);
  nand (_30174_, _30172_, _30168_);
  nor (_30175_, _29208_, _30567_);
  nor (_30176_, _29210_, _30512_);
  nor (_30177_, _30176_, _30175_);
  nand (_30178_, _30177_, _29224_);
  nor (_30179_, _29208_, _30546_);
  nor (_30180_, _29210_, _30392_);
  nor (_30181_, _30180_, _30179_);
  nand (_30182_, _30181_, _29232_);
  nand (_30183_, _30182_, _30178_);
  nor (_30184_, _30183_, _30174_);
  nand (_30185_, _30184_, _30164_);
  nand (_30186_, _29146_, _01703_);
  nand (_30187_, _29143_, _30705_);
  nand (_30188_, _30187_, _30186_);
  nor (_30189_, _30188_, _30185_);
  nand (_30190_, _30189_, _30156_);
  nand (_30191_, _30190_, _29305_);
  nand (_30192_, _29340_, _06128_);
  nand (_30193_, _30192_, _30191_);
  nor (_30194_, _30193_, _29041_);
  not (_30195_, _29653_);
  not (_30196_, _29935_);
  nand (_30197_, _30196_, _29934_);
  nand (_30198_, _29936_, _30197_);
  nand (_30199_, _30198_, _29938_);
  nor (_30200_, _30199_, _30195_);
  nand (_30201_, _29649_, _29536_);
  not (_30202_, _29608_);
  nor (_30203_, _30202_, _29605_);
  nor (_30204_, _30203_, _29548_);
  nand (_30205_, _30204_, _29606_);
  not (_30206_, _29606_);
  not (_30207_, _29548_);
  nand (_30208_, _29608_, _29630_);
  nand (_30209_, _30208_, _30207_);
  nand (_30210_, _30209_, _30206_);
  nand (_30211_, _30210_, _30205_);
  nand (_30212_, _30211_, _29614_);
  nand (_30213_, _30212_, _30201_);
  nand (_30215_, _30213_, _29345_);
  nor (_30216_, _30055_, _30021_);
  nor (_30217_, _30216_, _30057_);
  nor (_30218_, _30217_, _30016_);
  nor (_30219_, _28580_, _27083_);
  nor (_30220_, _30219_, _30001_);
  nor (_30221_, _30220_, _29998_);
  not (_30222_, _30221_);
  nand (_30223_, _30222_, _30010_);
  nor (_30224_, _30223_, _30000_);
  not (_30225_, _30089_);
  nand (_30226_, _30082_, _30225_);
  nor (_30227_, _30077_, _28393_);
  nor (_30228_, _30227_, _30072_);
  nand (_30229_, _30228_, _30226_);
  nor (_30230_, _30110_, _27016_);
  nor (_30231_, _30230_, _28595_);
  nor (_30232_, _30103_, _28391_);
  nor (_30233_, _30106_, _28452_);
  nor (_30234_, _30233_, _30232_);
  nand (_30235_, _30234_, _30231_);
  nor (_30236_, _30235_, _28592_);
  nand (_30237_, _30236_, _30229_);
  nor (_30238_, _30237_, _28590_);
  not (_30239_, _30238_);
  nor (_30240_, _30239_, _30224_);
  not (_30241_, _30240_);
  nor (_30242_, _30241_, _30218_);
  nand (_30243_, _30242_, _30215_);
  nor (_30244_, _30243_, _30200_);
  nand (_30245_, _30244_, _29041_);
  nand (_30246_, _30245_, _29344_);
  nor (_02158_, _30246_, _30194_);
  nand (_30247_, _29143_, _30655_);
  not (_30248_, _01710_);
  nor (_30249_, _29286_, _30248_);
  nor (_30250_, _29308_, _29123_);
  nor (_30251_, _29208_, _30564_);
  nor (_30252_, _29210_, _30490_);
  nor (_30253_, _30252_, _30251_);
  nand (_30255_, _30253_, _30250_);
  nor (_30256_, _28905_, _28781_);
  nand (_30257_, _29307_, _30256_);
  not (_30258_, _30257_);
  nor (_30259_, _29208_, _30543_);
  nor (_30260_, _29210_, _30374_);
  nor (_30261_, _30260_, _30259_);
  nand (_30262_, _30261_, _30258_);
  nand (_30263_, _30262_, _30255_);
  nor (_30264_, _30263_, _30249_);
  nand (_30265_, _30264_, _30247_);
  not (_30266_, _30806_);
  nor (_30267_, _29036_, _30266_);
  nand (_30268_, _29128_, _00784_);
  nand (_30269_, _29126_, _01029_);
  nand (_30270_, _30269_, _30268_);
  nor (_30271_, _30270_, _30267_);
  not (_30272_, _01627_);
  nor (_30273_, _29333_, _30272_);
  not (_30274_, _30777_);
  nor (_30275_, _29239_, _30274_);
  nor (_30276_, _30275_, _30273_);
  nand (_30278_, _30276_, _30271_);
  nor (_30280_, _30278_, _30265_);
  not (_30281_, _00022_);
  not (_30282_, _29118_);
  nor (_30284_, _30282_, _30281_);
  nand (_30286_, _29114_, _31031_);
  not (_30287_, _00256_);
  nor (_30289_, _29093_, _30287_);
  not (_30291_, _00230_);
  nor (_30292_, _29102_, _30291_);
  nor (_30293_, _30292_, _30289_);
  nand (_30294_, _30293_, _30286_);
  nor (_30295_, _30294_, _30284_);
  nand (_30296_, _29084_, _30975_);
  not (_30298_, _01453_);
  nor (_30299_, _29312_, _30298_);
  not (_30300_, _01291_);
  nor (_30302_, _29315_, _30300_);
  nor (_30304_, _30302_, _30299_);
  nand (_30305_, _30304_, _30296_);
  nand (_30306_, _29082_, _01482_);
  not (_30307_, _00888_);
  not (_30309_, _29070_);
  nor (_30310_, _30309_, _30307_);
  not (_30311_, _01374_);
  not (_30312_, _29074_);
  nor (_30314_, _30312_, _30311_);
  nor (_30315_, _30314_, _30310_);
  nand (_30317_, _30315_, _30306_);
  nor (_30318_, _30317_, _30305_);
  nand (_30319_, _30318_, _30295_);
  nor (_30320_, _29330_, _28775_);
  nor (_30322_, _29308_, _29100_);
  nor (_30323_, _29208_, _30607_);
  nor (_30324_, _29210_, _30471_);
  nor (_30326_, _30324_, _30323_);
  nand (_30327_, _30326_, _30322_);
  nor (_30328_, _29308_, _29091_);
  nor (_30329_, _29208_, _30585_);
  nor (_30330_, _29210_, _30483_);
  nor (_30332_, _30330_, _30329_);
  nand (_30333_, _30332_, _30328_);
  nand (_30334_, _30333_, _30327_);
  nor (_30335_, _30334_, _30320_);
  nand (_30336_, _29111_, _31022_);
  nand (_30337_, _29109_, _31135_);
  nand (_30338_, _30337_, _30336_);
  nand (_30340_, _29134_, _31066_);
  nand (_30341_, _29132_, _01193_);
  nand (_30342_, _30341_, _30340_);
  nor (_30343_, _30342_, _30338_);
  nand (_30344_, _30343_, _30335_);
  nor (_30345_, _30344_, _30319_);
  nand (_30347_, _30345_, _30280_);
  nand (_30348_, _30347_, _29305_);
  nand (_30349_, _29340_, _06125_);
  nand (_30350_, _30349_, _30348_);
  nor (_30351_, _30350_, _29041_);
  nand (_30353_, _30202_, _29605_);
  nand (_30354_, _30353_, _30208_);
  nand (_30355_, _30354_, _29614_);
  nand (_30356_, _29649_, _29547_);
  nand (_30357_, _30356_, _30355_);
  nor (_30359_, _30357_, _29346_);
  nor (_30360_, _29935_, _29972_);
  nor (_30361_, _30196_, _29934_);
  nor (_30362_, _30361_, _30360_);
  nand (_30363_, _30362_, _29653_);
  not (_30364_, _30054_);
  nor (_30365_, _30364_, _27085_);
  nor (_30366_, _30054_, _27087_);
  nor (_30367_, _30366_, _30365_);
  not (_30368_, _30367_);
  nor (_30369_, _30368_, _30016_);
  not (_30370_, _29997_);
  nor (_30371_, _30370_, _27085_);
  nor (_30372_, _30011_, _29998_);
  not (_30373_, _30372_);
  nor (_30375_, _30373_, _30371_);
  nor (_30376_, _30103_, _27016_);
  nor (_30377_, _30106_, _28391_);
  nor (_30378_, _30377_, _30376_);
  nor (_30380_, _30110_, _27403_);
  nor (_30381_, _30380_, _27578_);
  nand (_30382_, _30381_, _30378_);
  nor (_30383_, _30382_, _27552_);
  nor (_30384_, _30075_, _27018_);
  nor (_30385_, _30384_, _30080_);
  nand (_30386_, _30385_, _30069_);
  nand (_30387_, _30386_, _30383_);
  nor (_30388_, _30387_, _27538_);
  not (_30389_, _30388_);
  nor (_30390_, _30389_, _30375_);
  not (_30391_, _30390_);
  nor (_30393_, _30391_, _30369_);
  nand (_30394_, _30393_, _30363_);
  nor (_30395_, _30394_, _30359_);
  nand (_30397_, _30395_, _29041_);
  nand (_30399_, _30397_, _29344_);
  nor (_06159_, _30399_, _30351_);
  nand (_30400_, _29048_, _01450_);
  nand (_30401_, _29063_, _01405_);
  nand (_30403_, _30401_, _30400_);
  nand (_30404_, _29070_, _01224_);
  nand (_30405_, _29074_, _01415_);
  nand (_30406_, _30405_, _30404_);
  nor (_30407_, _30406_, _30403_);
  nand (_30408_, _29084_, _00512_);
  nand (_30410_, _29082_, _01479_);
  nand (_30411_, _30410_, _30408_);
  nand (_30412_, _29094_, _00224_);
  nand (_30413_, _29104_, _00246_);
  nand (_30414_, _30413_, _30412_);
  nor (_30415_, _30414_, _30411_);
  nand (_30416_, _30415_, _30407_);
  nand (_30417_, _29109_, _31246_);
  nand (_30418_, _29111_, _31158_);
  nand (_30419_, _30418_, _30417_);
  nand (_30420_, _29114_, _31232_);
  nand (_30421_, _29118_, _00162_);
  nand (_30422_, _30421_, _30420_);
  nor (_30423_, _30422_, _30419_);
  nand (_30425_, _29126_, _01025_);
  nand (_30426_, _29128_, _00941_);
  nand (_30427_, _30426_, _30425_);
  nand (_30429_, _29132_, _01191_);
  nand (_30430_, _29134_, _31176_);
  nand (_30431_, _30430_, _30429_);
  nor (_30432_, _30431_, _30427_);
  nand (_30433_, _30432_, _30423_);
  nor (_30434_, _30433_, _30416_);
  nand (_30435_, _29146_, _01714_);
  nand (_30436_, _29143_, _30691_);
  nand (_30437_, _30436_, _30435_);
  nand (_30438_, _29149_, _01620_);
  nand (_30439_, _29153_, _28914_);
  nand (_30441_, _30439_, _30438_);
  nand (_30442_, _29035_, _30803_);
  nand (_30444_, _29156_, _30773_);
  nand (_30445_, _30444_, _30442_);
  nor (_30446_, _30445_, _30441_);
  nor (_30447_, _29208_, _30582_);
  nor (_30448_, _29210_, _30456_);
  nor (_30449_, _30448_, _30447_);
  nand (_30450_, _30449_, _29163_);
  nor (_30452_, _29208_, _30604_);
  nor (_30453_, _29210_, _30396_);
  nor (_30454_, _30453_, _30452_);
  nand (_30455_, _30454_, _29218_);
  nand (_30457_, _30455_, _30450_);
  nor (_30458_, _29208_, _30561_);
  nor (_30460_, _29210_, _30478_);
  nor (_30461_, _30460_, _30458_);
  nand (_30462_, _30461_, _29224_);
  nor (_30463_, _29208_, _30540_);
  nor (_30464_, _29210_, _30358_);
  nor (_30465_, _30464_, _30463_);
  nand (_30467_, _30465_, _29232_);
  nand (_30468_, _30467_, _30462_);
  nor (_30469_, _30468_, _30457_);
  nand (_30470_, _30469_, _30446_);
  nor (_30472_, _30470_, _30437_);
  nand (_30473_, _30472_, _30434_);
  nand (_30474_, _30473_, _29305_);
  nand (_30475_, _29340_, _06122_);
  nand (_30476_, _30475_, _30474_);
  nor (_30477_, _30476_, _29041_);
  nor (_30479_, _29930_, _29964_);
  nor (_30480_, _30479_, _29855_);
  nor (_30481_, _30480_, _29856_);
  not (_30482_, _29857_);
  nor (_30484_, _30482_, _30481_);
  nor (_30485_, _30484_, _29934_);
  nand (_30486_, _30485_, _29653_);
  nand (_30487_, _30046_, _30033_);
  not (_30488_, _30487_);
  nor (_30489_, _30488_, _30047_);
  nor (_30491_, _30489_, _30016_);
  nor (_30494_, _30073_, _30072_);
  not (_30495_, _30494_);
  not (_30496_, _30666_);
  nor (_30498_, _27360_, _30496_);
  nor (_30499_, _30498_, _27405_);
  nor (_30500_, _30499_, _30495_);
  nor (_30501_, _30500_, _30491_);
  nand (_30502_, _30501_, _30486_);
  nand (_30503_, _29649_, _29558_);
  nor (_30504_, _29627_, _29596_);
  nor (_30505_, _30504_, _29566_);
  nand (_30506_, _30505_, _29574_);
  nor (_30507_, _30505_, _29574_);
  not (_30508_, _30507_);
  nand (_30509_, _30508_, _30506_);
  nand (_30510_, _30509_, _29614_);
  nand (_30511_, _30510_, _30503_);
  nand (_30513_, _30511_, _29345_);
  not (_30514_, _29985_);
  not (_30515_, _29992_);
  nor (_30516_, _30515_, _30514_);
  nor (_30518_, _30011_, _29993_);
  not (_30519_, _30518_);
  nor (_30520_, _30519_, _30516_);
  nor (_30521_, _30106_, _27016_);
  nor (_30522_, _30103_, _27403_);
  nor (_30523_, _30110_, _28510_);
  nor (_30524_, _30523_, _30522_);
  not (_30525_, _30524_);
  nor (_30526_, _30525_, _30521_);
  nand (_30527_, _30526_, _27714_);
  nor (_30528_, _30527_, _27736_);
  not (_30529_, _30528_);
  nor (_30530_, _30529_, _30520_);
  nand (_30532_, _30530_, _30513_);
  nor (_30533_, _30532_, _30502_);
  nand (_30535_, _30533_, _29041_);
  nand (_30536_, _30535_, _29344_);
  nor (_10626_, _30536_, _30477_);
  nand (_30538_, _29146_, _01718_);
  not (_30541_, _30677_);
  nor (_30542_, _29241_, _30541_);
  nor (_30544_, _29208_, _30558_);
  nor (_30545_, _29210_, _30466_);
  nor (_30547_, _30545_, _30544_);
  nand (_30548_, _30547_, _30250_);
  nor (_30550_, _29208_, _30537_);
  nor (_30551_, _29210_, _30339_);
  nor (_30553_, _30551_, _30550_);
  nand (_30554_, _30553_, _30258_);
  nand (_30556_, _30554_, _30548_);
  nor (_30557_, _30556_, _30542_);
  nand (_30559_, _30557_, _30538_);
  not (_30560_, _30769_);
  nor (_30562_, _29239_, _30560_);
  nand (_30563_, _29128_, _00929_);
  nand (_30565_, _29126_, _01022_);
  nand (_30566_, _30565_, _30563_);
  nor (_30568_, _30566_, _30562_);
  not (_30569_, _01606_);
  nor (_30571_, _29333_, _30569_);
  not (_30572_, _30800_);
  nor (_30574_, _29036_, _30572_);
  nor (_30575_, _30574_, _30571_);
  nand (_30577_, _30575_, _30568_);
  nor (_30578_, _30577_, _30559_);
  nand (_30580_, _29084_, _00315_);
  not (_30581_, _01447_);
  nor (_30583_, _29312_, _30581_);
  not (_30584_, _01409_);
  nor (_30586_, _29315_, _30584_);
  nor (_30587_, _30586_, _30583_);
  nand (_30589_, _30587_, _30580_);
  nand (_30590_, _29082_, _01476_);
  not (_30592_, _01238_);
  nor (_30593_, _30309_, _30592_);
  not (_30595_, _01383_);
  nor (_30596_, _30312_, _30595_);
  nor (_30598_, _30596_, _30593_);
  nand (_30599_, _30598_, _30590_);
  nor (_30602_, _30599_, _30589_);
  nand (_30603_, _29118_, _30961_);
  not (_30605_, _00236_);
  nor (_30606_, _29093_, _30605_);
  not (_30608_, _00495_);
  nor (_30609_, _29102_, _30608_);
  nor (_30611_, _30609_, _30606_);
  nand (_30612_, _30611_, _30603_);
  nand (_30614_, _29134_, _31178_);
  nand (_30615_, _29114_, _31144_);
  nand (_30616_, _30615_, _30614_);
  nor (_30617_, _30616_, _30612_);
  nand (_30618_, _30617_, _30602_);
  nor (_30619_, _29330_, _28978_);
  nor (_30620_, _29208_, _30601_);
  nor (_30621_, _29210_, _30331_);
  nor (_30622_, _30621_, _30620_);
  nand (_30623_, _30622_, _30322_);
  nor (_30624_, _29208_, _30579_);
  nor (_30625_, _29210_, _30428_);
  nor (_30626_, _30625_, _30624_);
  nand (_30627_, _30626_, _30328_);
  nand (_30628_, _30627_, _30623_);
  nor (_30629_, _30628_, _30619_);
  not (_30630_, _01189_);
  not (_30631_, _29132_);
  nor (_30632_, _30631_, _30630_);
  nand (_30633_, _29109_, _31243_);
  nand (_30634_, _29111_, _31285_);
  nand (_30635_, _30634_, _30633_);
  nor (_30636_, _30635_, _30632_);
  nand (_30637_, _30636_, _30629_);
  nor (_30638_, _30637_, _30618_);
  nand (_30639_, _30638_, _30578_);
  nand (_30640_, _30639_, _29305_);
  nand (_30641_, _29340_, _06119_);
  nand (_30642_, _30641_, _30640_);
  nor (_30643_, _30642_, _29041_);
  nor (_30644_, _29602_, _29625_);
  nor (_30645_, _30644_, _30504_);
  nor (_30647_, _30645_, _29649_);
  nor (_30648_, _29614_, _29600_);
  nor (_30649_, _30648_, _30647_);
  nand (_30650_, _30649_, _29345_);
  not (_30651_, _30481_);
  nand (_30652_, _30480_, _29856_);
  nand (_30653_, _30652_, _30651_);
  nor (_30654_, _30653_, _30195_);
  not (_30656_, _28531_);
  nor (_30657_, _29991_, _29988_);
  not (_30659_, _30657_);
  nand (_30660_, _30659_, _30010_);
  nor (_30661_, _30660_, _30515_);
  not (_30662_, _30036_);
  nor (_30663_, _30043_, _30662_);
  nor (_30664_, _30663_, _30045_);
  nor (_30665_, _30664_, _30016_);
  nand (_30667_, _27360_, _30666_);
  not (_30668_, _30667_);
  nor (_30669_, _30073_, _30666_);
  nor (_30671_, _30669_, _27318_);
  nor (_30672_, _30671_, _28510_);
  nor (_30673_, _30672_, _30668_);
  nor (_30674_, _30673_, _30072_);
  nor (_30675_, _30106_, _27403_);
  nor (_30676_, _30110_, _27476_);
  nor (_30678_, _30676_, _30675_);
  nor (_30679_, _30103_, _28510_);
  nor (_30680_, _30679_, _28537_);
  nand (_30681_, _30680_, _30678_);
  nor (_30682_, _30681_, _30674_);
  not (_30683_, _30682_);
  nor (_30684_, _30683_, _30665_);
  not (_30686_, _30684_);
  nor (_30687_, _30686_, _30661_);
  nand (_30688_, _30687_, _30656_);
  nor (_30690_, _30688_, _30654_);
  nand (_30692_, _30690_, _30650_);
  not (_30693_, _30692_);
  nand (_30694_, _30693_, _29041_);
  nand (_30696_, _30694_, _29344_);
  nor (_14540_, _30696_, _30643_);
  nand (_30697_, _29048_, _01444_);
  nand (_30698_, _29063_, _01412_);
  nand (_30699_, _30698_, _30697_);
  nand (_30700_, _29070_, _01229_);
  nand (_30701_, _29074_, _01421_);
  nand (_30703_, _30701_, _30700_);
  nor (_30704_, _30703_, _30699_);
  nand (_30706_, _29082_, _01473_);
  nand (_30707_, _29084_, _00517_);
  nand (_30708_, _30707_, _30706_);
  nand (_30709_, _29094_, _00250_);
  nand (_30710_, _29104_, _00435_);
  nand (_30711_, _30710_, _30709_);
  nor (_30712_, _30711_, _30708_);
  nand (_30713_, _30712_, _30704_);
  nand (_30714_, _29118_, _00155_);
  nand (_30715_, _29114_, _31208_);
  nand (_30716_, _30715_, _30714_);
  nand (_30717_, _29111_, _31275_);
  nand (_30718_, _29109_, _31202_);
  nand (_30719_, _30718_, _30717_);
  nor (_30720_, _30719_, _30716_);
  nand (_30721_, _29128_, _00920_);
  nand (_30722_, _29126_, _01018_);
  nand (_30723_, _30722_, _30721_);
  nand (_30724_, _29132_, _01187_);
  nand (_30725_, _29134_, _31216_);
  nand (_30726_, _30725_, _30724_);
  nor (_30727_, _30726_, _30723_);
  nand (_30728_, _30727_, _30720_);
  nor (_30729_, _30728_, _30713_);
  nand (_30730_, _29146_, _01722_);
  nand (_30731_, _29143_, _30670_);
  nand (_30732_, _30731_, _30730_);
  nand (_30733_, _29156_, _30765_);
  nand (_30734_, _29035_, _30797_);
  nand (_30735_, _30734_, _30733_);
  nand (_30737_, _29149_, _01597_);
  nand (_30739_, _29153_, _28187_);
  nand (_30740_, _30739_, _30737_);
  nor (_30741_, _30740_, _30735_);
  nor (_30742_, _29208_, _30576_);
  nor (_30744_, _29210_, _30402_);
  nor (_30745_, _30744_, _30742_);
  nand (_30746_, _30745_, _29163_);
  nor (_30747_, _29208_, _30597_);
  nor (_30748_, _29210_, _30497_);
  nor (_30749_, _30748_, _30747_);
  nand (_30750_, _30749_, _29218_);
  nand (_30751_, _30750_, _30746_);
  nor (_30752_, _29208_, _30555_);
  nor (_30753_, _29210_, _30451_);
  nor (_30754_, _30753_, _30752_);
  nand (_30755_, _30754_, _29224_);
  nor (_30756_, _29208_, _30534_);
  nor (_30757_, _29210_, _30325_);
  nor (_30758_, _30757_, _30756_);
  nand (_30759_, _30758_, _29232_);
  nand (_30760_, _30759_, _30755_);
  nor (_30762_, _30760_, _30751_);
  nand (_30763_, _30762_, _30741_);
  nor (_30764_, _30763_, _30732_);
  nand (_30766_, _30764_, _30729_);
  nand (_30767_, _30766_, _29305_);
  nand (_30768_, _29340_, _06117_);
  nand (_30770_, _30768_, _30767_);
  nor (_30771_, _30770_, _29041_);
  nor (_30772_, _29623_, _29622_);
  nor (_30774_, _30772_, _29595_);
  nor (_30775_, _30774_, _29649_);
  nor (_30776_, _29614_, _29587_);
  nor (_30778_, _30776_, _30775_);
  nand (_30779_, _30778_, _29345_);
  nor (_30781_, _29966_, _29964_);
  nor (_30782_, _30781_, _29853_);
  nor (_30784_, _30782_, _29929_);
  not (_30785_, _30782_);
  nor (_30786_, _30785_, _29967_);
  nor (_30788_, _30786_, _30784_);
  nor (_30789_, _30788_, _30195_);
  not (_30790_, _30039_);
  nor (_30791_, _30041_, _30790_);
  nor (_30792_, _30791_, _30043_);
  nor (_30793_, _30792_, _30016_);
  nor (_30795_, _28127_, _27851_);
  nor (_30796_, _30795_, _29978_);
  nor (_30798_, _30796_, _29986_);
  nor (_30799_, _30011_, _29988_);
  not (_30801_, _30799_);
  nor (_30802_, _30801_, _30798_);
  nor (_30804_, _30802_, _30793_);
  not (_30805_, _30804_);
  not (_30807_, _28141_);
  nand (_30808_, _30669_, _27318_);
  not (_30810_, _30808_);
  nor (_30811_, _30810_, _30671_);
  nor (_30813_, _30811_, _30072_);
  nor (_30814_, _30110_, _27271_);
  nor (_30815_, _30814_, _28151_);
  nor (_30816_, _30103_, _27476_);
  nor (_30817_, _30106_, _28510_);
  nor (_30818_, _30817_, _30816_);
  nand (_30819_, _30818_, _30815_);
  nor (_30820_, _30819_, _28145_);
  not (_30821_, _30820_);
  nor (_30823_, _30821_, _30813_);
  nand (_30824_, _30823_, _30807_);
  nor (_30825_, _30824_, _30805_);
  not (_30826_, _30825_);
  nor (_30827_, _30826_, _30789_);
  nand (_30828_, _30827_, _30779_);
  not (_30829_, _30828_);
  nand (_30830_, _30829_, _29041_);
  nand (_30831_, _30830_, _29344_);
  nor (_17402_, _30831_, _30771_);
  not (_30832_, _29593_);
  nor (_30833_, _29614_, _30832_);
  nor (_30834_, _29593_, _29484_);
  nor (_30836_, _30832_, _29453_);
  nor (_30837_, _30836_, _30834_);
  nand (_30838_, _29614_, _30837_);
  not (_30839_, _30838_);
  nor (_30840_, _30839_, _30833_);
  nor (_30841_, _30840_, _29346_);
  nor (_30842_, _29925_, _29920_);
  nor (_30843_, _30842_, _30781_);
  not (_30844_, _30843_);
  nor (_30845_, _30844_, _30195_);
  nor (_30846_, _30040_, _27225_);
  nor (_30847_, _30846_, _29986_);
  not (_30848_, _30847_);
  nor (_30849_, _30096_, _30848_);
  nor (_30850_, _27522_, _26913_);
  not (_30851_, _30850_);
  nor (_30852_, _30851_, _27466_);
  nor (_30853_, _30106_, _27476_);
  not (_30854_, _30853_);
  nor (_30856_, _26913_, _27494_);
  not (_30858_, _30856_);
  nor (_30859_, _30858_, _28313_);
  nor (_30860_, _30102_, _30069_);
  nor (_30861_, _30860_, _27271_);
  nor (_30862_, _30861_, _30859_);
  nand (_30863_, _30862_, _30854_);
  nor (_30864_, _30863_, _27855_);
  not (_30865_, _30864_);
  nor (_30866_, _30865_, _30852_);
  nand (_30867_, _30866_, _27884_);
  nor (_30869_, _30867_, _30849_);
  not (_30871_, _30869_);
  nor (_30872_, _30871_, _30845_);
  not (_30874_, _30872_);
  nor (_30876_, _30874_, _30841_);
  nand (_30877_, _30876_, _29041_);
  nand (_30879_, _30877_, _29344_);
  not (_30880_, _29305_);
  nor (_30881_, _26895_, _26777_);
  not (_30882_, _26751_);
  nor (_30884_, _26677_, _26640_);
  not (_30885_, _30884_);
  nor (_30886_, _30885_, _30882_);
  nand (_30887_, _30886_, _30881_);
  nor (_30888_, _30887_, _26789_);
  nor (_30889_, _30888_, _29290_);
  nor (_30890_, _30889_, _30395_);
  nor (_30891_, _28327_, _28315_);
  nor (_30892_, _28335_, _28331_);
  nor (_30893_, _28612_, _28452_);
  nor (_30895_, _30060_, _30893_);
  nor (_30896_, _30895_, _30066_);
  nor (_30897_, _30896_, _30892_);
  nor (_30898_, _30897_, _30891_);
  nor (_30899_, _30898_, _30016_);
  not (_30900_, _30892_);
  nor (_30901_, _30003_, _28614_);
  not (_30902_, _30901_);
  nor (_30903_, _30902_, _30012_);
  nor (_30904_, _30903_, _30900_);
  nor (_30905_, _30904_, _28335_);
  nor (_30906_, _30905_, _30011_);
  nor (_30907_, _27556_, _27411_);
  nand (_30908_, _30907_, _27221_);
  not (_30909_, _30908_);
  nor (_30910_, _27052_, _27504_);
  nor (_30911_, _30910_, _27556_);
  nor (_30912_, _30911_, _27466_);
  nor (_30913_, _30912_, _27221_);
  nor (_30914_, _27546_, _26925_);
  nor (_30915_, _27466_, _27462_);
  nand (_30916_, _30915_, _30914_);
  not (_30917_, _30916_);
  nor (_30918_, _30917_, _30913_);
  nor (_30919_, _30918_, _30856_);
  nor (_30920_, _30919_, _30909_);
  nor (_30921_, _30071_, _27466_);
  nor (_30922_, _30921_, _30073_);
  nor (_30923_, _30922_, _30072_);
  nor (_30924_, _30103_, _27466_);
  nand (_30926_, _30071_, _30069_);
  nand (_30927_, _30926_, _27576_);
  nand (_30928_, _30927_, _27466_);
  nor (_30929_, _26923_, _27504_);
  not (_30930_, _30929_);
  nor (_30931_, _30930_, _27271_);
  nor (_30932_, _30851_, _28313_);
  nor (_30933_, _30932_, _30931_);
  nand (_30934_, _30933_, _30928_);
  nor (_30935_, _30934_, _30924_);
  not (_30936_, _30935_);
  nor (_30937_, _30936_, _30923_);
  not (_30938_, _30937_);
  nor (_30939_, _30938_, _30920_);
  not (_30940_, _30939_);
  nor (_30941_, _30940_, _30906_);
  not (_30942_, _30941_);
  nor (_30943_, _30942_, _30899_);
  not (_30944_, _30943_);
  nor (_30945_, _26777_, _26721_);
  not (_30946_, _30945_);
  nor (_30947_, _30946_, _26640_);
  nor (_30948_, _26749_, _26677_);
  not (_30949_, _30948_);
  nor (_30950_, _30949_, _29297_);
  nand (_30952_, _30950_, _30947_);
  nor (_30953_, _26890_, _29267_);
  not (_30954_, _30953_);
  nor (_30955_, _30954_, _30952_);
  not (_30956_, _30955_);
  nor (_30957_, _30956_, _30944_);
  not (_30958_, _30889_);
  nor (_30959_, _30955_, _01710_);
  nor (_30960_, _30959_, _30958_);
  not (_30962_, _30960_);
  nor (_30963_, _30962_, _30957_);
  nor (_30965_, _30963_, _29287_);
  not (_30966_, _30965_);
  nor (_30967_, _30966_, _30890_);
  not (_30968_, _29287_);
  nor (_30972_, _03049_, _30773_);
  not (_30973_, _03049_);
  nor (_30974_, _03080_, _30973_);
  nor (_30976_, _30974_, _30972_);
  not (_30977_, _30905_);
  nor (_30979_, _03049_, _30761_);
  nor (_30980_, _03074_, _30973_);
  nor (_30982_, _30980_, _30979_);
  nand (_30983_, _30982_, _30977_);
  not (_30985_, _30983_);
  nor (_30986_, _03049_, _30765_);
  nor (_30987_, _03076_, _30973_);
  nor (_30988_, _30987_, _30986_);
  nand (_30989_, _30988_, _30985_);
  nor (_30991_, _03049_, _30769_);
  nor (_30992_, _03078_, _30973_);
  nor (_30993_, _30992_, _30991_);
  not (_30994_, _30993_);
  nor (_30996_, _30994_, _30989_);
  nand (_30998_, _30996_, _30976_);
  nor (_31000_, _03049_, _30777_);
  nor (_31001_, _03082_, _30973_);
  nor (_31002_, _31001_, _31000_);
  not (_31003_, _31002_);
  nor (_31004_, _31003_, _30998_);
  not (_31005_, _31004_);
  not (_31006_, _30998_);
  nor (_31007_, _31002_, _31006_);
  nor (_31008_, _31007_, _30011_);
  nand (_31009_, _31008_, _31005_);
  not (_31010_, _28345_);
  nor (_31011_, _30084_, _28315_);
  nand (_31012_, _31011_, _31010_);
  nor (_31013_, _29385_, _31012_);
  not (_31014_, _31013_);
  nor (_31015_, _31014_, _28096_);
  not (_31016_, _31015_);
  nor (_31017_, _31016_, _28500_);
  not (_31019_, _31017_);
  nor (_31020_, _31019_, _27645_);
  not (_31023_, _31020_);
  nor (_31024_, _31023_, _27466_);
  nor (_31025_, _27671_, _28521_);
  nor (_31026_, _27849_, _28313_);
  not (_31027_, _31026_);
  nor (_31028_, _31027_, _28452_);
  nand (_31030_, _31028_, _28401_);
  nor (_31032_, _31030_, _28123_);
  nand (_31033_, _31032_, _31025_);
  nor (_31034_, _31033_, _27225_);
  nor (_31035_, _31034_, _31024_);
  nor (_31036_, _31035_, _27081_);
  nand (_31038_, _31035_, _27081_);
  nand (_31039_, _31038_, _27506_);
  nor (_31040_, _31039_, _31036_);
  nor (_31041_, _29912_, _29907_);
  nor (_31042_, _31041_, _29957_);
  not (_31043_, _31042_);
  nor (_31044_, _31043_, _30195_);
  not (_31045_, _31044_);
  nor (_31046_, _27526_, _27225_);
  nor (_31047_, _31046_, _30102_);
  nor (_31048_, _31047_, _27081_);
  nor (_31049_, _27526_, _27016_);
  nand (_31050_, _31049_, _27225_);
  nor (_31051_, _30851_, _27271_);
  not (_31052_, _02619_);
  nor (_31053_, _29346_, _31052_);
  nor (_31054_, _31053_, _31051_);
  nand (_31055_, _31054_, _31050_);
  nor (_31056_, _31055_, _31048_);
  nand (_31057_, _31056_, _31045_);
  nor (_31058_, _31057_, _31040_);
  nand (_31059_, _31058_, _31009_);
  nor (_31060_, _31059_, _30968_);
  nor (_31061_, _31060_, _30967_);
  not (_31062_, _31061_);
  not (_31063_, _30242_);
  nor (_31065_, _31063_, _30200_);
  nand (_31067_, _31065_, _30215_);
  nand (_31069_, _30958_, _31067_);
  nor (_31070_, _29267_, _27959_);
  not (_31071_, _31070_);
  nor (_31072_, _31071_, _30952_);
  not (_31073_, _31072_);
  nor (_31074_, _31073_, _30944_);
  nor (_31075_, _31072_, _01703_);
  nor (_31076_, _31075_, _30958_);
  not (_31077_, _31076_);
  nor (_31079_, _31077_, _31074_);
  nor (_31080_, _31079_, _29287_);
  nand (_31081_, _31080_, _31069_);
  nor (_31083_, _03049_, _30780_);
  nor (_31084_, _03083_, _30973_);
  nor (_31085_, _31084_, _31083_);
  nor (_31086_, _31085_, _31004_);
  not (_31087_, _31086_);
  nand (_31088_, _31085_, _31004_);
  nand (_31089_, _31088_, _31087_);
  nor (_31090_, _31089_, _30011_);
  nor (_31091_, _31033_, _27081_);
  nand (_31092_, _31091_, _27466_);
  not (_31093_, _31092_);
  nor (_31094_, _31023_, _27040_);
  not (_31095_, _31094_);
  nor (_31096_, _31095_, _27466_);
  nor (_31097_, _31096_, _31093_);
  nor (_31098_, _31097_, _28578_);
  nand (_31099_, _31097_, _28578_);
  nand (_31100_, _31099_, _27506_);
  nor (_31101_, _31100_, _31098_);
  nor (_31102_, _29914_, _29883_);
  nor (_31103_, _31102_, _29959_);
  not (_31104_, _31103_);
  nor (_31105_, _31104_, _30195_);
  not (_31106_, _31105_);
  not (_31107_, _02855_);
  nor (_31108_, _29346_, _31107_);
  nor (_31109_, _28393_, _27466_);
  nor (_31110_, _28570_, _27225_);
  nor (_31112_, _31110_, _27526_);
  not (_31113_, _31112_);
  nor (_31114_, _31113_, _31109_);
  not (_31115_, _31114_);
  nor (_31116_, _30851_, _27476_);
  nor (_31117_, _30103_, _28578_);
  nor (_31118_, _31117_, _31116_);
  nand (_31119_, _31118_, _31115_);
  nor (_31120_, _31119_, _31108_);
  nand (_31121_, _31120_, _31106_);
  nor (_31122_, _31121_, _31101_);
  not (_31123_, _31122_);
  nor (_31124_, _31123_, _31090_);
  nand (_31125_, _31124_, _29287_);
  nand (_31126_, _31125_, _31081_);
  nand (_31127_, _31126_, _31062_);
  nor (_31128_, _30889_, _30244_);
  not (_31129_, _31080_);
  nor (_31130_, _31129_, _31128_);
  not (_31131_, _31125_);
  nor (_31132_, _31131_, _31130_);
  nand (_31133_, _31132_, _31061_);
  nand (_31134_, _31133_, _31127_);
  not (_31136_, _31088_);
  nor (_31137_, _03049_, _30783_);
  nor (_31138_, _03085_, _30973_);
  nor (_31139_, _31138_, _31137_);
  nor (_31140_, _31139_, _31136_);
  not (_31141_, _31139_);
  nor (_31142_, _31141_, _31088_);
  nor (_31143_, _31142_, _31140_);
  nand (_31145_, _31143_, _30010_);
  nor (_31146_, _31095_, _28570_);
  nor (_31147_, _31146_, _31093_);
  nor (_31148_, _31147_, _31110_);
  nor (_31149_, _31148_, _28612_);
  nand (_31151_, _31148_, _28612_);
  nand (_31152_, _31151_, _27506_);
  nor (_31153_, _31152_, _31149_);
  nor (_31154_, _29916_, _29875_);
  nor (_31156_, _31154_, _29961_);
  not (_31157_, _31156_);
  nor (_31159_, _31157_, _30195_);
  not (_31160_, _31159_);
  nand (_31161_, _29345_, _02809_);
  not (_31162_, _31161_);
  nor (_31163_, _28611_, _27225_);
  nor (_31164_, _31163_, _28458_);
  nor (_31165_, _31164_, _27526_);
  not (_31166_, _31165_);
  nor (_31167_, _30851_, _28510_);
  nor (_31168_, _30103_, _28611_);
  nor (_31169_, _31168_, _31167_);
  nand (_31170_, _31169_, _31166_);
  nor (_31171_, _31170_, _31162_);
  nand (_31172_, _31171_, _31160_);
  nor (_31173_, _31172_, _31153_);
  nand (_31174_, _31173_, _31145_);
  nand (_31175_, _31174_, _29287_);
  nand (_31177_, _30958_, _30122_);
  nor (_31179_, _26886_, _26856_);
  not (_31180_, _31179_);
  nor (_31181_, _31180_, _29267_);
  not (_31182_, _31181_);
  nor (_31183_, _31182_, _30952_);
  not (_31184_, _31183_);
  nor (_31185_, _31184_, _30943_);
  nand (_31186_, _31184_, _01740_);
  nand (_31187_, _31186_, _30889_);
  nor (_31188_, _31187_, _31185_);
  nor (_31189_, _31188_, _29287_);
  nand (_31190_, _31189_, _31177_);
  nand (_31191_, _31190_, _31175_);
  nor (_31192_, _29614_, _29507_);
  nor (_31193_, _29635_, _29527_);
  nor (_31194_, _31193_, _29519_);
  nor (_31195_, _31194_, _29642_);
  nor (_31196_, _31195_, _29649_);
  nor (_31197_, _31196_, _31192_);
  nand (_31198_, _31197_, _29345_);
  nand (_31200_, _29974_, _29940_);
  nor (_31201_, _31200_, _01880_);
  not (_31203_, _01880_);
  nor (_31205_, _29654_, _31203_);
  not (_31206_, _31205_);
  nor (_31207_, _31206_, _29939_);
  nor (_31209_, _31207_, _31201_);
  nor (_31211_, _31209_, _30195_);
  nand (_31212_, _30896_, _30892_);
  not (_31213_, _31212_);
  nor (_31214_, _31213_, _30897_);
  nor (_31215_, _31214_, _30016_);
  not (_31217_, _30903_);
  nor (_31218_, _31217_, _30892_);
  nor (_31219_, _30904_, _30011_);
  not (_31220_, _31219_);
  nor (_31221_, _31220_, _31218_);
  nor (_31222_, _30085_, _30078_);
  not (_31223_, _31222_);
  nor (_31224_, _31223_, _28315_);
  nor (_31225_, _31222_, _28313_);
  nor (_31226_, _31225_, _31224_);
  nor (_31227_, _31226_, _30072_);
  not (_31228_, _28474_);
  nor (_31229_, _30930_, _27466_);
  nor (_31230_, _30103_, _28313_);
  nand (_31231_, _30910_, _27861_);
  not (_31233_, _31231_);
  nor (_31234_, _31233_, _31230_);
  nor (_31235_, _30110_, _28452_);
  nor (_31236_, _31235_, _28478_);
  nand (_31237_, _31236_, _31234_);
  nor (_31238_, _31237_, _28475_);
  not (_31239_, _31238_);
  nor (_31240_, _31239_, _31229_);
  nand (_31241_, _31240_, _31228_);
  nor (_31242_, _31241_, _31227_);
  not (_31244_, _31242_);
  nor (_31245_, _31244_, _31221_);
  not (_31247_, _31245_);
  nor (_31249_, _31247_, _31215_);
  not (_31250_, _31249_);
  nor (_31252_, _31250_, _31211_);
  nand (_31253_, _31252_, _31198_);
  nand (_31255_, _31253_, _30958_);
  nor (_31256_, _26884_, _26856_);
  not (_31257_, _31256_);
  nor (_31258_, _31257_, _29267_);
  not (_31259_, _31258_);
  nor (_31260_, _31259_, _30952_);
  not (_31261_, _31260_);
  nor (_31262_, _31261_, _30944_);
  nor (_31263_, _31260_, _01678_);
  nor (_31264_, _31263_, _30958_);
  not (_31265_, _31264_);
  nor (_31266_, _31265_, _31262_);
  nor (_31267_, _31266_, _29287_);
  nand (_31269_, _31267_, _31255_);
  nor (_31270_, _03049_, _30736_);
  nor (_31272_, _30973_, _03047_);
  nor (_31273_, _31272_, _31270_);
  not (_31274_, _31273_);
  nand (_31276_, _31274_, _31142_);
  not (_31278_, _31276_);
  nor (_31279_, _31274_, _31142_);
  nor (_31280_, _31279_, _31278_);
  nor (_31281_, _31280_, _30011_);
  nor (_31282_, _29918_, _29867_);
  nor (_31283_, _31282_, _29963_);
  not (_31284_, _31283_);
  nor (_31286_, _31284_, _30195_);
  nand (_31287_, _31146_, _28625_);
  not (_31288_, _28401_);
  nor (_31289_, _28452_, _31288_);
  nand (_31291_, _31026_, _31289_);
  nor (_31292_, _31291_, _28123_);
  nand (_31293_, _31292_, _28500_);
  nor (_31294_, _31293_, _27671_);
  nand (_31295_, _31294_, _27040_);
  nor (_31296_, _31295_, _28578_);
  nand (_31298_, _31163_, _31296_);
  nand (_31299_, _31298_, _31287_);
  not (_31300_, _31299_);
  nor (_31301_, _31300_, _28327_);
  nor (_31302_, _31299_, _28329_);
  nor (_31303_, _31302_, _27508_);
  not (_31304_, _31303_);
  nor (_31305_, _31304_, _31301_);
  not (_31306_, _31047_);
  nand (_31307_, _31306_, _28329_);
  nand (_31308_, _27524_, _28315_);
  nor (_31309_, _31308_, _27466_);
  nor (_31310_, _30851_, _27403_);
  not (_31311_, _31310_);
  nand (_31312_, _29345_, _02586_);
  nand (_31313_, _31312_, _31311_);
  nor (_31314_, _31313_, _31309_);
  nand (_31315_, _31314_, _31307_);
  nor (_31316_, _31315_, _31305_);
  not (_31317_, _31316_);
  nor (_31318_, _31317_, _31286_);
  not (_31319_, _31318_);
  nor (_31320_, _31319_, _31281_);
  nand (_31321_, _31320_, _29287_);
  nand (_31322_, _31321_, _31269_);
  nand (_31323_, _31322_, _31191_);
  not (_31324_, _31175_);
  not (_31325_, _30015_);
  nand (_31326_, _30118_, _29977_);
  nor (_31327_, _31326_, _29652_);
  nand (_31328_, _31327_, _31325_);
  nor (_31329_, _30889_, _31328_);
  not (_31330_, _31189_);
  nor (_31331_, _31330_, _31329_);
  nor (_31332_, _31331_, _31324_);
  not (_31333_, _31192_);
  nand (_31334_, _29633_, _29520_);
  nand (_31335_, _31334_, _29524_);
  nand (_31336_, _31335_, _29614_);
  nand (_31337_, _31336_, _31333_);
  nor (_31339_, _31337_, _29346_);
  nand (_31340_, _29939_, _31203_);
  nand (_31341_, _31205_, _31200_);
  nand (_31342_, _31341_, _31340_);
  nand (_31343_, _31342_, _29653_);
  nand (_31344_, _31249_, _31343_);
  nor (_31345_, _31344_, _31339_);
  nor (_31346_, _31345_, _30889_);
  not (_31347_, _31267_);
  nor (_31348_, _31347_, _31346_);
  not (_31349_, _31279_);
  nand (_31350_, _31349_, _31276_);
  nand (_31351_, _31350_, _30010_);
  nand (_31352_, _31318_, _31351_);
  nor (_31353_, _31352_, _30968_);
  nor (_31354_, _31353_, _31348_);
  nand (_31355_, _31354_, _31332_);
  nand (_31356_, _31355_, _31323_);
  nand (_31357_, _31356_, _31134_);
  nor (_31358_, _31132_, _31061_);
  nor (_31359_, _31126_, _31062_);
  nor (_31360_, _31359_, _31358_);
  nor (_31361_, _31354_, _31332_);
  nor (_31362_, _31322_, _31191_);
  nor (_31363_, _31362_, _31361_);
  nand (_31364_, _31363_, _31360_);
  nand (_31365_, _31364_, _31357_);
  nor (_31366_, _30988_, _30985_);
  not (_31367_, _31366_);
  nand (_31368_, _31367_, _30989_);
  nor (_31369_, _31368_, _30011_);
  nor (_31370_, _27526_, _27476_);
  nor (_31371_, _29502_, _29346_);
  not (_31372_, _31371_);
  nor (_31373_, _31014_, _27466_);
  nor (_31374_, _31030_, _27225_);
  nor (_31375_, _31374_, _31373_);
  nor (_31376_, _31375_, _28096_);
  nand (_31377_, _31375_, _28096_);
  not (_31378_, _31377_);
  nor (_31380_, _31378_, _31376_);
  nor (_31381_, _31380_, _27508_);
  nor (_31382_, _29686_, _27271_);
  nor (_31383_, _31382_, _29767_);
  nor (_31384_, _31383_, _29787_);
  not (_31385_, _31384_);
  nor (_31386_, _31385_, _30195_);
  not (_31387_, _31386_);
  nor (_31388_, _30851_, _28391_);
  nor (_31389_, _30103_, _28123_);
  nor (_31390_, _31389_, _31388_);
  nand (_31391_, _31390_, _31387_);
  nor (_31392_, _31391_, _31381_);
  nand (_31393_, _31392_, _31372_);
  nor (_31394_, _31393_, _31370_);
  not (_31395_, _31394_);
  nor (_31396_, _31395_, _31369_);
  nor (_31397_, _31396_, _30968_);
  nor (_31398_, _30889_, _30828_);
  not (_31399_, _27961_);
  nor (_31400_, _30943_, _31399_);
  nor (_31401_, _26826_, _26886_);
  nand (_31402_, _31401_, _01722_);
  not (_31403_, _31402_);
  nor (_31404_, _31403_, _31400_);
  nor (_31405_, _31404_, _30952_);
  not (_31406_, _30952_);
  nor (_31407_, _31256_, _26826_);
  nand (_31408_, _31407_, _31406_);
  nand (_31409_, _31408_, _01722_);
  not (_31410_, _31409_);
  nor (_31411_, _31410_, _31405_);
  nand (_31412_, _31411_, _30889_);
  nand (_31413_, _31412_, _30968_);
  nor (_31414_, _31413_, _31398_);
  nor (_31415_, _31414_, _31397_);
  not (_31416_, _30833_);
  nand (_31417_, _30838_, _31416_);
  nand (_31418_, _31417_, _29345_);
  nand (_31419_, _30872_, _31418_);
  nand (_00003_, _30958_, _31419_);
  nor (_00004_, _30952_, _26895_);
  not (_00005_, _00004_);
  nor (_00006_, _00005_, _30944_);
  nor (_00007_, _00004_, _01728_);
  nor (_00008_, _00007_, _30958_);
  not (_00009_, _00008_);
  nor (_00010_, _00009_, _00006_);
  nor (_00011_, _00010_, _29287_);
  nand (_00012_, _00011_, _00003_);
  nor (_00013_, _29649_, _29346_);
  nor (_00014_, _30982_, _30977_);
  not (_00015_, _00014_);
  nand (_00016_, _00015_, _30983_);
  nor (_00017_, _00016_, _30011_);
  nor (_00019_, _31289_, _27225_);
  nand (_00020_, _31012_, _27225_);
  not (_00021_, _00020_);
  nor (_00023_, _00021_, _28469_);
  not (_00024_, _00023_);
  nor (_00025_, _00024_, _00019_);
  not (_00026_, _00025_);
  nor (_00027_, _00026_, _27849_);
  nor (_00028_, _00025_, _29385_);
  nor (_00029_, _00028_, _00027_);
  nand (_00030_, _00029_, _27506_);
  nor (_00031_, _27526_, _27271_);
  nor (_00032_, _30195_, _29786_);
  not (_00033_, _00032_);
  nor (_00034_, _30851_, _27016_);
  nor (_00035_, _30103_, _27849_);
  nor (_00036_, _00035_, _00034_);
  nand (_00037_, _00036_, _00033_);
  nor (_00038_, _00037_, _00031_);
  nand (_00039_, _00038_, _00030_);
  nor (_00040_, _00039_, _00017_);
  not (_00041_, _00040_);
  nor (_00042_, _00041_, _00013_);
  nand (_00043_, _00042_, _29287_);
  nand (_00044_, _00043_, _00012_);
  nand (_00046_, _00044_, _31415_);
  not (_00047_, _31415_);
  nor (_00048_, _30889_, _30876_);
  not (_00049_, _00011_);
  nor (_00050_, _00049_, _00048_);
  not (_00051_, _00043_);
  nor (_00052_, _00051_, _00050_);
  nand (_00053_, _00052_, _00047_);
  nand (_00054_, _00053_, _00046_);
  not (_00055_, _30989_);
  nor (_00056_, _30993_, _00055_);
  nor (_00057_, _30996_, _30011_);
  not (_00058_, _00057_);
  nor (_00059_, _00058_, _00056_);
  nor (_00060_, _29898_, _29896_);
  nor (_00061_, _00060_, _29900_);
  not (_00062_, _00061_);
  nor (_00063_, _00062_, _30195_);
  nor (_00064_, _31016_, _27466_);
  nand (_00065_, _31032_, _27466_);
  not (_00066_, _00065_);
  nor (_00067_, _00066_, _00064_);
  not (_00068_, _00067_);
  nor (_00069_, _00068_, _28500_);
  nor (_00070_, _00067_, _28521_);
  nor (_00071_, _00070_, _27508_);
  not (_00072_, _00071_);
  nor (_00073_, _00072_, _00069_);
  not (_00074_, _00073_);
  nor (_00075_, _27526_, _28510_);
  nor (_00076_, _30103_, _28521_);
  not (_00077_, _00076_);
  nor (_00078_, _30851_, _28452_);
  not (_00079_, _02686_);
  nor (_00080_, _29346_, _00079_);
  nor (_00081_, _00080_, _00078_);
  nand (_00082_, _00081_, _00077_);
  nor (_00083_, _00082_, _00075_);
  nand (_00084_, _00083_, _00074_);
  nor (_00085_, _00084_, _00063_);
  not (_00087_, _00085_);
  nor (_00088_, _00087_, _00059_);
  nand (_00089_, _00088_, _29287_);
  nand (_00090_, _30958_, _30692_);
  nor (_00091_, _31180_, _26826_);
  not (_00092_, _00091_);
  nor (_00093_, _00092_, _30952_);
  not (_00094_, _00093_);
  nor (_00095_, _00094_, _30944_);
  nor (_00096_, _00093_, _01718_);
  nor (_00097_, _00096_, _30958_);
  not (_00098_, _00097_);
  nor (_00099_, _00098_, _00095_);
  nor (_00100_, _00099_, _29287_);
  nand (_00101_, _00100_, _00090_);
  nand (_00102_, _00101_, _00089_);
  nor (_00103_, _30889_, _30533_);
  nor (_00104_, _31257_, _26826_);
  not (_00105_, _00104_);
  nor (_00106_, _00105_, _30952_);
  not (_00107_, _00106_);
  nor (_00108_, _00107_, _30944_);
  nor (_00109_, _00106_, _01714_);
  nor (_00110_, _00109_, _30958_);
  not (_00111_, _00110_);
  nor (_00112_, _00111_, _00108_);
  nor (_00113_, _00112_, _29287_);
  not (_00114_, _00113_);
  nor (_00115_, _00114_, _00103_);
  nor (_00116_, _30996_, _30976_);
  not (_00117_, _00116_);
  nand (_00118_, _00117_, _30998_);
  nor (_00119_, _00118_, _30011_);
  nor (_00120_, _31019_, _27466_);
  nor (_00121_, _31293_, _27225_);
  nor (_00122_, _00121_, _00120_);
  not (_00123_, _00122_);
  nor (_00124_, _00123_, _27645_);
  nor (_00125_, _00122_, _27671_);
  nor (_00126_, _00125_, _27508_);
  not (_00128_, _00126_);
  nor (_00129_, _00128_, _00124_);
  nor (_00130_, _29905_, _29900_);
  nor (_00131_, _00130_, _29953_);
  not (_00132_, _00131_);
  nor (_00133_, _00132_, _30195_);
  not (_00134_, _00133_);
  nor (_00135_, _30103_, _27671_);
  not (_00136_, _30932_);
  nor (_00137_, _27526_, _27403_);
  not (_00138_, _02652_);
  nor (_00139_, _29346_, _00138_);
  nor (_00140_, _00139_, _00137_);
  nand (_00141_, _00140_, _00136_);
  nor (_00142_, _00141_, _00135_);
  nand (_00143_, _00142_, _00134_);
  nor (_00144_, _00143_, _00129_);
  not (_00145_, _00144_);
  nor (_00146_, _00145_, _00119_);
  nand (_00147_, _00146_, _29287_);
  not (_00148_, _00147_);
  nor (_00149_, _00148_, _00115_);
  nor (_00150_, _00149_, _00102_);
  not (_00151_, _00102_);
  not (_00152_, _30502_);
  nor (_00153_, _29614_, _29572_);
  not (_00154_, _30506_);
  nor (_00156_, _30507_, _00154_);
  nor (_00157_, _00156_, _29649_);
  nor (_00159_, _00157_, _00153_);
  nor (_00160_, _00159_, _29346_);
  not (_00161_, _30530_);
  nor (_00163_, _00161_, _00160_);
  nand (_00164_, _00163_, _00152_);
  nand (_00165_, _30958_, _00164_);
  nand (_00166_, _00113_, _00165_);
  nand (_00167_, _00147_, _00166_);
  nor (_00168_, _00167_, _00151_);
  nor (_00169_, _00168_, _00150_);
  nand (_00170_, _00169_, _00054_);
  nor (_00172_, _00052_, _00047_);
  nor (_00173_, _00044_, _31415_);
  nor (_00174_, _00173_, _00172_);
  nand (_00175_, _00167_, _00151_);
  nand (_00176_, _00149_, _00102_);
  nand (_00177_, _00176_, _00175_);
  nand (_00178_, _00177_, _00174_);
  nand (_00179_, _00178_, _00170_);
  nand (_00180_, _00179_, _31365_);
  nor (_00181_, _31363_, _31360_);
  nor (_00182_, _31356_, _31134_);
  nor (_00183_, _00182_, _00181_);
  nor (_00184_, _00177_, _00174_);
  nor (_00185_, _00169_, _00054_);
  nor (_00186_, _00185_, _00184_);
  nand (_00187_, _00186_, _00183_);
  nand (_00188_, _00187_, _00180_);
  not (_00189_, _00188_);
  nor (_00190_, _00189_, _29241_);
  not (_00191_, _30531_);
  nand (_00192_, _29210_, _00191_);
  not (_00193_, _30301_);
  nand (_00194_, _29208_, _00193_);
  nand (_00195_, _00194_, _00192_);
  nor (_00196_, _00195_, _30257_);
  nand (_00197_, _29146_, _01728_);
  nor (_00198_, _29208_, _30552_);
  nor (_00199_, _29210_, _30440_);
  nor (_00200_, _00199_, _00198_);
  nand (_00202_, _00200_, _30250_);
  nand (_00203_, _00202_, _00197_);
  nor (_00205_, _00203_, _00196_);
  nand (_00206_, _29149_, _01589_);
  nand (_00208_, _29153_, _28011_);
  nand (_00209_, _00208_, _00206_);
  nor (_00210_, _29208_, _30594_);
  nor (_00211_, _29210_, _30459_);
  nor (_00212_, _00211_, _00210_);
  nand (_00213_, _00212_, _30322_);
  nor (_00214_, _29208_, _30573_);
  nor (_00216_, _29210_, _30379_);
  nor (_00217_, _00216_, _00214_);
  nand (_00218_, _00217_, _30328_);
  nand (_00219_, _00218_, _00213_);
  nor (_00220_, _00219_, _00209_);
  nand (_00221_, _00220_, _00205_);
  not (_00222_, _00158_);
  nor (_00223_, _30282_, _00222_);
  nand (_00225_, _29114_, _31210_);
  not (_00226_, _00508_);
  nor (_00227_, _29093_, _00226_);
  not (_00228_, _00464_);
  nor (_00229_, _29102_, _00228_);
  nor (_00231_, _00229_, _00227_);
  nand (_00232_, _00231_, _00225_);
  nor (_00233_, _00232_, _00223_);
  nand (_00234_, _29084_, _00289_);
  not (_00235_, _01441_);
  nor (_00237_, _29312_, _00235_);
  not (_00238_, _01295_);
  nor (_00239_, _29315_, _00238_);
  nor (_00240_, _00239_, _00237_);
  nand (_00241_, _00240_, _00234_);
  nand (_00242_, _29082_, _01469_);
  not (_00243_, _01252_);
  nor (_00244_, _30309_, _00243_);
  not (_00245_, _01423_);
  nor (_00247_, _30312_, _00245_);
  nor (_00248_, _00247_, _00244_);
  nand (_00249_, _00248_, _00242_);
  nor (_00251_, _00249_, _00241_);
  nand (_00252_, _00251_, _00233_);
  nor (_00253_, _00252_, _00221_);
  nand (_00254_, _29156_, _30761_);
  not (_00255_, _30794_);
  nor (_00257_, _29036_, _00255_);
  nand (_00258_, _29126_, _01015_);
  nand (_00259_, _29128_, _00818_);
  nand (_00260_, _00259_, _00258_);
  nor (_00261_, _00260_, _00257_);
  nand (_00263_, _00261_, _00254_);
  not (_00265_, _31277_);
  not (_00266_, _29111_);
  nor (_00267_, _00266_, _00265_);
  not (_00268_, _31204_);
  not (_00269_, _29109_);
  nor (_00271_, _00269_, _00268_);
  nor (_00272_, _00271_, _00267_);
  not (_00273_, _01185_);
  nor (_00274_, _30631_, _00273_);
  not (_00275_, _31037_);
  not (_00276_, _29134_);
  nor (_00278_, _00276_, _00275_);
  nor (_00279_, _00278_, _00274_);
  nand (_00280_, _00279_, _00272_);
  nor (_00281_, _00280_, _00263_);
  nand (_00282_, _00281_, _00253_);
  nor (_00283_, _00282_, _00190_);
  nor (_00284_, _00283_, _30880_);
  not (_00285_, _29041_);
  nand (_00286_, _29340_, _06114_);
  nand (_00287_, _00286_, _00285_);
  nor (_00288_, _00287_, _00284_);
  nor (_20930_, _00288_, _30879_);
  nand (_00290_, _06940_, _06938_);
  nor (_00292_, _00290_, _06971_);
  nand (_00293_, _00292_, _07283_);
  not (_00294_, _00292_);
  nand (_00295_, _00290_, _06971_);
  nand (_00296_, _00295_, _00294_);
  nand (_00297_, _00296_, _00293_);
  nor (_23346_, _00297_, _23698_);
  nor (_00298_, _06940_, _06938_);
  nand (_00299_, _00290_, _29344_);
  nor (_23699_, _00299_, _00298_);
  nor (_24110_, _06940_, _23698_);
  nand (_00300_, _29063_, _01263_);
  nand (_00301_, _29048_, _01303_);
  nand (_00302_, _00301_, _00300_);
  nand (_00303_, _29070_, _01345_);
  nand (_00305_, _29074_, _01268_);
  nand (_00306_, _00305_, _00303_);
  nor (_00307_, _00306_, _00302_);
  nand (_00308_, _29094_, _00327_);
  nand (_00309_, _29104_, _00453_);
  nand (_00310_, _00309_, _00308_);
  nand (_00311_, _29084_, _00382_);
  nand (_00312_, _29082_, _01307_);
  nand (_00313_, _00312_, _00311_);
  nor (_00314_, _00313_, _00310_);
  nand (_00316_, _00314_, _00307_);
  nand (_00317_, _29109_, _31150_);
  nand (_00319_, _29111_, _31078_);
  nand (_00320_, _00319_, _00317_);
  nand (_00321_, _29114_, _31082_);
  nand (_00322_, _29118_, _30978_);
  nand (_00323_, _00322_, _00321_);
  nor (_00324_, _00323_, _00320_);
  nand (_00325_, _29126_, _00878_);
  nand (_00326_, _29128_, _00916_);
  nand (_00328_, _00326_, _00325_);
  nand (_00329_, _29132_, _00834_);
  nand (_00330_, _29134_, _30999_);
  nand (_00331_, _00330_, _00329_);
  nor (_00332_, _00331_, _00328_);
  nand (_00333_, _00332_, _00324_);
  nor (_00334_, _00333_, _00316_);
  nand (_00335_, _29143_, _30702_);
  nand (_00336_, _29146_, _01678_);
  nand (_00337_, _00336_, _00335_);
  nand (_00338_, _29149_, _01617_);
  nand (_00339_, _29153_, _28664_);
  nand (_00341_, _00339_, _00338_);
  nand (_00342_, _29035_, _30743_);
  nand (_00344_, _29156_, _30736_);
  nand (_00346_, _00344_, _00342_);
  nor (_00348_, _00346_, _00341_);
  nor (_00349_, _29208_, _30283_);
  nor (_00351_, _29210_, _30285_);
  nor (_00352_, _00351_, _00349_);
  nand (_00354_, _00352_, _29163_);
  nor (_00355_, _29208_, _30288_);
  nor (_00356_, _29210_, _30290_);
  nor (_00357_, _00356_, _00355_);
  nand (_00358_, _00357_, _29218_);
  nand (_00359_, _00358_, _00354_);
  nor (_00360_, _29208_, _30277_);
  nor (_00361_, _29210_, _30279_);
  nor (_00362_, _00361_, _00360_);
  nand (_00363_, _00362_, _29224_);
  nor (_00364_, _29208_, _06713_);
  nor (_00365_, _29210_, _30424_);
  nor (_00366_, _00365_, _00364_);
  nand (_00367_, _00366_, _29232_);
  nand (_00368_, _00367_, _00363_);
  nor (_00369_, _00368_, _00359_);
  nand (_00370_, _00369_, _00348_);
  nor (_00371_, _00370_, _00337_);
  nand (_00372_, _00371_, _00334_);
  nand (_00373_, _00372_, _29305_);
  nand (_00375_, _29340_, _04368_);
  nand (_00376_, _00375_, _00373_);
  nor (_00377_, _00376_, _29041_);
  nand (_00378_, _31345_, _29041_);
  nand (_00379_, _00378_, _29344_);
  nor (_24521_, _00379_, _00377_);
  nand (_00380_, _00285_, _29344_);
  nor (_24932_, _00380_, _29305_);
  nor (_00381_, _28780_, _28718_);
  not (_00383_, _00381_);
  nor (_00384_, _00383_, _28971_);
  nand (_00385_, _00384_, _29046_);
  nor (_00386_, _00188_, _29030_);
  nand (_00387_, _29030_, _26644_);
  nand (_00388_, _00387_, _29066_);
  nor (_00389_, _00388_, _00386_);
  nand (_00391_, _29055_, _30705_);
  nand (_00392_, _28262_, _30666_);
  nand (_00393_, _00392_, _00391_);
  nand (_00394_, _00393_, _29030_);
  nor (_00396_, _29057_, _27095_);
  nor (_00397_, _29030_, _27627_);
  nor (_00398_, _00397_, _00396_);
  nor (_00399_, _00398_, _29079_);
  not (_00400_, _30670_);
  nor (_00401_, _29056_, _00400_);
  nor (_00403_, _28264_, _30541_);
  nor (_00404_, _00403_, _00401_);
  nor (_00405_, _00404_, _29030_);
  nor (_00406_, _00405_, _00399_);
  nand (_00407_, _00406_, _00394_);
  nor (_00409_, _00407_, _00389_);
  nor (_00410_, _00409_, _00385_);
  nor (_00411_, _29047_, _28970_);
  nand (_00412_, _28970_, _28782_);
  nor (_00413_, _00412_, _29046_);
  nand (_00414_, _28971_, _29087_);
  nor (_00415_, _00384_, _27457_);
  nand (_00416_, _00415_, _00414_);
  nor (_00418_, _00416_, _00413_);
  nor (_00419_, _00418_, _00411_);
  not (_00420_, _00411_);
  not (_00421_, _01249_);
  nor (_00422_, _29057_, _00421_);
  nor (_00423_, _29030_, _30592_);
  nor (_00424_, _00423_, _00422_);
  nor (_00425_, _00424_, _28264_);
  nor (_00426_, _29057_, _30307_);
  nor (_00427_, _29030_, _00243_);
  nor (_00428_, _00427_, _00426_);
  nor (_00429_, _00428_, _29067_);
  nor (_00430_, _00429_, _00425_);
  not (_00431_, _00841_);
  nor (_00432_, _29057_, _00431_);
  not (_00433_, _01229_);
  nor (_00434_, _29030_, _00433_);
  nor (_00436_, _00434_, _00432_);
  nor (_00437_, _00436_, _29056_);
  not (_00438_, _01345_);
  nor (_00439_, _29057_, _00438_);
  not (_00442_, _01224_);
  nor (_00443_, _29030_, _00442_);
  nor (_00444_, _00443_, _00439_);
  nor (_00445_, _00444_, _29079_);
  nor (_00446_, _00445_, _00437_);
  nand (_00447_, _00446_, _00430_);
  nor (_00448_, _00447_, _00420_);
  nor (_00449_, _00448_, _00419_);
  nor (_00450_, _29089_, _28845_);
  not (_00451_, _00412_);
  nand (_00452_, _00451_, _00450_);
  nand (_00454_, _00352_, _29030_);
  nand (_00455_, _30449_, _29057_);
  nand (_00456_, _00455_, _00454_);
  nand (_00457_, _00456_, _29078_);
  nand (_00458_, _30167_, _29030_);
  nand (_00459_, _30745_, _29057_);
  nand (_00460_, _00459_, _00458_);
  nand (_00461_, _00460_, _29055_);
  nand (_00462_, _00461_, _00457_);
  nand (_00463_, _30332_, _29030_);
  nand (_00465_, _00217_, _29057_);
  nand (_00466_, _00465_, _00463_);
  nand (_00467_, _00466_, _29066_);
  nand (_00468_, _29212_, _29030_);
  nand (_00469_, _30626_, _29057_);
  nand (_00470_, _00469_, _00468_);
  nand (_00471_, _00470_, _28262_);
  nand (_00472_, _00471_, _00467_);
  nor (_00474_, _00472_, _00462_);
  nor (_00475_, _00474_, _00452_);
  nor (_00476_, _00383_, _28970_);
  nand (_00477_, _00476_, _00450_);
  not (_00478_, _00453_);
  nor (_00479_, _29057_, _00478_);
  not (_00480_, _00246_);
  nor (_00481_, _29030_, _00480_);
  nor (_00482_, _00481_, _00479_);
  nor (_00483_, _00482_, _29079_);
  nor (_00484_, _29057_, _30291_);
  nor (_00486_, _29030_, _00228_);
  nor (_00487_, _00486_, _00484_);
  nor (_00488_, _00487_, _29067_);
  not (_00489_, _00402_);
  nor (_00490_, _29057_, _00489_);
  nor (_00491_, _29030_, _30608_);
  nor (_00492_, _00491_, _00490_);
  nor (_00493_, _00492_, _28264_);
  nor (_00494_, _00493_, _00488_);
  nand (_00496_, _29030_, _00204_);
  nand (_00497_, _29057_, _00435_);
  nand (_00498_, _00497_, _00496_);
  nand (_00499_, _00498_, _29055_);
  nand (_00500_, _00499_, _00494_);
  nor (_00501_, _00500_, _00483_);
  nor (_00502_, _00501_, _00477_);
  nor (_00503_, _00502_, _00475_);
  nor (_00504_, _29282_, _29293_);
  nand (_00505_, _00476_, _28906_);
  not (_00506_, _00762_);
  nor (_00507_, _29057_, _00506_);
  not (_00509_, _00920_);
  nor (_00510_, _29030_, _00509_);
  nor (_00511_, _00510_, _00507_);
  nor (_00513_, _00511_, _29056_);
  not (_00514_, _00784_);
  nor (_00515_, _29057_, _00514_);
  not (_00516_, _00818_);
  nor (_00518_, _29030_, _00516_);
  nor (_00519_, _00518_, _00515_);
  nor (_00520_, _00519_, _29067_);
  not (_00521_, _00801_);
  nor (_00522_, _29057_, _00521_);
  not (_00523_, _00929_);
  nor (_00524_, _29030_, _00523_);
  nor (_00525_, _00524_, _00522_);
  nor (_00526_, _00525_, _28264_);
  nor (_00527_, _00526_, _00520_);
  nand (_00528_, _29030_, _00916_);
  nand (_00529_, _29057_, _00941_);
  nand (_00531_, _00529_, _00528_);
  nand (_00532_, _00531_, _29078_);
  nand (_00533_, _00532_, _00527_);
  nor (_00534_, _00533_, _00513_);
  nor (_00535_, _00534_, _00505_);
  nor (_00536_, _00535_, _00504_);
  nand (_00537_, _00536_, _00503_);
  nor (_00538_, _00537_, _00449_);
  not (_00539_, _28906_);
  not (_00540_, _00384_);
  nand (_00541_, _30253_, _29030_);
  nand (_00542_, _00200_, _29057_);
  nand (_00543_, _00542_, _00541_);
  nand (_00544_, _00543_, _29066_);
  nand (_00545_, _00362_, _29030_);
  nand (_00547_, _30461_, _29057_);
  nand (_00548_, _00547_, _00545_);
  nand (_00550_, _00548_, _29078_);
  nand (_00552_, _00550_, _00544_);
  nand (_00553_, _30177_, _29030_);
  nand (_00555_, _30754_, _29057_);
  nand (_00557_, _00555_, _00553_);
  nand (_00558_, _00557_, _29055_);
  nand (_00560_, _29223_, _29030_);
  nand (_00562_, _30547_, _29057_);
  nand (_00563_, _00562_, _00560_);
  nand (_00564_, _00563_, _28262_);
  nand (_00566_, _00564_, _00558_);
  nor (_00567_, _00566_, _00552_);
  nor (_00568_, _00567_, _00540_);
  nand (_00569_, _30261_, _29030_);
  nor (_00570_, _29208_, _30531_);
  nor (_00571_, _29210_, _30301_);
  nor (_00572_, _00571_, _00570_);
  nand (_00573_, _00572_, _29057_);
  nand (_00574_, _00573_, _00569_);
  nand (_00575_, _00574_, _29066_);
  nand (_00576_, _00366_, _29030_);
  nand (_00577_, _30465_, _29057_);
  nand (_00578_, _00577_, _00576_);
  nand (_00580_, _00578_, _29078_);
  nand (_00581_, _00580_, _00575_);
  nand (_00582_, _30181_, _29030_);
  nand (_00583_, _30758_, _29057_);
  nand (_00584_, _00583_, _00582_);
  nand (_00585_, _00584_, _29055_);
  nand (_00586_, _29231_, _29030_);
  nand (_00587_, _30553_, _29057_);
  nand (_00588_, _00587_, _00586_);
  nand (_00589_, _00588_, _28262_);
  nand (_00590_, _00589_, _00585_);
  nor (_00591_, _00590_, _00581_);
  nor (_00592_, _00591_, _00412_);
  nor (_00593_, _00592_, _00568_);
  nor (_00594_, _00593_, _00539_);
  nand (_00595_, _28971_, _28782_);
  not (_00596_, _00343_);
  nor (_00597_, _29057_, _00596_);
  not (_00598_, _00517_);
  nor (_00599_, _29030_, _00598_);
  nor (_00600_, _00599_, _00597_);
  nor (_00601_, _00600_, _29056_);
  not (_00602_, _30981_);
  nor (_00603_, _29057_, _00602_);
  not (_00604_, _00315_);
  nor (_00605_, _29030_, _00604_);
  nor (_00606_, _00605_, _00603_);
  nor (_00607_, _00606_, _28264_);
  not (_00608_, _30975_);
  nor (_00609_, _29057_, _00608_);
  not (_00610_, _00289_);
  nor (_00611_, _29030_, _00610_);
  nor (_00612_, _00611_, _00609_);
  nor (_00613_, _00612_, _29067_);
  nor (_00614_, _00613_, _00607_);
  nand (_00615_, _29030_, _00382_);
  nand (_00616_, _29057_, _00512_);
  nand (_00617_, _00616_, _00615_);
  nand (_00618_, _00617_, _29078_);
  nand (_00619_, _00618_, _00614_);
  nor (_00621_, _00619_, _00601_);
  nor (_00622_, _00621_, _00539_);
  not (_00623_, _00450_);
  not (_00624_, _00327_);
  nor (_00625_, _29057_, _00624_);
  not (_00626_, _00224_);
  nor (_00628_, _29030_, _00626_);
  nor (_00629_, _00628_, _00625_);
  nor (_00630_, _00629_, _29079_);
  not (_00631_, _00390_);
  nor (_00632_, _29057_, _00631_);
  nor (_00633_, _29030_, _30605_);
  nor (_00634_, _00633_, _00632_);
  nor (_00635_, _00634_, _28264_);
  nor (_00636_, _29057_, _30287_);
  nor (_00637_, _29030_, _00226_);
  nor (_00638_, _00637_, _00636_);
  nor (_00639_, _00638_, _29067_);
  nor (_00640_, _00639_, _00635_);
  nand (_00642_, _29030_, _00207_);
  nand (_00643_, _29057_, _00250_);
  nand (_00644_, _00643_, _00642_);
  nand (_00645_, _00644_, _29055_);
  nand (_00646_, _00645_, _00640_);
  nor (_00647_, _00646_, _00630_);
  nor (_00648_, _00647_, _00623_);
  nor (_00649_, _00648_, _00622_);
  nor (_00650_, _00649_, _00595_);
  nand (_00651_, _00450_, _00384_);
  nand (_00652_, _30326_, _29030_);
  nand (_00653_, _00212_, _29057_);
  nand (_00654_, _00653_, _00652_);
  nand (_00655_, _00654_, _29066_);
  nand (_00656_, _00357_, _29030_);
  nand (_00657_, _30454_, _29057_);
  nand (_00658_, _00657_, _00656_);
  nand (_00659_, _00658_, _29078_);
  nand (_00660_, _00659_, _00655_);
  nand (_00661_, _30171_, _29030_);
  nand (_00662_, _30749_, _29057_);
  nand (_00664_, _00662_, _00661_);
  nand (_00665_, _00664_, _29055_);
  nand (_00666_, _29216_, _29030_);
  nand (_00667_, _30622_, _29057_);
  nand (_00668_, _00667_, _00666_);
  nand (_00669_, _00668_, _28262_);
  nand (_00670_, _00669_, _00665_);
  nor (_00671_, _00670_, _00660_);
  nor (_00672_, _00671_, _00651_);
  nor (_00673_, _00672_, _00650_);
  nor (_00674_, _29089_, _28844_);
  nand (_00675_, _00674_, _00384_);
  not (_00676_, _01617_);
  nor (_00677_, _29057_, _00676_);
  not (_00678_, _01620_);
  nor (_00679_, _29030_, _00678_);
  nor (_00680_, _00679_, _00677_);
  nor (_00681_, _00680_, _29079_);
  nor (_00682_, _29057_, _30272_);
  not (_00683_, _01589_);
  nor (_00684_, _29030_, _00683_);
  nor (_00685_, _00684_, _00682_);
  nor (_00686_, _00685_, _29067_);
  not (_00687_, _01609_);
  nor (_00688_, _29057_, _00687_);
  nor (_00689_, _29030_, _30569_);
  nor (_00690_, _00689_, _00688_);
  nor (_00691_, _00690_, _28264_);
  nor (_00692_, _00691_, _00686_);
  nand (_00693_, _29030_, _01585_);
  nand (_00694_, _29057_, _01597_);
  nand (_00695_, _00694_, _00693_);
  nand (_00696_, _00695_, _29055_);
  nand (_00697_, _00696_, _00692_);
  nor (_00698_, _00697_, _00681_);
  nor (_00699_, _00698_, _00675_);
  nand (_00700_, _00674_, _00451_);
  nor (_00701_, _29057_, _28301_);
  nor (_00702_, _29030_, _27391_);
  nor (_00703_, _00702_, _00701_);
  nor (_00705_, _00703_, _29079_);
  nor (_00706_, _29057_, _30248_);
  not (_00707_, _01728_);
  nor (_00708_, _29030_, _00707_);
  nor (_00709_, _00708_, _00706_);
  nor (_00710_, _00709_, _29067_);
  nor (_00711_, _29057_, _28436_);
  nor (_00712_, _29030_, _27340_);
  nor (_00713_, _00712_, _00711_);
  nor (_00714_, _00713_, _28264_);
  nor (_00715_, _00714_, _00710_);
  nand (_00716_, _29030_, _01703_);
  nand (_00717_, _29057_, _01722_);
  nand (_00718_, _00717_, _00716_);
  nand (_00719_, _00718_, _29055_);
  nand (_00720_, _00719_, _00715_);
  nor (_00721_, _00720_, _00705_);
  nor (_00722_, _00721_, _00700_);
  nor (_00723_, _00722_, _00699_);
  nand (_00724_, _00723_, _00673_);
  nor (_00725_, _00724_, _00594_);
  nand (_00726_, _00725_, _00538_);
  nor (_00727_, _00726_, _00410_);
  nor (_00728_, _31258_, _26789_);
  nand (_00729_, _00728_, _29265_);
  not (_00730_, _00729_);
  nor (_00731_, _00700_, _29289_);
  nor (_00732_, _00731_, _00730_);
  nand (_00733_, _00504_, _30943_);
  nand (_00734_, _00733_, _00732_);
  nor (_00735_, _00734_, _00727_);
  nor (_00736_, _29057_, _28481_);
  nor (_00737_, _29030_, _27718_);
  nor (_00738_, _00737_, _00736_);
  nor (_00739_, _00738_, _29079_);
  nor (_00740_, _29057_, _28639_);
  nor (_00741_, _29030_, _28540_);
  nor (_00742_, _00741_, _00740_);
  nor (_00743_, _00742_, _28264_);
  nor (_00744_, _29057_, _27584_);
  nor (_00746_, _29030_, _27888_);
  nor (_00747_, _00746_, _00744_);
  nor (_00748_, _00747_, _29067_);
  nor (_00749_, _00748_, _00743_);
  not (_00750_, _28598_);
  nand (_00751_, _29030_, _00750_);
  nand (_00752_, _29057_, _28244_);
  nand (_00753_, _00752_, _00751_);
  nand (_00754_, _00753_, _29055_);
  nand (_00755_, _00754_, _00749_);
  nor (_00756_, _00755_, _00739_);
  nor (_00757_, _00756_, _00732_);
  nor (_00758_, _00757_, _00735_);
  nor (_25343_, _00758_, _23698_);
  nand (_00759_, _00294_, _29344_);
  not (_00760_, _07283_);
  nand (_00761_, _00290_, _00760_);
  not (_00763_, _00290_);
  nand (_00764_, _00763_, _07283_);
  nand (_00766_, _00764_, _00761_);
  nor (_25917_, _00766_, _00759_);
  nor (_26728_, _00293_, _23698_);
  nor (_00767_, _27726_, _26642_);
  not (_00768_, _00767_);
  nor (_00769_, _27610_, _26677_);
  nand (_00770_, _00769_, _29298_);
  nor (_00771_, _00770_, _00768_);
  nand (_00772_, _00771_, _31258_);
  nor (_00773_, _00772_, _30944_);
  nor (_00774_, _26677_, _26642_);
  nand (_00775_, _00774_, _27953_);
  not (_00777_, _00775_);
  nor (_00778_, _31259_, _26793_);
  nand (_00779_, _00778_, _00777_);
  nand (_00780_, _00772_, _00478_);
  nand (_00781_, _00780_, _00779_);
  nor (_00782_, _00781_, _00773_);
  nor (_00783_, _30946_, _26642_);
  nand (_00785_, _00783_, _00769_);
  nor (_00786_, _00785_, _31259_);
  nand (_00788_, _00786_, _26787_);
  nor (_00789_, _00788_, _28481_);
  nor (_00790_, _00789_, _00782_);
  nor (_27539_, _00790_, _23698_);
  not (_00792_, _27951_);
  nor (_00793_, _27614_, _00792_);
  nor (_00794_, _31399_, _27726_);
  not (_00795_, _00794_);
  nor (_00796_, _00795_, _26785_);
  nand (_00797_, _00796_, _00793_);
  nand (_00798_, _00797_, _28740_);
  nand (_00799_, _00798_, _29344_);
  not (_00800_, _27584_);
  nor (_00802_, _00797_, _00800_);
  nor (_28350_, _00802_, _00799_);
  nand (_00804_, _00797_, _28919_);
  nand (_00805_, _00804_, _29344_);
  nor (_00807_, _00797_, _27742_);
  nor (_28815_, _00807_, _00805_);
  nand (_00808_, _00797_, _28990_);
  nand (_00809_, _00808_, _29344_);
  not (_00811_, _28540_);
  nor (_00812_, _00797_, _00811_);
  nor (_29227_, _00812_, _00809_);
  nand (_00815_, _00797_, _28232_);
  nand (_00816_, _00815_, _29344_);
  nor (_00817_, _00797_, _28244_);
  nor (_29639_, _00817_, _00816_);
  nor (_00819_, _00797_, _27886_);
  nand (_00820_, _00797_, _27782_);
  nand (_00821_, _00820_, _29344_);
  nor (_30050_, _00821_, _00819_);
  nand (_00822_, _26783_, _26777_);
  nor (_00823_, _00822_, _26895_);
  nand (_00825_, _00823_, _00793_);
  nand (_00826_, _00825_, _28795_);
  nand (_00827_, _00826_, _29344_);
  not (_00828_, _28639_);
  nor (_00829_, _00825_, _00828_);
  nor (_30492_, _00829_, _00827_);
  nand (_00832_, _00825_, _28863_);
  nand (_00833_, _00832_, _29344_);
  nor (_00835_, _00825_, _00750_);
  nor (_30969_, _00835_, _00833_);
  nand (_00836_, _00825_, _28756_);
  nand (_00837_, _00836_, _29344_);
  nor (_00838_, _00825_, _00800_);
  nor (_00001_, _00838_, _00837_);
  nand (_00840_, _00825_, _28935_);
  nand (_00842_, _00840_, _29344_);
  nor (_00843_, _00825_, _27742_);
  nor (_00440_, _00843_, _00842_);
  nand (_00844_, _00825_, _29001_);
  nand (_00845_, _00844_, _29344_);
  nor (_00846_, _00825_, _00811_);
  nor (_00871_, _00846_, _00845_);
  nand (_00849_, _00825_, _28206_);
  nand (_00850_, _00849_, _29344_);
  nor (_00851_, _00825_, _28244_);
  nor (_01281_, _00851_, _00850_);
  nor (_00852_, _26895_, _27726_);
  not (_00853_, _00852_);
  nor (_00854_, _00853_, _26785_);
  nand (_00855_, _00854_, _00793_);
  nor (_00856_, _00855_, _27886_);
  nand (_00857_, _00855_, _27809_);
  nand (_00858_, _00857_, _29344_);
  nor (_01726_, _00858_, _00856_);
  nor (_00860_, _27963_, _26785_);
  nand (_00861_, _00860_, _00793_);
  nor (_00862_, _00861_, _00828_);
  nand (_00863_, _00861_, _28803_);
  nand (_00864_, _00863_, _29344_);
  nor (_02159_, _00864_, _00862_);
  nor (_00865_, _00861_, _00750_);
  nand (_00866_, _00861_, _28853_);
  nand (_00867_, _00866_, _29344_);
  nor (_02541_, _00867_, _00865_);
  nor (_00868_, _00861_, _00800_);
  nand (_00870_, _00861_, _28742_);
  nand (_00873_, _00870_, _29344_);
  nor (_02878_, _00873_, _00868_);
  nor (_00874_, _00861_, _27742_);
  nand (_00875_, _00861_, _28921_);
  nand (_00876_, _00875_, _29344_);
  nor (_03289_, _00876_, _00874_);
  nor (_00879_, _00861_, _00811_);
  nand (_00880_, _00861_, _28994_);
  nand (_00881_, _00880_, _29344_);
  nor (_03630_, _00881_, _00879_);
  nor (_00882_, _00861_, _28244_);
  nand (_00883_, _00861_, _28222_);
  nand (_00884_, _00883_, _29344_);
  nor (_04029_, _00884_, _00882_);
  nor (_00885_, _00861_, _27886_);
  nand (_00886_, _00861_, _27793_);
  nand (_00887_, _00886_, _29344_);
  nor (_04419_, _00887_, _00885_);
  not (_00889_, _30881_);
  nor (_00890_, _00889_, _26785_);
  nand (_00891_, _00890_, _00793_);
  nor (_00892_, _00891_, _00828_);
  nand (_00893_, _00891_, _28797_);
  nand (_00895_, _00893_, _29344_);
  nor (_04830_, _00895_, _00892_);
  nor (_00896_, _00891_, _00750_);
  nand (_00897_, _00891_, _28858_);
  nand (_00898_, _00897_, _29344_);
  nor (_05287_, _00898_, _00896_);
  nor (_00899_, _00891_, _00800_);
  nand (_00901_, _00891_, _28751_);
  nand (_00902_, _00901_, _29344_);
  nor (_05725_, _00902_, _00899_);
  nor (_00903_, _00891_, _27742_);
  nand (_00905_, _00891_, _28930_);
  nand (_00906_, _00905_, _29344_);
  nor (_06160_, _00906_, _00903_);
  nor (_00907_, _00891_, _00811_);
  nand (_00908_, _00891_, _28996_);
  nand (_00909_, _00908_, _29344_);
  nor (_06634_, _00909_, _00907_);
  nor (_00911_, _00891_, _28244_);
  nand (_00912_, _00891_, _28200_);
  nand (_00913_, _00912_, _29344_);
  nor (_07049_, _00913_, _00911_);
  nor (_00914_, _00891_, _27886_);
  nand (_00915_, _00891_, _27799_);
  nand (_00917_, _00915_, _29344_);
  nor (_07422_, _00917_, _00914_);
  nor (_00918_, _27614_, _26683_);
  nand (_00919_, _00918_, _00796_);
  nand (_00921_, _00919_, _28848_);
  nand (_00922_, _00921_, _29344_);
  nor (_00923_, _00919_, _00750_);
  nor (_07840_, _00923_, _00922_);
  nand (_00924_, _00919_, _28745_);
  nand (_00925_, _00924_, _29344_);
  nor (_00926_, _00919_, _00800_);
  nor (_08287_, _00926_, _00925_);
  nand (_00927_, _00919_, _28924_);
  nand (_00928_, _00927_, _29344_);
  nor (_00930_, _00919_, _27742_);
  nor (_08791_, _00930_, _00928_);
  nand (_00931_, _00919_, _28988_);
  nand (_00932_, _00931_, _29344_);
  nor (_00933_, _00919_, _00811_);
  nor (_09311_, _00933_, _00932_);
  nand (_00934_, _00919_, _28196_);
  nand (_00935_, _00934_, _29344_);
  nor (_00936_, _00919_, _28244_);
  nor (_09801_, _00936_, _00935_);
  nor (_00937_, _00919_, _27886_);
  nand (_00938_, _00919_, _27764_);
  nand (_00939_, _00938_, _29344_);
  nor (_10212_, _00939_, _00937_);
  nand (_00940_, _00918_, _00860_);
  nor (_00942_, _00940_, _00800_);
  nand (_00943_, _00940_, _28747_);
  nand (_00944_, _00943_, _29344_);
  nor (_10627_, _00944_, _00942_);
  nor (_00946_, _00940_, _27742_);
  nand (_00948_, _00940_, _28937_);
  nand (_00949_, _00948_, _29344_);
  nor (_11040_, _00949_, _00946_);
  nand (_00950_, _00918_, _00823_);
  nand (_00951_, _00950_, _28806_);
  nand (_00952_, _00951_, _29344_);
  nor (_00954_, _00950_, _00828_);
  nor (_11450_, _00954_, _00952_);
  nand (_00955_, _00950_, _28851_);
  nand (_00956_, _00955_, _29344_);
  nor (_00957_, _00950_, _00750_);
  nor (_11861_, _00957_, _00956_);
  nor (_00958_, _00940_, _00811_);
  nand (_00959_, _00940_, _28983_);
  nand (_00960_, _00959_, _29344_);
  nor (_12271_, _00960_, _00958_);
  nor (_00962_, _00940_, _28244_);
  nand (_00964_, _00940_, _28210_);
  nand (_00965_, _00964_, _29344_);
  nor (_12683_, _00965_, _00962_);
  nand (_00966_, _00950_, _28753_);
  nand (_00967_, _00966_, _29344_);
  nor (_00968_, _00950_, _00800_);
  nor (_13094_, _00968_, _00967_);
  nand (_00969_, _00950_, _28932_);
  nand (_00970_, _00969_, _29344_);
  nor (_00972_, _00950_, _27742_);
  nor (_13505_, _00972_, _00970_);
  nor (_00974_, _00940_, _27886_);
  nand (_00975_, _00940_, _27774_);
  nand (_00976_, _00975_, _29344_);
  nor (_13872_, _00976_, _00974_);
  nand (_00977_, _00918_, _00890_);
  nor (_00979_, _00977_, _00828_);
  nand (_00980_, _00977_, _28801_);
  nand (_00982_, _00980_, _29344_);
  nor (_14206_, _00982_, _00979_);
  nand (_00984_, _00950_, _28999_);
  nand (_00986_, _00984_, _29344_);
  nor (_00989_, _00950_, _00811_);
  nor (_14541_, _00989_, _00986_);
  nand (_00991_, _00950_, _28228_);
  nand (_00993_, _00991_, _29344_);
  nor (_00994_, _00950_, _28244_);
  nor (_14862_, _00994_, _00993_);
  nand (_00997_, _00918_, _00854_);
  nor (_00998_, _00997_, _27886_);
  nand (_00999_, _00997_, _27756_);
  nand (_01001_, _00999_, _29344_);
  nor (_15140_, _01001_, _00998_);
  nor (_01002_, _00940_, _00828_);
  nand (_01003_, _00940_, _28792_);
  nand (_01004_, _01003_, _29344_);
  nor (_15412_, _01004_, _01002_);
  nor (_01005_, _00940_, _00750_);
  nand (_01006_, _00940_, _28865_);
  nand (_01007_, _01006_, _29344_);
  nor (_15688_, _01007_, _01005_);
  nand (_01008_, _00919_, _28790_);
  nand (_01009_, _01008_, _29344_);
  nor (_01010_, _00919_, _00828_);
  nor (_15972_, _01010_, _01009_);
  nor (_01011_, _00891_, _28482_);
  nand (_01012_, _00891_, _28689_);
  nand (_01014_, _01012_, _29344_);
  nor (_16254_, _01014_, _01011_);
  nand (_01017_, _00797_, _28860_);
  nand (_01019_, _01017_, _29344_);
  nor (_01021_, _00797_, _00750_);
  nor (_16542_, _01021_, _01019_);
  nand (_01024_, _00797_, _28808_);
  nand (_01026_, _01024_, _29344_);
  nor (_01028_, _00797_, _00828_);
  nor (_16828_, _01028_, _01026_);
  nor (_01031_, _00977_, _27886_);
  nand (_01033_, _00977_, _27815_);
  nand (_01035_, _01033_, _29344_);
  nor (_17114_, _01035_, _01031_);
  nor (_01037_, _00977_, _28244_);
  nand (_01040_, _00977_, _28218_);
  nand (_01041_, _01040_, _29344_);
  nor (_17403_, _01041_, _01037_);
  nor (_01043_, _00977_, _00811_);
  nand (_01044_, _00977_, _28985_);
  nand (_01045_, _01044_, _29344_);
  nor (_17689_, _01045_, _01043_);
  nor (_01046_, _00977_, _27742_);
  nand (_01047_, _00977_, _28926_);
  nand (_01048_, _01047_, _29344_);
  nor (_17976_, _01048_, _01046_);
  nor (_01049_, _00977_, _00800_);
  nand (_01050_, _00977_, _28758_);
  nand (_01051_, _01050_, _29344_);
  nor (_18264_, _01051_, _01049_);
  nor (_01052_, _00977_, _00750_);
  nand (_01053_, _00977_, _28846_);
  nand (_01054_, _01053_, _29344_);
  nor (_18551_, _01054_, _01052_);
  nand (_01055_, _00919_, _28701_);
  nand (_01056_, _01055_, _29344_);
  nor (_01057_, _00919_, _28482_);
  nor (_18911_, _01057_, _01056_);
  nand (_01058_, _00950_, _28699_);
  nand (_01059_, _01058_, _29344_);
  nor (_01060_, _00950_, _28482_);
  nor (_19310_, _01060_, _01059_);
  nor (_01061_, _00940_, _28482_);
  nand (_01062_, _00940_, _28706_);
  nand (_01063_, _01062_, _29344_);
  nor (_19712_, _01063_, _01061_);
  nor (_01064_, _00977_, _28482_);
  nand (_01065_, _00977_, _28704_);
  nand (_01066_, _01065_, _29344_);
  nor (_20122_, _01066_, _01064_);
  nand (_01067_, _00797_, _28693_);
  nand (_01068_, _01067_, _29344_);
  nor (_01069_, _00797_, _28482_);
  nor (_20533_, _01069_, _01068_);
  nand (_01070_, _00825_, _28695_);
  nand (_01072_, _01070_, _29344_);
  nor (_01073_, _00825_, _28482_);
  nor (_20931_, _01073_, _01072_);
  nor (_01074_, _00861_, _28482_);
  nand (_01075_, _00861_, _28687_);
  nand (_01076_, _01075_, _29344_);
  nor (_21320_, _01076_, _01074_);
  nor (_21708_, _28260_, _23698_);
  nor (_22100_, _29053_, _23698_);
  nor (_01077_, _27103_, _29293_);
  nand (_01078_, _01077_, _27166_);
  nor (_01079_, _01078_, _30943_);
  nand (_01080_, _00828_, _29293_);
  nand (_01081_, _27166_, _06243_);
  nor (_01082_, _27176_, _29293_);
  nand (_01083_, _01082_, _01081_);
  nand (_01084_, _01083_, _01080_);
  nor (_01085_, _01084_, _01079_);
  nor (_22521_, _01085_, _23698_);
  nand (_01086_, _01077_, _27138_);
  nor (_01087_, _01086_, _30943_);
  nand (_01088_, _00750_, _29293_);
  nand (_01089_, _27138_, _06243_);
  nor (_01090_, _27148_, _29293_);
  nand (_01091_, _01090_, _01089_);
  nand (_01092_, _01091_, _01088_);
  nor (_01093_, _01092_, _01087_);
  nor (_22942_, _01093_, _23698_);
  nand (_01094_, _01077_, _27117_);
  nor (_01095_, _01094_, _30943_);
  nand (_01096_, _00800_, _29293_);
  nor (_01097_, _27429_, _29293_);
  nand (_01098_, _01097_, _26980_);
  nand (_01099_, _01098_, _01096_);
  nor (_01100_, _01099_, _01095_);
  nor (_23263_, _01100_, _23698_);
  not (_01101_, _27200_);
  nor (_01102_, _06243_, _29293_);
  nand (_01103_, _01102_, _01101_);
  nor (_01104_, _01103_, _30943_);
  nand (_01106_, _27742_, _29293_);
  nor (_01107_, _27425_, _29293_);
  nand (_01108_, _01107_, _27206_);
  nand (_01109_, _01108_, _01106_);
  nor (_01110_, _01109_, _01104_);
  nor (_23284_, _01110_, _23698_);
  nand (_01111_, _01102_, _27166_);
  nor (_01112_, _01111_, _30943_);
  nand (_01113_, _00811_, _29293_);
  nand (_01114_, _01102_, _27164_);
  not (_01115_, _01103_);
  nor (_01116_, _01115_, _01077_);
  nand (_01117_, _01116_, _01114_);
  nand (_01118_, _01117_, _27160_);
  nand (_01119_, _01118_, _01113_);
  nor (_01120_, _01119_, _01112_);
  nor (_23304_, _01120_, _23698_);
  nand (_01121_, _01102_, _27138_);
  nor (_01122_, _01121_, _30943_);
  nand (_01123_, _28244_, _29293_);
  nand (_01124_, _27138_, _27103_);
  nor (_01125_, _28111_, _29293_);
  nand (_01126_, _01125_, _01124_);
  nand (_01127_, _01126_, _01123_);
  nor (_01128_, _01127_, _01122_);
  nor (_23325_, _01128_, _23698_);
  nor (_01129_, _01114_, _06269_);
  not (_01130_, _01129_);
  nor (_01131_, _01130_, _30943_);
  nand (_01132_, _27886_, _29293_);
  nor (_01133_, _27435_, _29293_);
  nand (_01134_, _01133_, _27251_);
  nand (_01135_, _01134_, _01132_);
  nor (_01136_, _01135_, _01131_);
  nor (_23347_, _01136_, _23698_);
  not (_01137_, _26306_);
  nor (_01138_, _26290_, _25601_);
  nor (_01139_, _01138_, _01137_);
  nor (_01140_, _01139_, _26464_);
  not (_01141_, _26237_);
  nor (_01143_, _29189_, _29181_);
  nand (_01144_, _01143_, _01141_);
  not (_01145_, _26270_);
  nor (_01146_, _26412_, _01145_);
  nor (_01147_, _26156_, _26244_);
  nor (_01148_, _01147_, _26357_);
  nand (_01149_, _01148_, _01146_);
  nor (_01150_, _01149_, _01144_);
  nor (_01151_, _01150_, _25601_);
  nor (_01152_, _01151_, _01140_);
  nor (_23376_, _01152_, _23698_);
  nor (_01153_, _28482_, _30308_);
  nand (_01154_, _01077_, _01101_);
  nand (_01155_, _27196_, _30308_);
  nand (_01156_, _01155_, _01154_);
  nor (_01157_, _01156_, _01153_);
  nor (_01158_, _01154_, _30943_);
  nor (_01159_, _01158_, _01157_);
  nor (_23417_, _01159_, _23698_);
  nor (_01160_, _27608_, _29293_);
  not (_01161_, _01160_);
  nor (_01162_, _01161_, _26642_);
  nor (_01163_, _26856_, _30308_);
  nor (_01164_, _01163_, _01162_);
  not (_01165_, _01164_);
  nor (_01166_, _26171_, _26306_);
  nor (_01167_, _26266_, _26244_);
  nor (_01168_, _01167_, _29181_);
  not (_01169_, _01168_);
  nor (_01170_, _01169_, _01145_);
  not (_01171_, _01170_);
  nand (_01172_, _26296_, _26290_);
  not (_01173_, _01172_);
  nor (_01174_, _25884_, _25708_);
  nand (_01175_, _01174_, _26148_);
  nor (_01176_, _01175_, _26244_);
  nor (_01177_, _01176_, _26304_);
  nand (_01178_, _01177_, _01173_);
  nor (_01179_, _01178_, _01171_);
  not (_01180_, _01179_);
  not (_01182_, _26365_);
  nor (_01183_, _01182_, _26235_);
  nor (_01184_, _01175_, _26181_);
  nand (_01186_, _26377_, _26150_);
  nor (_01188_, _01186_, _26244_);
  nor (_01190_, _01188_, _01184_);
  nand (_01192_, _01190_, _01183_);
  nor (_01194_, _01192_, _01180_);
  nor (_01196_, _01194_, _25601_);
  nor (_01198_, _01196_, _01166_);
  not (_01199_, _01198_);
  nor (_01200_, _01199_, _28260_);
  nor (_01201_, _01198_, _28717_);
  not (_01202_, _01201_);
  nor (_01203_, _01202_, _28780_);
  nor (_01204_, _01203_, _01200_);
  nor (_01205_, _01204_, _01165_);
  not (_01206_, _01204_);
  nor (_01207_, _01206_, _01164_);
  nor (_01208_, _01207_, _01205_);
  not (_01209_, _01208_);
  nor (_01210_, _01160_, _26749_);
  not (_01211_, _01210_);
  not (_01212_, _01166_);
  nor (_01213_, _01172_, _26304_);
  nor (_01214_, _01213_, _25601_);
  not (_01215_, _01183_);
  nor (_01216_, _01215_, _01145_);
  nor (_01217_, _25892_, _26244_);
  nor (_01218_, _29189_, _26237_);
  not (_01219_, _01218_);
  nor (_01220_, _01219_, _01217_);
  nand (_01221_, _01220_, _01216_);
  nor (_01222_, _01221_, _01169_);
  nor (_01223_, _01222_, _25601_);
  nor (_01225_, _01223_, _01214_);
  nand (_01227_, _01225_, _01212_);
  nand (_01228_, _01227_, _28718_);
  not (_01230_, _01228_);
  nor (_01231_, _01230_, _28844_);
  nor (_01233_, _01231_, _01211_);
  not (_01235_, _01231_);
  nor (_01236_, _01235_, _01210_);
  nor (_01237_, _01236_, _01233_);
  nor (_01239_, _01160_, _26642_);
  not (_01240_, _01239_);
  nor (_01241_, _01230_, _28780_);
  nor (_01242_, _01241_, _01240_);
  nor (_01243_, _01160_, _26679_);
  nor (_01244_, _01230_, _28905_);
  not (_01245_, _01244_);
  nand (_01246_, _01245_, _01243_);
  not (_01247_, _01246_);
  nor (_01248_, _01247_, _01242_);
  nand (_01250_, _01248_, _01237_);
  nor (_01251_, _01250_, _01209_);
  nor (_01253_, _01161_, _26677_);
  nor (_01254_, _29267_, _30308_);
  nor (_01255_, _01254_, _01253_);
  not (_01256_, _01255_);
  nor (_01257_, _01199_, _29057_);
  nor (_01258_, _01202_, _29089_);
  nor (_01260_, _01258_, _01257_);
  nor (_01261_, _01260_, _01256_);
  not (_01262_, _01260_);
  nor (_01264_, _01262_, _01255_);
  nor (_01266_, _01264_, _01261_);
  nor (_01267_, _01161_, _26749_);
  nor (_01269_, _01160_, _27726_);
  nor (_01270_, _01269_, _01267_);
  not (_01271_, _01270_);
  nor (_01272_, _01230_, _28971_);
  nor (_01273_, _01228_, _28845_);
  nor (_01274_, _01273_, _01272_);
  not (_01275_, _01274_);
  nor (_01276_, _01275_, _01271_);
  nor (_01277_, _01274_, _01270_);
  nor (_01278_, _01277_, _01276_);
  nand (_01279_, _01278_, _01266_);
  nor (_01280_, _01161_, _27726_);
  nor (_01283_, _26884_, _30308_);
  nor (_01285_, _01283_, _01280_);
  not (_01286_, _01285_);
  nor (_01288_, _01199_, _29053_);
  nor (_01289_, _01202_, _28970_);
  nor (_01290_, _01289_, _01288_);
  nor (_01292_, _01290_, _01286_);
  nand (_01293_, _01198_, _28028_);
  nand (_01294_, _01201_, _28971_);
  nand (_01296_, _01294_, _01293_);
  nor (_01297_, _01296_, _01285_);
  nor (_01298_, _01297_, _01292_);
  nor (_01300_, _01245_, _01243_);
  nor (_01301_, _26721_, _26779_);
  nor (_01302_, _01301_, _26781_);
  not (_01304_, _01302_);
  nor (_01305_, _01304_, _29255_);
  not (_01306_, _01305_);
  not (_01308_, _01241_);
  nor (_01309_, _01308_, _01239_);
  nor (_01310_, _01309_, _01306_);
  not (_01311_, _01310_);
  nor (_01312_, _01311_, _01300_);
  nand (_01313_, _01312_, _01298_);
  nor (_01314_, _01313_, _01279_);
  nand (_01315_, _01314_, _01251_);
  nor (_23458_, _01315_, _23698_);
  nor (_23499_, _29057_, _23698_);
  nor (_01316_, _25603_, _23698_);
  nand (_01317_, _01316_, _04390_);
  nor (_01318_, _25611_, _30658_);
  not (_01319_, _04390_);
  nor (_01320_, _04945_, _04617_);
  not (_01321_, _01320_);
  nor (_01322_, _01321_, _04950_);
  not (_01323_, _01322_);
  nor (_01324_, _01323_, _04879_);
  not (_01325_, _01324_);
  nor (_01326_, _01325_, _04877_);
  not (_01327_, _01326_);
  nor (_01329_, _01327_, _04956_);
  not (_01330_, _01329_);
  not (_01331_, _04510_);
  nor (_01332_, _01331_, _25639_);
  not (_01333_, _04684_);
  nor (_01334_, _01333_, _25671_);
  not (_01335_, _04680_);
  nor (_01336_, _01335_, _25653_);
  not (_01337_, _01336_);
  nor (_01338_, _04684_, _04412_);
  nor (_01339_, _01338_, _01334_);
  not (_01340_, _01339_);
  nor (_01341_, _01340_, _01337_);
  nor (_01342_, _01341_, _01334_);
  nor (_01343_, _04510_, _04417_);
  nor (_01344_, _01343_, _01332_);
  not (_01346_, _01344_);
  nor (_01347_, _01346_, _01342_);
  nor (_01348_, _01347_, _01332_);
  not (_01349_, _01348_);
  nor (_01350_, _01349_, _01330_);
  not (_01351_, _01350_);
  nor (_01352_, _01351_, _04960_);
  nor (_01353_, _01352_, _01319_);
  nor (_01354_, _01330_, _04960_);
  nand (_01355_, _01354_, _01319_);
  nor (_01356_, _01355_, _01349_);
  nor (_01357_, _01356_, _01353_);
  not (_01358_, _04960_);
  nor (_01359_, _01350_, _01358_);
  nor (_01360_, _01359_, _01352_);
  not (_01361_, _01360_);
  nor (_01362_, _01349_, _01327_);
  not (_01363_, _04877_);
  nor (_01364_, _01349_, _01325_);
  nor (_01365_, _01364_, _01363_);
  nor (_01366_, _01365_, _01362_);
  not (_01367_, _01366_);
  not (_01368_, _04879_);
  nor (_01370_, _01349_, _01323_);
  nor (_01372_, _01370_, _01368_);
  nor (_01373_, _01372_, _01364_);
  not (_01375_, _04950_);
  nor (_01376_, _01349_, _01321_);
  nor (_01377_, _01376_, _01375_);
  nor (_01378_, _01377_, _01370_);
  not (_01379_, _01378_);
  nor (_01380_, _01349_, _04945_);
  not (_01381_, _04945_);
  nor (_01382_, _01348_, _01381_);
  nor (_01384_, _01382_, _01380_);
  not (_01385_, _01384_);
  nor (_01386_, _26059_, _26001_);
  not (_01387_, _01386_);
  nor (_01388_, _01387_, _26118_);
  not (_01390_, _01388_);
  nor (_01391_, _01390_, _25938_);
  not (_01392_, _01391_);
  nor (_01393_, _25817_, _25759_);
  not (_01394_, _01393_);
  nor (_01395_, _25872_, _25698_);
  not (_01396_, _01395_);
  nor (_01397_, _01396_, _01394_);
  not (_01398_, _01397_);
  nor (_01399_, _01398_, _01392_);
  not (_01400_, _26118_);
  nor (_01401_, _01400_, _25938_);
  nand (_01402_, _01401_, _01386_);
  not (_01403_, _01402_);
  nor (_01404_, _25870_, _25698_);
  not (_01406_, _01404_);
  nor (_01407_, _01406_, _01394_);
  nand (_01408_, _01407_, _01403_);
  not (_01410_, _25698_);
  nor (_01411_, _25872_, _01410_);
  not (_01413_, _01411_);
  nor (_01414_, _01413_, _01394_);
  nand (_01416_, _01414_, _01391_);
  nand (_01417_, _01416_, _01408_);
  nor (_01418_, _01417_, _01399_);
  nor (_01420_, _25817_, _25757_);
  not (_01422_, _01420_);
  nor (_01424_, _01422_, _01406_);
  not (_01425_, _01424_);
  nor (_01426_, _26118_, _25998_);
  nor (_01427_, _01426_, _26059_);
  nor (_01428_, _01427_, _01425_);
  nor (_01429_, _01411_, _01404_);
  nand (_01430_, _01429_, _01393_);
  nor (_01431_, _01430_, _01402_);
  nor (_01433_, _01431_, _01428_);
  nor (_01434_, _01422_, _01396_);
  not (_01435_, _01434_);
  nor (_01436_, _01435_, _01402_);
  nor (_01437_, _01390_, _25936_);
  not (_01438_, _01437_);
  nor (_01439_, _25815_, _25759_);
  not (_01440_, _01439_);
  nor (_01442_, _01440_, _01396_);
  nor (_01443_, _01440_, _01410_);
  nor (_01445_, _01443_, _01442_);
  nor (_01446_, _01445_, _01438_);
  nor (_01448_, _01446_, _01436_);
  nand (_01449_, _01448_, _01433_);
  nor (_01451_, _26059_, _25998_);
  nand (_01452_, _01451_, _26118_);
  nor (_01454_, _01452_, _25936_);
  nor (_01455_, _25815_, _25757_);
  not (_01457_, _01455_);
  nor (_01458_, _01457_, _01396_);
  nand (_01460_, _01458_, _01454_);
  not (_01461_, _01460_);
  nor (_01462_, _01452_, _01425_);
  nor (_01463_, _01462_, _01461_);
  not (_01464_, _01463_);
  not (_01465_, _01454_);
  nor (_01466_, _01422_, _01413_);
  nor (_01467_, _01440_, _01406_);
  nor (_01468_, _01467_, _01466_);
  nor (_01470_, _01468_, _01465_);
  nor (_01472_, _01470_, _01464_);
  not (_01474_, _01472_);
  nor (_01475_, _01474_, _01449_);
  nand (_01477_, _01475_, _01418_);
  not (_01478_, _01442_);
  not (_01480_, _01452_);
  nor (_01481_, _01480_, _01391_);
  nor (_01483_, _01481_, _01478_);
  not (_01484_, _01443_);
  nor (_01486_, _01452_, _25938_);
  nor (_01487_, _01486_, _01391_);
  nor (_01489_, _01487_, _01484_);
  nor (_01490_, _01422_, _01410_);
  nor (_01491_, _01490_, _01467_);
  nor (_01492_, _01491_, _01427_);
  nor (_01493_, _01492_, _01489_);
  not (_01494_, _01493_);
  nor (_01495_, _01494_, _01483_);
  not (_01496_, _01495_);
  nor (_01497_, _01440_, _01402_);
  not (_01498_, _01486_);
  not (_01499_, _01467_);
  nor (_01500_, _01499_, _01498_);
  nor (_01501_, _01500_, _01497_);
  nor (_01502_, _01440_, _01413_);
  nor (_01503_, _01457_, _25870_);
  nor (_01504_, _01503_, _01502_);
  nor (_01505_, _01504_, _01465_);
  nor (_01506_, _01457_, _25872_);
  nor (_01507_, _01490_, _01506_);
  nor (_01508_, _01507_, _01402_);
  nor (_01509_, _01508_, _01505_);
  nand (_01510_, _01509_, _01501_);
  nor (_01511_, _01400_, _25936_);
  nand (_01512_, _01511_, _01386_);
  nand (_01513_, _01458_, _26059_);
  nand (_01514_, _01513_, _01512_);
  nor (_01515_, _01425_, _01402_);
  nor (_01516_, _01394_, _25870_);
  not (_01517_, _01516_);
  nor (_01519_, _01452_, _01517_);
  nor (_01520_, _01452_, _01435_);
  nor (_01521_, _01520_, _01519_);
  not (_01522_, _01521_);
  nor (_01523_, _01522_, _01515_);
  not (_01524_, _01523_);
  nor (_01525_, _01524_, _01514_);
  not (_01526_, _01525_);
  nor (_01527_, _01526_, _01510_);
  nand (_01528_, _25872_, _25817_);
  nor (_01529_, _01528_, _25759_);
  nor (_01530_, _01529_, _01506_);
  nor (_01531_, _01392_, _25698_);
  nor (_01532_, _01465_, _01410_);
  nor (_01533_, _01532_, _01531_);
  nor (_01534_, _01533_, _01530_);
  nor (_01535_, _01394_, _25872_);
  nand (_01536_, _01454_, _01535_);
  nand (_01537_, _01429_, _01420_);
  nor (_01538_, _01537_, _01392_);
  nor (_01539_, _01413_, _25757_);
  nor (_01540_, _01539_, _01424_);
  nor (_01541_, _01540_, _01392_);
  nor (_01542_, _01541_, _01538_);
  nand (_01543_, _01542_, _01536_);
  nor (_01544_, _01543_, _01534_);
  nand (_01545_, _01544_, _01527_);
  nor (_01546_, _01545_, _01496_);
  not (_01547_, _01546_);
  nor (_01548_, _01547_, _01477_);
  nor (_01549_, _01339_, _01336_);
  nor (_01550_, _01549_, _01341_);
  not (_01551_, _01550_);
  nor (_01552_, _01551_, _01548_);
  nor (_01553_, _04680_, _04414_);
  nor (_01554_, _01553_, _01336_);
  not (_01555_, _01554_);
  nor (_01556_, _01555_, _01547_);
  not (_01557_, _01548_);
  nor (_01558_, _01550_, _01557_);
  nor (_01560_, _01558_, _01552_);
  nand (_01561_, _01560_, _01556_);
  not (_01562_, _01561_);
  nor (_01563_, _01562_, _01552_);
  nand (_01564_, _01346_, _01342_);
  not (_01565_, _01564_);
  nor (_01566_, _01565_, _01347_);
  not (_01567_, _01566_);
  nor (_01568_, _01567_, _01563_);
  nand (_01569_, _01568_, _01385_);
  not (_01570_, _04617_);
  nor (_01571_, _01380_, _01570_);
  nor (_01572_, _01571_, _01376_);
  nor (_01573_, _01572_, _01569_);
  nand (_01574_, _01573_, _01379_);
  nor (_01575_, _01574_, _01373_);
  nand (_01576_, _01575_, _01367_);
  not (_01577_, _04956_);
  nor (_01578_, _01362_, _01577_);
  nor (_01579_, _01578_, _01350_);
  nor (_01580_, _01579_, _01576_);
  nand (_01581_, _01580_, _01361_);
  nor (_01582_, _01581_, _01357_);
  not (_01583_, _01582_);
  nand (_01584_, _01581_, _01357_);
  nand (_01586_, _01584_, _01583_);
  nand (_01587_, _01586_, _01318_);
  nor (_01588_, _01318_, _03078_);
  nor (_01590_, _04344_, _23698_);
  not (_01591_, _01590_);
  nor (_01592_, _01591_, _01588_);
  nand (_01593_, _01592_, _01587_);
  nand (_23540_, _01593_, _01317_);
  nand (_01594_, _01316_, _04960_);
  not (_01595_, _01580_);
  nand (_01596_, _01595_, _01360_);
  nand (_01598_, _01596_, _01581_);
  nand (_01599_, _01598_, _01318_);
  nor (_01600_, _01318_, _03076_);
  nor (_01601_, _01600_, _01591_);
  nand (_01603_, _01601_, _01599_);
  nand (_23581_, _01603_, _01594_);
  nand (_01604_, _01316_, _04956_);
  nand (_01605_, _01579_, _01576_);
  nand (_01607_, _01605_, _01595_);
  nand (_01608_, _01607_, _01318_);
  nor (_01610_, _01318_, _03074_);
  nor (_01611_, _01610_, _01591_);
  nand (_01612_, _01611_, _01608_);
  nand (_23622_, _01612_, _01604_);
  not (_01613_, _01575_);
  nand (_01614_, _01613_, _01366_);
  nand (_01615_, _01614_, _01576_);
  nand (_01616_, _01615_, _01318_);
  nor (_01618_, _01318_, _03131_);
  nor (_01619_, _01618_, _01591_);
  nand (_01621_, _01619_, _01616_);
  nand (_01622_, _01316_, _04877_);
  nand (_23663_, _01622_, _01621_);
  nand (_01623_, _01316_, _04879_);
  nand (_01624_, _01574_, _01373_);
  nand (_01625_, _01624_, _01613_);
  nand (_01626_, _01625_, _01318_);
  nor (_01628_, _01318_, _03122_);
  nor (_01629_, _01628_, _01591_);
  nand (_01630_, _01629_, _01626_);
  nand (_23685_, _01630_, _01623_);
  nand (_01631_, _01316_, _04950_);
  not (_01632_, _01573_);
  nand (_01633_, _01632_, _01378_);
  nand (_01634_, _01633_, _01574_);
  nand (_01635_, _01634_, _01318_);
  nor (_01636_, _01318_, _03119_);
  nor (_01637_, _01636_, _01591_);
  nand (_01638_, _01637_, _01635_);
  nand (_23700_, _01638_, _01631_);
  nand (_01639_, _01572_, _01569_);
  nand (_01640_, _01639_, _01632_);
  nand (_01641_, _01640_, _01318_);
  nor (_01642_, _01318_, _03188_);
  nor (_01644_, _01642_, _01591_);
  nand (_01645_, _01644_, _01641_);
  nand (_01646_, _01316_, _04617_);
  nand (_23741_, _01646_, _01645_);
  nand (_01647_, _01316_, _04945_);
  not (_01648_, _01568_);
  nand (_01649_, _01648_, _01384_);
  nand (_01650_, _01649_, _01569_);
  nand (_01651_, _01650_, _01318_);
  nor (_01652_, _01318_, _03128_);
  nor (_01653_, _01652_, _01591_);
  nand (_01654_, _01653_, _01651_);
  nand (_23782_, _01654_, _01647_);
  nand (_01655_, _01567_, _01563_);
  nand (_01656_, _01655_, _01648_);
  nand (_01657_, _01656_, _01318_);
  nor (_01658_, _01318_, _03301_);
  nor (_01659_, _01658_, _01591_);
  nand (_01660_, _01659_, _01657_);
  nand (_01661_, _01316_, _04510_);
  nand (_23823_, _01661_, _01660_);
  nand (_01662_, _01316_, _04684_);
  not (_01663_, _01318_);
  nor (_01664_, _01560_, _01556_);
  nor (_01665_, _01664_, _01562_);
  nor (_01666_, _01665_, _01663_);
  nor (_01667_, _01318_, _03299_);
  nor (_01668_, _01667_, _01666_);
  nand (_01669_, _01668_, _01590_);
  nand (_23864_, _01669_, _01662_);
  not (_01670_, _01556_);
  nand (_01671_, _01555_, _01547_);
  nand (_01672_, _01671_, _01670_);
  nand (_01673_, _01672_, _01318_);
  nor (_01674_, _01318_, _03297_);
  nor (_01675_, _01674_, _01591_);
  nand (_01676_, _01675_, _01673_);
  nand (_01677_, _01316_, _04680_);
  nand (_23905_, _01677_, _01676_);
  not (_01679_, _26171_);
  nand (_01681_, _26434_, _26329_);
  nor (_01682_, _25888_, _25706_);
  nand (_01683_, _26314_, _29171_);
  nand (_01684_, _01683_, _01682_);
  nand (_01685_, _01684_, _01681_);
  nor (_01686_, _29168_, _26266_);
  nor (_01687_, _01686_, _01685_);
  nand (_01688_, _01687_, _01213_);
  nand (_01689_, _01688_, _01679_);
  nor (_01690_, _26292_, _26244_);
  nand (_01691_, _01690_, _25599_);
  nand (_01692_, _26179_, _25599_);
  nor (_01693_, _01692_, _26286_);
  nor (_01694_, _01693_, _26472_);
  nand (_01695_, _01694_, _01691_);
  not (_01696_, _01695_);
  nand (_01697_, _01696_, _01689_);
  nor (_01698_, _25609_, _26713_);
  not (_01699_, _04514_);
  nor (_01700_, _25712_, _01699_);
  not (_01701_, _04658_);
  nor (_01702_, _25643_, _01701_);
  nor (_01704_, _25657_, _28673_);
  nor (_01705_, _01704_, _01702_);
  not (_01706_, _01705_);
  nor (_01707_, _25631_, _25714_);
  nor (_01708_, _25663_, _28677_);
  nor (_01709_, _01708_, _01707_);
  nor (_01711_, _25621_, _28667_);
  nor (_01712_, _25676_, _25736_);
  nor (_01713_, _01712_, _01711_);
  nand (_01715_, _01713_, _01709_);
  nor (_01716_, _01715_, _01706_);
  nor (_01717_, _01716_, _25684_);
  nor (_01719_, _01717_, _01700_);
  nor (_01720_, _01719_, _25611_);
  nor (_01721_, _01720_, _01698_);
  nand (_01723_, _01721_, _01697_);
  not (_01724_, _01723_);
  nor (_01725_, _01697_, _28684_);
  nor (_01729_, _01725_, _01724_);
  not (_01730_, _01729_);
  nor (_01731_, _01730_, _28266_);
  not (_01732_, _01731_);
  nor (_01733_, _01729_, _03131_);
  nor (_01734_, _01733_, _01731_);
  nand (_01735_, _01682_, _26173_);
  not (_01736_, _01735_);
  not (_01737_, _26290_);
  nor (_01738_, _01186_, _26327_);
  nor (_01739_, _01738_, _01737_);
  nand (_01741_, _01739_, _26306_);
  nor (_01742_, _01741_, _01736_);
  nor (_01743_, _01742_, _26171_);
  nor (_01744_, _01695_, _01743_);
  nor (_01745_, _25609_, _26741_);
  not (_01746_, _05350_);
  nor (_01747_, _25712_, _01746_);
  not (_01748_, _05636_);
  nor (_01749_, _25643_, _01748_);
  nor (_01750_, _25657_, _28829_);
  nor (_01751_, _01750_, _01749_);
  not (_01752_, _01751_);
  nor (_01753_, _25631_, _25771_);
  nor (_01754_, _25663_, _25791_);
  nor (_01755_, _01754_, _01753_);
  nor (_01756_, _25621_, _28823_);
  nor (_01757_, _25676_, _25777_);
  nor (_01758_, _01757_, _01756_);
  nand (_01759_, _01758_, _01755_);
  nor (_01760_, _01759_, _01752_);
  nor (_01761_, _01760_, _25684_);
  nor (_01762_, _01761_, _01747_);
  nor (_01763_, _01762_, _25611_);
  nor (_01764_, _01763_, _01745_);
  not (_01765_, _01764_);
  nor (_01766_, _01765_, _01744_);
  nand (_01767_, _01744_, _28838_);
  not (_01768_, _01767_);
  nor (_01769_, _01768_, _01766_);
  not (_01771_, _01769_);
  nor (_01772_, _01771_, _28407_);
  not (_01773_, _01772_);
  nor (_01774_, _01769_, _03122_);
  nor (_01775_, _01774_, _01772_);
  nor (_01776_, _25609_, _26669_);
  not (_01777_, _05348_);
  nor (_01778_, _25712_, _01777_);
  not (_01779_, _05631_);
  nor (_01780_, _25643_, _01779_);
  nor (_01781_, _25657_, _28882_);
  nor (_01782_, _01781_, _01780_);
  not (_01783_, _01782_);
  nor (_01784_, _25631_, _28877_);
  nor (_01785_, _25663_, _25846_);
  nor (_01786_, _01785_, _01784_);
  nor (_01787_, _25621_, _28875_);
  nor (_01788_, _25676_, _25835_);
  nor (_01789_, _01788_, _01787_);
  nand (_01790_, _01789_, _01786_);
  nor (_01791_, _01790_, _01783_);
  nor (_01792_, _01791_, _25684_);
  nor (_01793_, _01792_, _01778_);
  nor (_01794_, _01793_, _25611_);
  nor (_01795_, _01794_, _01776_);
  not (_01796_, _01795_);
  nor (_01797_, _01796_, _01744_);
  not (_01798_, _28891_);
  nor (_01799_, _01697_, _01798_);
  nor (_01800_, _01799_, _01797_);
  not (_01801_, _01800_);
  nor (_01802_, _01801_, _28347_);
  not (_01803_, _01802_);
  nor (_01804_, _01800_, _03119_);
  nor (_01805_, _01804_, _01802_);
  nor (_01806_, _25609_, _26594_);
  not (_01807_, _05346_);
  nor (_01808_, _25712_, _01807_);
  nor (_01809_, _25631_, _25637_);
  nor (_01810_, _25657_, _25625_);
  nor (_01812_, _01810_, _01809_);
  nor (_01813_, _25621_, _28721_);
  nor (_01814_, _25676_, _25617_);
  nor (_01815_, _01814_, _01813_);
  nand (_01816_, _01815_, _01812_);
  not (_01817_, _05627_);
  nor (_01818_, _25643_, _01817_);
  nor (_01819_, _25663_, _25669_);
  nor (_01820_, _01819_, _01818_);
  not (_01821_, _01820_);
  nor (_01822_, _01821_, _01816_);
  nor (_01823_, _01822_, _25684_);
  nor (_01824_, _01823_, _01808_);
  nor (_01825_, _01824_, _25611_);
  nor (_01826_, _01825_, _01806_);
  not (_01827_, _01826_);
  nor (_01828_, _01827_, _01744_);
  not (_01829_, _28736_);
  nor (_01830_, _01697_, _01829_);
  nor (_01831_, _01830_, _01828_);
  not (_01832_, _01831_);
  nor (_01833_, _01832_, _26929_);
  not (_01834_, _01833_);
  nor (_01835_, _25609_, _26753_);
  not (_01836_, _05344_);
  nor (_01837_, _25712_, _01836_);
  nor (_01838_, _25621_, _28951_);
  nor (_01839_, _25657_, _26017_);
  nor (_01840_, _01839_, _01838_);
  not (_01841_, _01840_);
  not (_01842_, _05623_);
  nor (_01843_, _25643_, _01842_);
  nor (_01844_, _25676_, _26039_);
  nor (_01845_, _01844_, _01843_);
  nor (_01846_, _25663_, _26025_);
  nor (_01847_, _25631_, _28953_);
  nor (_01848_, _01847_, _01846_);
  nand (_01849_, _01848_, _01845_);
  nor (_01850_, _01849_, _01841_);
  nor (_01851_, _01850_, _25684_);
  nor (_01853_, _01851_, _01837_);
  nor (_01854_, _01853_, _25611_);
  nor (_01855_, _01854_, _01835_);
  not (_01856_, _01855_);
  nor (_01857_, _01856_, _01744_);
  nor (_01858_, _01697_, _28967_);
  nor (_01859_, _01858_, _01857_);
  nor (_01860_, _01859_, _03128_);
  not (_01861_, _01859_);
  nor (_01862_, _01861_, _27364_);
  nor (_01863_, _25609_, _26809_);
  not (_01864_, _05342_);
  nor (_01865_, _25712_, _01864_);
  nor (_01867_, _25621_, _29011_);
  nor (_01868_, _25663_, _25966_);
  nor (_01869_, _01868_, _01867_);
  not (_01870_, _01869_);
  not (_01871_, _05618_);
  nor (_01872_, _25643_, _01871_);
  nor (_01873_, _25676_, _25980_);
  nor (_01874_, _01873_, _01872_);
  nor (_01875_, _25657_, _25958_);
  nor (_01876_, _25631_, _29013_);
  nor (_01877_, _01876_, _01875_);
  nand (_01878_, _01877_, _01874_);
  nor (_01879_, _01878_, _01870_);
  nor (_01881_, _01879_, _25684_);
  nor (_01882_, _01881_, _01865_);
  nor (_01883_, _01882_, _25611_);
  nor (_01884_, _01883_, _01863_);
  not (_01885_, _01884_);
  nor (_01886_, _01885_, _01744_);
  not (_01887_, _29027_);
  nor (_01888_, _01697_, _01887_);
  nor (_01889_, _01888_, _01886_);
  not (_01890_, _01889_);
  nor (_01891_, _01890_, _28503_);
  not (_01892_, _01891_);
  nor (_01893_, _25609_, _26844_);
  not (_01894_, _05341_);
  nor (_01896_, _25712_, _01894_);
  nor (_01897_, _25631_, _26098_);
  nor (_01898_, _25657_, _26077_);
  nor (_01899_, _01898_, _01897_);
  nor (_01900_, _25621_, _28032_);
  nor (_01901_, _25676_, _26073_);
  nor (_01902_, _01901_, _01900_);
  nand (_01903_, _01902_, _01899_);
  not (_01905_, _05614_);
  nor (_01906_, _25643_, _01905_);
  nor (_01907_, _25663_, _26084_);
  nor (_01908_, _01907_, _01906_);
  not (_01909_, _01908_);
  nor (_01910_, _01909_, _01903_);
  nor (_01911_, _01910_, _25684_);
  nor (_01912_, _01911_, _01896_);
  nor (_01913_, _01912_, _25611_);
  nor (_01914_, _01913_, _01893_);
  not (_01915_, _01914_);
  nor (_01916_, _01915_, _01744_);
  not (_01917_, _28060_);
  nor (_01918_, _01697_, _01917_);
  nor (_01919_, _01918_, _01916_);
  nand (_01920_, _01919_, _03299_);
  nor (_01921_, _25609_, _26860_);
  not (_01922_, _05339_);
  nor (_01923_, _25712_, _01922_);
  not (_01924_, _05608_);
  nor (_01925_, _25643_, _01924_);
  nor (_01926_, _25657_, _25900_);
  nor (_01927_, _01926_, _01925_);
  not (_01928_, _01927_);
  nor (_01929_, _25631_, _27914_);
  nor (_01930_, _25663_, _25914_);
  nor (_01931_, _01930_, _01929_);
  nor (_01932_, _25621_, _27910_);
  nor (_01933_, _25676_, _25904_);
  nor (_01934_, _01933_, _01932_);
  nand (_01935_, _01934_, _01931_);
  nor (_01936_, _01935_, _01928_);
  nor (_01938_, _01936_, _25684_);
  nor (_01939_, _01938_, _01923_);
  nor (_01940_, _01939_, _25611_);
  nor (_01941_, _01940_, _01921_);
  nand (_01942_, _01941_, _01697_);
  not (_01943_, _27940_);
  nor (_01944_, _01697_, _01943_);
  not (_01945_, _01944_);
  nand (_01946_, _01945_, _01942_);
  nor (_01947_, _01946_, _27231_);
  nand (_01948_, _01914_, _01697_);
  nand (_01949_, _01744_, _28060_);
  nand (_01950_, _01949_, _01948_);
  nor (_01951_, _01950_, _27281_);
  nor (_01952_, _01919_, _03299_);
  nor (_01953_, _01952_, _01951_);
  nand (_01954_, _01953_, _01947_);
  nand (_01955_, _01954_, _01920_);
  nor (_01956_, _01889_, _03301_);
  nor (_01957_, _01956_, _01891_);
  nand (_01958_, _01957_, _01955_);
  nand (_01959_, _01958_, _01892_);
  nor (_01960_, _01959_, _01862_);
  nor (_01961_, _01960_, _01860_);
  nor (_01962_, _01831_, _03188_);
  nor (_01963_, _01962_, _01833_);
  nand (_01964_, _01963_, _01961_);
  nand (_01965_, _01964_, _01834_);
  nand (_01966_, _01965_, _01805_);
  nand (_01967_, _01966_, _01803_);
  nand (_01968_, _01967_, _01775_);
  nand (_01969_, _01968_, _01773_);
  nand (_01970_, _01969_, _01734_);
  nand (_01971_, _01970_, _01732_);
  nand (_01972_, _03076_, _03074_);
  nand (_01973_, _03080_, _03078_);
  nor (_01974_, _01973_, _01972_);
  nand (_01975_, _01974_, _01971_);
  nor (_01976_, _01975_, _26939_);
  nor (_01978_, _01976_, _01729_);
  not (_01980_, _01978_);
  nor (_01982_, _01971_, _03074_);
  nand (_01984_, _01982_, _27306_);
  nand (_01986_, _27368_, _27346_);
  nor (_01987_, _01986_, _01984_);
  nand (_01989_, _01987_, _26939_);
  nand (_01990_, _01989_, _01729_);
  nand (_01992_, _01990_, _01980_);
  nor (_01994_, _01730_, _03083_);
  nor (_01996_, _01729_, _28353_);
  nor (_01997_, _01996_, _01994_);
  nor (_01999_, _01997_, _01992_);
  nor (_02001_, _01999_, _03085_);
  not (_02003_, _26325_);
  nor (_02004_, _02003_, _26173_);
  nor (_02006_, _02004_, _01690_);
  nor (_02007_, _02006_, _25601_);
  not (_02009_, _26146_);
  nor (_02010_, _26126_, _25950_);
  nand (_02011_, _02010_, _26071_);
  nor (_02012_, _02011_, _02009_);
  not (_02013_, _02012_);
  nor (_02014_, _02013_, _26171_);
  nor (_02015_, _02014_, _02007_);
  nor (_02016_, _02015_, _01697_);
  not (_02017_, _01693_);
  nor (_02018_, _26134_, _02009_);
  nor (_02019_, _26199_, _26181_);
  nor (_02020_, _02019_, _02018_);
  not (_02021_, _26191_);
  nand (_02022_, _26420_, _25708_);
  nor (_02023_, _02022_, _29171_);
  nor (_02024_, _02023_, _02021_);
  nand (_02025_, _02024_, _02020_);
  nand (_02026_, _02025_, _01679_);
  nand (_02027_, _02026_, _02017_);
  nor (_02028_, _02027_, _01743_);
  nor (_02029_, _02028_, _02016_);
  nand (_02030_, _01999_, _03085_);
  nand (_02031_, _02030_, _02029_);
  nor (_02033_, _02031_, _02001_);
  nand (_02034_, _31328_, _26472_);
  not (_02035_, _26189_);
  nor (_02036_, _02035_, _26171_);
  nor (_02037_, _02036_, _26308_);
  nor (_02038_, _02037_, _26464_);
  nor (_02039_, _02038_, _26193_);
  nor (_02040_, _02039_, _26193_);
  not (_02041_, _02040_);
  nor (_02042_, _02041_, _00729_);
  not (_02043_, _30067_);
  not (_02044_, _30217_);
  nand (_02045_, _30792_, _30848_);
  nand (_02046_, _30664_, _30489_);
  nor (_02047_, _02046_, _02045_);
  nand (_02048_, _02047_, _30368_);
  nor (_02049_, _02048_, _02044_);
  nand (_02050_, _02049_, _02039_);
  nor (_02051_, _02050_, _02043_);
  nand (_02052_, _02051_, _31214_);
  nor (_02053_, _02041_, _27462_);
  not (_02054_, _02036_);
  nor (_02055_, _02054_, _27095_);
  nor (_02056_, _01728_, _01722_);
  nor (_02057_, _01740_, _01718_);
  nand (_02058_, _02057_, _02056_);
  nor (_02059_, _01703_, _01678_);
  nor (_02060_, _01714_, _01710_);
  nand (_02061_, _02060_, _02059_);
  nor (_02062_, _02061_, _02058_);
  nand (_02063_, _02062_, _26491_);
  not (_02064_, _02063_);
  nor (_02065_, _02064_, _02055_);
  not (_02066_, _02065_);
  nor (_02067_, _02066_, _02053_);
  nand (_02068_, _02067_, _02052_);
  not (_02069_, _02068_);
  nor (_02070_, _01686_, _26304_);
  not (_02071_, _02070_);
  nor (_02072_, _02071_, _02023_);
  nor (_02074_, _26272_, _26146_);
  nor (_02075_, _02074_, _26181_);
  nor (_02076_, _02075_, _01685_);
  nand (_02077_, _02076_, _02072_);
  nand (_02078_, _02077_, _02069_);
  not (_02079_, _02078_);
  nand (_02080_, _02020_, _26432_);
  nor (_02081_, _02080_, _02079_);
  nand (_02082_, _29164_, _26248_);
  nand (_02083_, _02082_, _26179_);
  nand (_02084_, _02083_, _01173_);
  nand (_02085_, _02084_, _02068_);
  nand (_02086_, _02085_, _02081_);
  nand (_02087_, _02086_, _01679_);
  nor (_02088_, _02007_, _26472_);
  nand (_02089_, _02088_, _02087_);
  not (_02090_, _02089_);
  not (_02092_, _29242_);
  nor (_02094_, _02092_, _26901_);
  nor (_02095_, _26749_, _26679_);
  not (_02097_, _02095_);
  nor (_02098_, _02097_, _29297_);
  nand (_02099_, _02098_, _00783_);
  nand (_02100_, _02099_, _02094_);
  nand (_02101_, _02100_, _02036_);
  nor (_02102_, _31406_, _29287_);
  nand (_02103_, _02102_, _30889_);
  nand (_02104_, _02103_, _26491_);
  nand (_02105_, _02104_, _02101_);
  nor (_02106_, _02105_, _02090_);
  nand (_02107_, _02106_, _29285_);
  nor (_02108_, _02107_, _02042_);
  not (_02109_, _02108_);
  not (_02110_, _02018_);
  nor (_02111_, _02110_, _26171_);
  nand (_02112_, _02111_, _31174_);
  not (_02113_, _04449_);
  nor (_02114_, _26126_, _26011_);
  nor (_02115_, _26069_, _25950_);
  nand (_02116_, _02115_, _02114_);
  nor (_02118_, _02116_, _02009_);
  not (_02119_, _02118_);
  nor (_02120_, _02119_, _26171_);
  nand (_02121_, _29172_, _26420_);
  nand (_02122_, _02121_, _26489_);
  nor (_02123_, _02019_, _02118_);
  nand (_02124_, _02123_, _02035_);
  nor (_02125_, _02124_, _02122_);
  nor (_02126_, _02125_, _26171_);
  nand (_02127_, _02017_, _01689_);
  nor (_02128_, _02127_, _02126_);
  nor (_02129_, _02128_, _02016_);
  nor (_02130_, _02129_, _26472_);
  nand (_02131_, _02130_, _01691_);
  nor (_02132_, _02131_, _02120_);
  not (_02133_, _02132_);
  nor (_02134_, _02133_, _02113_);
  nor (_02135_, _01691_, _28838_);
  nor (_02136_, _02135_, _02134_);
  nand (_02137_, _02136_, _02112_);
  nor (_02138_, _02137_, _02109_);
  nand (_02139_, _02138_, _02034_);
  nor (_02140_, _02139_, _02033_);
  not (_02141_, _04868_);
  not (_02142_, _04861_);
  not (_02143_, _04388_);
  nand (_02144_, _25627_, _25639_);
  nand (_02145_, _02144_, _25609_);
  nand (_02146_, _02145_, _25603_);
  not (_02147_, _02146_);
  nor (_02148_, _02147_, _01331_);
  not (_02149_, _02148_);
  nor (_02150_, _02149_, _01381_);
  not (_02151_, _02150_);
  nor (_02152_, _02151_, _01570_);
  not (_02153_, _02152_);
  nor (_02154_, _02153_, _01375_);
  not (_02155_, _02154_);
  nor (_02156_, _02155_, _01368_);
  not (_02157_, _02156_);
  nor (_02161_, _02157_, _01363_);
  not (_02162_, _02161_);
  nor (_02163_, _02162_, _01577_);
  not (_02164_, _02163_);
  nor (_02165_, _02164_, _01358_);
  not (_02166_, _02165_);
  nor (_02167_, _02166_, _01319_);
  not (_02168_, _02167_);
  nor (_02169_, _02168_, _02143_);
  not (_02170_, _02169_);
  nor (_02171_, _02170_, _02142_);
  not (_02172_, _02171_);
  nor (_02173_, _02172_, _02141_);
  not (_02174_, _02173_);
  nor (_02175_, _02174_, _02113_);
  not (_02176_, _02175_);
  nand (_02177_, _02174_, _02113_);
  nand (_02178_, _02177_, _02176_);
  nand (_02179_, _02178_, _02109_);
  nand (_02180_, _02179_, _29344_);
  nor (_23946_, _02180_, _02140_);
  not (_02181_, _02029_);
  not (_02182_, _01992_);
  nor (_02183_, _02182_, _28353_);
  nor (_02184_, _01992_, _03083_);
  nor (_02185_, _02184_, _02183_);
  nor (_02186_, _02185_, _02181_);
  nand (_02187_, _31067_, _26472_);
  not (_02188_, _02111_);
  nor (_02189_, _02188_, _31124_);
  nand (_02190_, _02132_, _04868_);
  not (_02191_, _01691_);
  nand (_02192_, _02191_, _01798_);
  nand (_02193_, _02192_, _02190_);
  nor (_02194_, _02193_, _02189_);
  nand (_02195_, _02194_, _02187_);
  nor (_02196_, _02195_, _02186_);
  nor (_02197_, _02196_, _02109_);
  nand (_02198_, _02172_, _02141_);
  nand (_02199_, _02198_, _02174_);
  nor (_02201_, _02199_, _02108_);
  nor (_02202_, _02201_, _02197_);
  nor (_23987_, _02202_, _23698_);
  nor (_02203_, _01975_, _03082_);
  not (_02204_, _01975_);
  nor (_02205_, _02204_, _26939_);
  nor (_02206_, _02205_, _02203_);
  nor (_02207_, _02206_, _01729_);
  not (_02208_, _01989_);
  nor (_02209_, _01987_, _26939_);
  nor (_02210_, _02209_, _02208_);
  nor (_02211_, _02210_, _01730_);
  nor (_02213_, _02211_, _02207_);
  nor (_02215_, _02213_, _02181_);
  not (_02217_, _30395_);
  nand (_02219_, _02217_, _26472_);
  not (_02221_, _31059_);
  nor (_02223_, _02188_, _02221_);
  nand (_02225_, _02132_, _04861_);
  nand (_02226_, _02191_, _01829_);
  nand (_02227_, _02226_, _02225_);
  nor (_02228_, _02227_, _02223_);
  nand (_02229_, _02228_, _02219_);
  nor (_02230_, _02229_, _02215_);
  nor (_02231_, _02230_, _02109_);
  nand (_02232_, _02170_, _02142_);
  nand (_02233_, _02232_, _02172_);
  nor (_02234_, _02233_, _02108_);
  nor (_02235_, _02234_, _02231_);
  nor (_24028_, _02235_, _23698_);
  not (_02236_, _01734_);
  not (_02237_, _01775_);
  not (_02238_, _01805_);
  not (_02239_, _01942_);
  nor (_02240_, _01944_, _02239_);
  nand (_02241_, _02240_, _03297_);
  nand (_02242_, _01950_, _27281_);
  nand (_02243_, _02242_, _01920_);
  nor (_02244_, _02243_, _02241_);
  nor (_02245_, _02244_, _01951_);
  not (_02247_, _01957_);
  nor (_02248_, _02247_, _02245_);
  nor (_02249_, _02248_, _01891_);
  nor (_02250_, _02249_, _01860_);
  nor (_02251_, _02250_, _01862_);
  not (_02252_, _01963_);
  nor (_02253_, _02252_, _02251_);
  nor (_02254_, _02253_, _01833_);
  nor (_02255_, _02254_, _02238_);
  nor (_02256_, _02255_, _01802_);
  nor (_02257_, _02256_, _02237_);
  nor (_02258_, _02257_, _01772_);
  nor (_02259_, _02258_, _02236_);
  nor (_02260_, _02259_, _01731_);
  nor (_02261_, _01972_, _02260_);
  nand (_02262_, _02261_, _03078_);
  nand (_02263_, _02262_, _01730_);
  not (_02264_, _02263_);
  nor (_02265_, _01984_, _03078_);
  nor (_02266_, _02265_, _01730_);
  nor (_02267_, _02266_, _02264_);
  nor (_02268_, _02267_, _27368_);
  not (_02269_, _02267_);
  nor (_02270_, _02269_, _03080_);
  nor (_02271_, _02270_, _02268_);
  nor (_02272_, _02271_, _02181_);
  nand (_02273_, _00164_, _26472_);
  nor (_02274_, _02188_, _00146_);
  nand (_02275_, _02132_, _04388_);
  nand (_02276_, _02191_, _28967_);
  nand (_02277_, _02276_, _02275_);
  nor (_02278_, _02277_, _02274_);
  nand (_02279_, _02278_, _02273_);
  nor (_02280_, _02279_, _02272_);
  nor (_02281_, _02280_, _02109_);
  nand (_02282_, _02168_, _02143_);
  nand (_02283_, _02282_, _02170_);
  nor (_02284_, _02283_, _02108_);
  nor (_02285_, _02284_, _02281_);
  nor (_24069_, _02285_, _23698_);
  nand (_02287_, _02132_, _02007_);
  nor (_02288_, _02287_, _25757_);
  nand (_02289_, _30692_, _26472_);
  not (_02290_, _02287_);
  nor (_02291_, _02290_, _02131_);
  not (_02292_, _02291_);
  nor (_02293_, _02292_, _02014_);
  nand (_02294_, _02293_, _04390_);
  nand (_02295_, _02191_, _01887_);
  nand (_02296_, _02295_, _02294_);
  not (_02297_, _02120_);
  nor (_02298_, _02297_, _00088_);
  nor (_02299_, _02298_, _02296_);
  nand (_02300_, _02299_, _02289_);
  nor (_02301_, _02300_, _02288_);
  nand (_02302_, _02260_, _27227_);
  nor (_02303_, _02302_, _03076_);
  nor (_02304_, _02303_, _01730_);
  nor (_02305_, _02261_, _01729_);
  nor (_02306_, _02305_, _02304_);
  not (_02307_, _02306_);
  nand (_02308_, _02307_, _03078_);
  nand (_02309_, _02306_, _27346_);
  nand (_02310_, _02309_, _02308_);
  nand (_02311_, _02310_, _02029_);
  nand (_02312_, _02311_, _02301_);
  nor (_02313_, _02312_, _02109_);
  nand (_02314_, _02166_, _01319_);
  nand (_02315_, _02314_, _02168_);
  nand (_02316_, _02315_, _02109_);
  nand (_02317_, _02316_, _29344_);
  nor (_24111_, _02317_, _02313_);
  nor (_02318_, _02260_, _27227_);
  nor (_02319_, _02318_, _01729_);
  nor (_02320_, _01982_, _01730_);
  nor (_02321_, _02320_, _02319_);
  nor (_02322_, _02321_, _27306_);
  not (_02323_, _02321_);
  nor (_02324_, _02323_, _03076_);
  nor (_02325_, _02324_, _02322_);
  nor (_02327_, _02325_, _02181_);
  nand (_02328_, _30828_, _26472_);
  nor (_02329_, _02188_, _31396_);
  nand (_02330_, _02290_, _25817_);
  not (_02331_, _02293_);
  nor (_02332_, _02331_, _01358_);
  nor (_02333_, _01691_, _28060_);
  nor (_02334_, _02333_, _02332_);
  nand (_02335_, _02334_, _02330_);
  nor (_02336_, _02335_, _02329_);
  nand (_02337_, _02336_, _02328_);
  nor (_02338_, _02337_, _02327_);
  nor (_02339_, _02338_, _02109_);
  nand (_02340_, _02164_, _01358_);
  nand (_02341_, _02340_, _02166_);
  nor (_02342_, _02341_, _02108_);
  nor (_02343_, _02342_, _02339_);
  nor (_24152_, _02343_, _23698_);
  nand (_02344_, _02162_, _01577_);
  nand (_02345_, _02344_, _02164_);
  nand (_02346_, _02345_, _02109_);
  nand (_02347_, _02346_, _29344_);
  nor (_02348_, _02287_, _25870_);
  nand (_02349_, _31419_, _26472_);
  nand (_02350_, _02293_, _04956_);
  nand (_02351_, _02191_, _01943_);
  nand (_02352_, _02351_, _02350_);
  nor (_02353_, _02297_, _00042_);
  nor (_02354_, _02353_, _02352_);
  nand (_02355_, _02354_, _02349_);
  nor (_02356_, _02355_, _02348_);
  nor (_02357_, _02260_, _03074_);
  nor (_02358_, _01971_, _27227_);
  nor (_02359_, _02358_, _02357_);
  nand (_02360_, _02359_, _01729_);
  nand (_02361_, _02302_, _02319_);
  nand (_02362_, _02361_, _02360_);
  nand (_02363_, _02362_, _02129_);
  nand (_02364_, _02363_, _02356_);
  nor (_02365_, _02364_, _02109_);
  nor (_24193_, _02365_, _02347_);
  nand (_02367_, _02291_, _31253_);
  nor (_02368_, _01969_, _01734_);
  nand (_02369_, _02029_, _01970_);
  nor (_02370_, _02369_, _02368_);
  nand (_02371_, _02290_, _28684_);
  nor (_02372_, _01721_, _01691_);
  nor (_02373_, _26487_, _01363_);
  nor (_02374_, _02373_, _02372_);
  nand (_02375_, _02374_, _02371_);
  nor (_02376_, _02375_, _02370_);
  nand (_02377_, _02376_, _02367_);
  nor (_02378_, _02377_, _02109_);
  nand (_02379_, _02157_, _01363_);
  nand (_02380_, _02379_, _02162_);
  nand (_02381_, _02380_, _02109_);
  nand (_02382_, _02381_, _29344_);
  nor (_24234_, _02382_, _02378_);
  nor (_02383_, _02292_, _30122_);
  nor (_02384_, _02287_, _28838_);
  nand (_02385_, _01765_, _02191_);
  nand (_02386_, _26472_, _04879_);
  nand (_02387_, _02386_, _02385_);
  nor (_02388_, _02387_, _02384_);
  nand (_02389_, _02256_, _02237_);
  nor (_02390_, _02181_, _02257_);
  nand (_02391_, _02390_, _02389_);
  nand (_02392_, _02391_, _02388_);
  nor (_02393_, _02392_, _02383_);
  nor (_02394_, _02393_, _02109_);
  nand (_02395_, _02155_, _01368_);
  nand (_02396_, _02395_, _02157_);
  nor (_02397_, _02396_, _02108_);
  nor (_02398_, _02397_, _02394_);
  nor (_24275_, _02398_, _23698_);
  nor (_02399_, _02292_, _30244_);
  nand (_02400_, _02254_, _02238_);
  nor (_02401_, _02181_, _02255_);
  nand (_02402_, _02401_, _02400_);
  nor (_02403_, _02287_, _28891_);
  nand (_02405_, _01796_, _02191_);
  nand (_02406_, _26472_, _04950_);
  nand (_02407_, _02406_, _02405_);
  nor (_02408_, _02407_, _02403_);
  nand (_02409_, _02408_, _02402_);
  nor (_02410_, _02409_, _02399_);
  nor (_02411_, _02410_, _02109_);
  nand (_02412_, _02153_, _01375_);
  nand (_02413_, _02412_, _02155_);
  nor (_02414_, _02413_, _02108_);
  nor (_02415_, _02414_, _02411_);
  nor (_24316_, _02415_, _23698_);
  nor (_02416_, _02292_, _30395_);
  nor (_02417_, _02287_, _28736_);
  nand (_02418_, _01827_, _02191_);
  nand (_02419_, _26472_, _04617_);
  nand (_02420_, _02419_, _02418_);
  nor (_02421_, _02420_, _02417_);
  nand (_02422_, _02252_, _02251_);
  nor (_02423_, _02181_, _02253_);
  nand (_02424_, _02423_, _02422_);
  nand (_02425_, _02424_, _02421_);
  nor (_02426_, _02425_, _02416_);
  nor (_02427_, _02426_, _02109_);
  nand (_02428_, _02151_, _01570_);
  nand (_02429_, _02428_, _02153_);
  nor (_02430_, _02429_, _02108_);
  nor (_02431_, _02430_, _02427_);
  nor (_24357_, _02431_, _23698_);
  nor (_02432_, _02292_, _30533_);
  nor (_02433_, _02287_, _28966_);
  nand (_02434_, _01856_, _02191_);
  nand (_02435_, _26472_, _04945_);
  nand (_02436_, _02435_, _02434_);
  nor (_02437_, _02436_, _02433_);
  nor (_02438_, _01860_, _01862_);
  nand (_02439_, _02438_, _01959_);
  nor (_02440_, _02438_, _01959_);
  nor (_02441_, _02440_, _02181_);
  nand (_02442_, _02441_, _02439_);
  nand (_02444_, _02442_, _02437_);
  nor (_02445_, _02444_, _02432_);
  nor (_02446_, _02445_, _02109_);
  nor (_02447_, _02148_, _04945_);
  nor (_02448_, _02447_, _02150_);
  not (_02449_, _02448_);
  nor (_02450_, _02449_, _02108_);
  nor (_02451_, _02450_, _02446_);
  nor (_24398_, _02451_, _23698_);
  nor (_02452_, _02146_, _04510_);
  nor (_02453_, _02452_, _02148_);
  nor (_02454_, _02453_, _02108_);
  nor (_02455_, _02292_, _30693_);
  nand (_02456_, _02247_, _02245_);
  nor (_02457_, _02181_, _02248_);
  nand (_02458_, _02457_, _02456_);
  nor (_02459_, _02287_, _29027_);
  nand (_02460_, _01885_, _02191_);
  nand (_02461_, _26472_, _04510_);
  nand (_02462_, _02461_, _02460_);
  nor (_02463_, _02462_, _02459_);
  nand (_02464_, _02463_, _02458_);
  nor (_02465_, _02464_, _02455_);
  nand (_02466_, _02465_, _02108_);
  nand (_02467_, _02466_, _29344_);
  nor (_24439_, _02467_, _02454_);
  nor (_02468_, _02109_, _26472_);
  nor (_02469_, _02468_, _01333_);
  nor (_02470_, _02292_, _30829_);
  nor (_02471_, _01914_, _01691_);
  nor (_02472_, _02287_, _28060_);
  nor (_02473_, _02472_, _02471_);
  nand (_02474_, _02243_, _02241_);
  nor (_02475_, _02181_, _02244_);
  nand (_02476_, _02475_, _02474_);
  nand (_02477_, _02476_, _02473_);
  nor (_02478_, _02477_, _02470_);
  nor (_02479_, _02478_, _02109_);
  nor (_02480_, _02479_, _02469_);
  nor (_24480_, _02480_, _23698_);
  nor (_02482_, _02468_, _01335_);
  nor (_02483_, _02292_, _30876_);
  nand (_02484_, _02290_, _01943_);
  nor (_02485_, _01941_, _01691_);
  nor (_02486_, _02240_, _03297_);
  nand (_02487_, _02029_, _02241_);
  nor (_02488_, _02487_, _02486_);
  nor (_02489_, _02488_, _02485_);
  nand (_02490_, _02489_, _02484_);
  nor (_02491_, _02490_, _02483_);
  nor (_02492_, _02491_, _02109_);
  nor (_02493_, _02492_, _02482_);
  nor (_24522_, _02493_, _23698_);
  nor (_24563_, _28817_, _23698_);
  nor (_24604_, _28872_, _23698_);
  nor (_24645_, _28765_, _23698_);
  nor (_24686_, _28946_, _23698_);
  nor (_24727_, _29008_, _23698_);
  nor (_24768_, _28250_, _23698_);
  nor (_24809_, _27894_, _23698_);
  nor (_24850_, _27722_, _23698_);
  nor (_24891_, _26201_, _23698_);
  nor (_24933_, _26126_, _23698_);
  nor (_24974_, _25950_, _23698_);
  nor (_02494_, _01547_, _25653_);
  nor (_02495_, _01548_, _25671_);
  nor (_02496_, _01557_, _04412_);
  nor (_02497_, _02496_, _02495_);
  nand (_02498_, _02497_, _02494_);
  not (_02499_, _02498_);
  nor (_02500_, _02497_, _02494_);
  nor (_02501_, _02500_, _02499_);
  nor (_02502_, _02501_, _25611_);
  nand (_02503_, _25611_, _25671_);
  nand (_02504_, _02503_, _01590_);
  nor (_25015_, _02504_, _02502_);
  nor (_02505_, _02147_, _25682_);
  nor (_02506_, _02505_, _05413_);
  nand (_02507_, _02505_, _01871_);
  nand (_02508_, _02507_, _29344_);
  nor (_25056_, _02508_, _02506_);
  nor (_02510_, _02505_, _26039_);
  not (_02511_, _04901_);
  not (_02512_, _02505_);
  nor (_02513_, _02512_, _02511_);
  nor (_02514_, _02513_, _02510_);
  nor (_25097_, _02514_, _23698_);
  nor (_02515_, _30316_, _23698_);
  nand (_02516_, _02515_, _06045_);
  nor (_02517_, _02511_, _25682_);
  not (_02518_, _30316_);
  nor (_30303_, _02518_, _23698_);
  nand (_02519_, _30303_, _02517_);
  nand (_25138_, _02519_, _02516_);
  nor (_02520_, _02505_, _05392_);
  nand (_02521_, _02505_, _29011_);
  nand (_02522_, _02521_, _29344_);
  nor (_25179_, _02522_, _02520_);
  nor (_02523_, _02505_, _05608_);
  not (_02524_, _04778_);
  nand (_02525_, _02505_, _02524_);
  nand (_02526_, _02525_, _29344_);
  nor (_25220_, _02526_, _02523_);
  nor (_02527_, _02505_, _05409_);
  nand (_02528_, _02505_, _01905_);
  nand (_02529_, _02528_, _29344_);
  nor (_25261_, _02529_, _02527_);
  nand (_02530_, _02515_, _06040_);
  not (_02531_, _04889_);
  nor (_02532_, _02531_, _25682_);
  nand (_02533_, _02532_, _30303_);
  nand (_25302_, _02533_, _02530_);
  nor (_02534_, _02505_, _05897_);
  nand (_02535_, _02505_, _25904_);
  nand (_02536_, _02535_, _29344_);
  nor (_25344_, _02536_, _02534_);
  nor (_02537_, _02505_, _05618_);
  not (_02538_, _04786_);
  nand (_02539_, _02505_, _02538_);
  nand (_02540_, _02539_, _29344_);
  nor (_25385_, _02540_, _02537_);
  nor (_02543_, _02505_, _05394_);
  nand (_02544_, _02505_, _28951_);
  nand (_02545_, _02544_, _29344_);
  nor (_25426_, _02545_, _02543_);
  nor (_02546_, _02505_, _05900_);
  nand (_02547_, _02505_, _26073_);
  nand (_02548_, _02547_, _29344_);
  nor (_25467_, _02548_, _02546_);
  nor (_02549_, _02505_, _05367_);
  nand (_02550_, _02505_, _28953_);
  nand (_02551_, _02550_, _29344_);
  nor (_25508_, _02551_, _02549_);
  nor (_02552_, _02505_, _05403_);
  nand (_02553_, _02505_, _28875_);
  nand (_02554_, _02553_, _29344_);
  nor (_25549_, _02554_, _02552_);
  not (_02555_, _04814_);
  not (_02556_, _04811_);
  nand (_02557_, _04820_, _04817_);
  not (_02558_, _02557_);
  nor (_02559_, _02558_, _02556_);
  nor (_02560_, _02559_, _02555_);
  not (_02561_, _02559_);
  nor (_02562_, _02561_, _04814_);
  nor (_02563_, _02562_, _02560_);
  nor (_25593_, _02563_, _23698_);
  not (_02564_, _04817_);
  nor (_02565_, _02555_, _02556_);
  not (_02566_, _02565_);
  nor (_02567_, _02566_, _02564_);
  nor (_02568_, _02565_, _04817_);
  nor (_02569_, _02568_, _02567_);
  nor (_02570_, _02569_, _02558_);
  nor (_25674_, _02570_, _23698_);
  nand (_02571_, _02515_, _06047_);
  not (_02572_, _04905_);
  nor (_02573_, _02572_, _25682_);
  nand (_02574_, _02573_, _30303_);
  nand (_25755_, _02574_, _02571_);
  nor (_02576_, _02505_, _05459_);
  not (_02577_, _04736_);
  nand (_02578_, _02505_, _02577_);
  nand (_02579_, _02578_, _29344_);
  nor (_25836_, _02579_, _02576_);
  nand (_02580_, _02515_, _06051_);
  not (_02581_, _04912_);
  nor (_02582_, _02581_, _25682_);
  nand (_02583_, _02582_, _30303_);
  nand (_25918_, _02583_, _02580_);
  nand (_02584_, _02558_, _02556_);
  nand (_02585_, _02584_, _02561_);
  nor (_25999_, _02585_, _23698_);
  nand (_02587_, _00546_, _29344_);
  not (_02588_, _00551_);
  not (_02589_, _00561_);
  nor (_02590_, _00559_, _00556_);
  nand (_02591_, _02590_, _02589_);
  nor (_02592_, _00546_, _00350_);
  nor (_02593_, _00554_, _00549_);
  nand (_02594_, _02593_, _02592_);
  nor (_02595_, _02594_, _02591_);
  nand (_02596_, _02595_, _02588_);
  not (_02597_, _02596_);
  nor (_02598_, _01746_, _23698_);
  nand (_02599_, _02598_, _02597_);
  nand (_26080_, _02599_, _02587_);
  nand (_02600_, _02515_, _06049_);
  not (_02601_, _04908_);
  nor (_02602_, _02601_, _25682_);
  nand (_02603_, _02602_, _30303_);
  nand (_26161_, _02603_, _02600_);
  nor (_02604_, _02505_, _05382_);
  nand (_02605_, _02505_, _25771_);
  nand (_02606_, _02605_, _29344_);
  nor (_26242_, _02606_, _02604_);
  nor (_02607_, _02505_, _05493_);
  not (_02608_, _04768_);
  nand (_02609_, _02505_, _02608_);
  nand (_02610_, _02609_, _29344_);
  nor (_26323_, _02610_, _02607_);
  nand (_02612_, _02515_, _06043_);
  not (_02613_, _04897_);
  nor (_02614_, _02613_, _25682_);
  nand (_02615_, _02614_, _30303_);
  nand (_26404_, _02615_, _02612_);
  nor (_02616_, _02505_, _05355_);
  nand (_02617_, _02505_, _27914_);
  nand (_02618_, _02617_, _29344_);
  nor (_26485_, _02618_, _02616_);
  nor (_02620_, _02505_, _05407_);
  nand (_02621_, _02505_, _01924_);
  nand (_02622_, _02621_, _29344_);
  nor (_26566_, _02622_, _02620_);
  nand (_02623_, _02515_, _06042_);
  not (_02624_, _04893_);
  nor (_02625_, _02624_, _25682_);
  nand (_02626_, _02625_, _30303_);
  nand (_26647_, _02626_, _02623_);
  nor (_02627_, _02505_, _05379_);
  nand (_02628_, _02505_, _28877_);
  nand (_02629_, _02628_, _29344_);
  nor (_26729_, _02629_, _02627_);
  nor (_02630_, _02505_, _05918_);
  nand (_02631_, _02505_, _26039_);
  nand (_02632_, _02631_, _29344_);
  nor (_26810_, _02632_, _02630_);
  nor (_02633_, _02505_, _05915_);
  nand (_02634_, _02505_, _25980_);
  nand (_02635_, _02634_, _29344_);
  nor (_26891_, _02635_, _02633_);
  nor (_02636_, _02505_, _05457_);
  not (_02637_, _04731_);
  nand (_02638_, _02505_, _02637_);
  nand (_02639_, _02638_, _29344_);
  nor (_26972_, _02639_, _02636_);
  nor (_02640_, _02505_, _06067_);
  not (_02641_, _04748_);
  nand (_02642_, _02505_, _02641_);
  nand (_02643_, _02642_, _29344_);
  nor (_27053_, _02643_, _02640_);
  nor (_02645_, _02505_, _05623_);
  not (_02646_, _04790_);
  nand (_02647_, _02505_, _02646_);
  nand (_02648_, _02647_, _29344_);
  nor (_27134_, _02648_, _02645_);
  nor (_02649_, _02505_, _05390_);
  nand (_02650_, _02505_, _28032_);
  nand (_02651_, _02650_, _29344_);
  nor (_27215_, _02651_, _02649_);
  nor (_02653_, _02505_, _05359_);
  nand (_02654_, _02505_, _26098_);
  nand (_02655_, _02654_, _29344_);
  nor (_27296_, _02655_, _02653_);
  nor (_02656_, _02505_, _05388_);
  nand (_02657_, _02505_, _27910_);
  nand (_02658_, _02657_, _29344_);
  nor (_27377_, _02658_, _02656_);
  nor (_02659_, _02505_, _05375_);
  nand (_02660_, _02505_, _25637_);
  nand (_02661_, _02660_, _29344_);
  nor (_27458_, _02661_, _02659_);
  nor (_02662_, _02505_, _05452_);
  not (_02663_, _04720_);
  nand (_02664_, _02505_, _02663_);
  nand (_02665_, _02664_, _29344_);
  nor (_27540_, _02665_, _02662_);
  nor (_02666_, _02505_, _05420_);
  nand (_02667_, _02505_, _01817_);
  nand (_02668_, _02667_, _29344_);
  nor (_27621_, _02668_, _02666_);
  nor (_02669_, _02505_, _06072_);
  not (_02670_, _04774_);
  nand (_02671_, _02505_, _02670_);
  nand (_02672_, _02671_, _29344_);
  nor (_27702_, _02672_, _02669_);
  nor (_02673_, _02505_, _05453_);
  not (_02674_, _04724_);
  nand (_02675_, _02505_, _02674_);
  nand (_02676_, _02675_, _29344_);
  nor (_27783_, _02676_, _02673_);
  nor (_02678_, _02505_, _05455_);
  not (_02679_, _04728_);
  nand (_02680_, _02505_, _02679_);
  nand (_02681_, _02680_, _29344_);
  nor (_27864_, _02681_, _02678_);
  nor (_02682_, _06094_, _06091_);
  nand (_02683_, _02682_, _04696_);
  nor (_02684_, _02683_, _31419_);
  not (_02685_, _04682_);
  nand (_02687_, _02683_, _02685_);
  nand (_02688_, _02687_, _29344_);
  nor (_27945_, _02688_, _02684_);
  nor (_02689_, _01547_, _25611_);
  nand (_02690_, _02689_, _04414_);
  not (_02691_, _02689_);
  nand (_02692_, _02691_, _25653_);
  nand (_02693_, _02692_, _02690_);
  nor (_28026_, _02693_, _01591_);
  nor (_02694_, _02505_, _25736_);
  not (_02695_, _04717_);
  nor (_02696_, _02512_, _02695_);
  nor (_02697_, _02696_, _02694_);
  nor (_28107_, _02697_, _23698_);
  nor (_02698_, _02505_, _05478_);
  not (_02699_, _04761_);
  nand (_02700_, _02505_, _02699_);
  nand (_02701_, _02700_, _29344_);
  nor (_28188_, _02701_, _02698_);
  nor (_02702_, _02505_, _05497_);
  not (_02703_, _04772_);
  nand (_02704_, _02505_, _02703_);
  nand (_02705_, _02704_, _29344_);
  nor (_28269_, _02705_, _02702_);
  nor (_02706_, _02505_, _05415_);
  nand (_02707_, _02505_, _01842_);
  nand (_02708_, _02707_, _29344_);
  nor (_28351_, _02708_, _02706_);
  nor (_02709_, _02505_, _05921_);
  nand (_02710_, _02505_, _25617_);
  nand (_02712_, _02710_, _29344_);
  nor (_28432_, _02712_, _02709_);
  nor (_02713_, _02505_, _05362_);
  nand (_02714_, _02505_, _29013_);
  nand (_02715_, _02714_, _29344_);
  nor (_28487_, _02715_, _02713_);
  nor (_02716_, _02505_, _05614_);
  not (_02717_, _04782_);
  nand (_02718_, _02505_, _02717_);
  nand (_02719_, _02718_, _29344_);
  nor (_28528_, _02719_, _02716_);
  nor (_02720_, _02505_, _25617_);
  nor (_02721_, _02512_, _02572_);
  nor (_02722_, _02721_, _02720_);
  nor (_28569_, _02722_, _23698_);
  nor (_02723_, _02505_, _05631_);
  not (_02724_, _04798_);
  nand (_02725_, _02505_, _02724_);
  nand (_02726_, _02725_, _29344_);
  nor (_28610_, _02726_, _02723_);
  nor (_02727_, _02505_, _06063_);
  nand (_02728_, _02505_, _28667_);
  nand (_02729_, _02728_, _29344_);
  nor (_28651_, _02729_, _02727_);
  nor (_02730_, _02512_, _02601_);
  nor (_02731_, _02505_, _25835_);
  nor (_02732_, _02731_, _02730_);
  nor (_28692_, _02732_, _23698_);
  nor (_02733_, _02505_, _05627_);
  not (_02734_, _04794_);
  nand (_02735_, _02505_, _02734_);
  nand (_02736_, _02735_, _29344_);
  nor (_28733_, _02736_, _02733_);
  nor (_02737_, _02505_, _05636_);
  not (_02738_, _04801_);
  nand (_02739_, _02505_, _02738_);
  nand (_02740_, _02739_, _29344_);
  nor (_28774_, _02740_, _02737_);
  nor (_02741_, _02596_, _01807_);
  nor (_02742_, _02741_, _00551_);
  nor (_28816_, _02742_, _23698_);
  nor (_02744_, _02505_, _26073_);
  nor (_02745_, _02512_, _02624_);
  nor (_02746_, _02745_, _02744_);
  nor (_28857_, _02746_, _23698_);
  nor (_02747_, _02505_, _25980_);
  nor (_02748_, _02512_, _02613_);
  nor (_02749_, _02748_, _02747_);
  nor (_28898_, _02749_, _23698_);
  nor (_02750_, _02512_, _02531_);
  nor (_02751_, _02505_, _25904_);
  nor (_02752_, _02751_, _02750_);
  nor (_28939_, _02752_, _23698_);
  nor (_02753_, _02596_, _01777_);
  nor (_02754_, _02753_, _00549_);
  nor (_28980_, _02754_, _23698_);
  nor (_02755_, _02505_, _05427_);
  nand (_02756_, _02505_, _01748_);
  nand (_02757_, _02756_, _29344_);
  nor (_29021_, _02757_, _02755_);
  nor (_02758_, _02505_, _05472_);
  not (_02759_, _04757_);
  nand (_02760_, _02505_, _02759_);
  nand (_02761_, _02760_, _29344_);
  nor (_29062_, _02761_, _02758_);
  nor (_02762_, _02505_, _05422_);
  nand (_02763_, _02505_, _01779_);
  nand (_02764_, _02763_, _29344_);
  nor (_29103_, _02764_, _02762_);
  nor (_02765_, _02683_, _30828_);
  not (_02766_, _04686_);
  nand (_02767_, _02683_, _02766_);
  nand (_02768_, _02767_, _29344_);
  nor (_29144_, _02768_, _02765_);
  nor (_02769_, _02683_, _00164_);
  not (_02770_, _04693_);
  nand (_02771_, _02683_, _02770_);
  nand (_02772_, _02771_, _29344_);
  nor (_29185_, _02772_, _02769_);
  nor (_02773_, _01355_, _04388_);
  not (_02775_, _02773_);
  nor (_02776_, _02775_, _01349_);
  nor (_02777_, _02776_, _02142_);
  nor (_02778_, _02775_, _04861_);
  not (_02779_, _02778_);
  nor (_02780_, _02779_, _01349_);
  nor (_02781_, _02780_, _02777_);
  nor (_02782_, _01356_, _02143_);
  nor (_02783_, _02782_, _02776_);
  not (_02784_, _02783_);
  nand (_02785_, _02784_, _01582_);
  nor (_02786_, _02785_, _02781_);
  not (_02787_, _02786_);
  nand (_02788_, _02785_, _02781_);
  nand (_02789_, _02788_, _02787_);
  nand (_02790_, _02789_, _01318_);
  nor (_02791_, _01318_, _03082_);
  nor (_02792_, _02791_, _01591_);
  nand (_02793_, _02792_, _02790_);
  nand (_02794_, _01316_, _04861_);
  nand (_29228_, _02794_, _02793_);
  nor (_02795_, _02780_, _02141_);
  nor (_02796_, _02779_, _04868_);
  nand (_02797_, _02796_, _01348_);
  not (_02798_, _02797_);
  nor (_02799_, _02798_, _02795_);
  not (_02800_, _02799_);
  nand (_02801_, _02800_, _02786_);
  nand (_02802_, _02799_, _02787_);
  nand (_02803_, _02802_, _02801_);
  nand (_02804_, _02803_, _01318_);
  nor (_02805_, _01318_, _03083_);
  nor (_02806_, _02805_, _01591_);
  nand (_02807_, _02806_, _02804_);
  nand (_02808_, _01316_, _04868_);
  nand (_29269_, _02808_, _02807_);
  nor (_02810_, _02798_, _02113_);
  nor (_02811_, _02797_, _04449_);
  nor (_02812_, _02811_, _02810_);
  nor (_02813_, _02812_, _02801_);
  not (_02815_, _02813_);
  nand (_02816_, _02812_, _02801_);
  nand (_02817_, _02816_, _02815_);
  nand (_02818_, _02817_, _01318_);
  nor (_02819_, _01318_, _03085_);
  nor (_02820_, _02819_, _01591_);
  nand (_02821_, _02820_, _02818_);
  nand (_02822_, _01316_, _04449_);
  nand (_29311_, _02822_, _02821_);
  nor (_02823_, _02596_, _01922_);
  nor (_02824_, _02823_, _00561_);
  nor (_29352_, _02824_, _23698_);
  nor (_02825_, _02596_, _01894_);
  nor (_02826_, _02825_, _00559_);
  nor (_29393_, _02826_, _23698_);
  nor (_02827_, _02596_, _01836_);
  nor (_02828_, _02827_, _00554_);
  nor (_29434_, _02828_, _23698_);
  nand (_02829_, _00556_, _29344_);
  nor (_02830_, _01864_, _23698_);
  nand (_02831_, _02830_, _02597_);
  nand (_29475_, _02831_, _02829_);
  nor (_02832_, _02505_, _06061_);
  nand (_02833_, _02505_, _25714_);
  nand (_02834_, _02833_, _29344_);
  nor (_29516_, _02834_, _02832_);
  nor (_02835_, _02505_, _25777_);
  nor (_02836_, _02512_, _02581_);
  nor (_02837_, _02836_, _02835_);
  nor (_29557_, _02837_, _23698_);
  nor (_02838_, _02505_, _05405_);
  nand (_02839_, _02505_, _28823_);
  nand (_02840_, _02839_, _29344_);
  nor (_29598_, _02840_, _02838_);
  nor (_02841_, _02505_, _05468_);
  not (_02842_, _04754_);
  nand (_02843_, _02505_, _02842_);
  nand (_02844_, _02843_, _29344_);
  nor (_29640_, _02844_, _02841_);
  nor (_02845_, _02505_, _05464_);
  not (_02847_, _04751_);
  nand (_02848_, _02505_, _02847_);
  nand (_02849_, _02848_, _29344_);
  nor (_29681_, _02849_, _02845_);
  nor (_02850_, _02505_, _04349_);
  not (_02851_, _04744_);
  nand (_02852_, _02505_, _02851_);
  nand (_02853_, _02852_, _29344_);
  nor (_29722_, _02853_, _02850_);
  nor (_02854_, _02683_, _30692_);
  not (_02856_, _04689_);
  nand (_02857_, _02683_, _02856_);
  nand (_02858_, _02857_, _29344_);
  nor (_29763_, _02858_, _02854_);
  nor (_02859_, _02505_, _05398_);
  nand (_02860_, _02505_, _28721_);
  nand (_02861_, _02860_, _29344_);
  nor (_29804_, _02861_, _02859_);
  nor (_02862_, _02505_, _05491_);
  not (_02863_, _04764_);
  nand (_02864_, _02505_, _02863_);
  nand (_02865_, _02864_, _29344_);
  nor (_29845_, _02865_, _02862_);
  nor (_02866_, _02505_, _06059_);
  nand (_02867_, _02505_, _25736_);
  nand (_02868_, _02867_, _29344_);
  nor (_29886_, _02868_, _02866_);
  nor (_02869_, _02505_, _05946_);
  nand (_02870_, _02505_, _25777_);
  nand (_02871_, _02870_, _29344_);
  nor (_29927_, _02871_, _02869_);
  nor (_29968_, _27944_, _23698_);
  not (_02872_, _02683_);
  not (_02873_, _04342_);
  nor (_02874_, _04376_, _02873_);
  nor (_02875_, _02874_, _02872_);
  nor (_30009_, _02875_, _23698_);
  nand (_02876_, _02872_, _29344_);
  nand (_02877_, _30303_, _04342_);
  nand (_30051_, _02877_, _02876_);
  not (_02880_, _04696_);
  nor (_02881_, _02880_, _04340_);
  nor (_30092_, _02881_, _23698_);
  nor (_02882_, _02505_, _04660_);
  nand (_02883_, _02505_, _01701_);
  nand (_02884_, _02883_, _29344_);
  nor (_30132_, _02884_, _02882_);
  nor (_02885_, _02505_, _04658_);
  not (_02886_, _04386_);
  nand (_02887_, _02505_, _02886_);
  nand (_02888_, _02887_, _29344_);
  nor (_30173_, _02888_, _02885_);
  nor (_02889_, _02567_, _04820_);
  nor (_30214_, _02889_, _23698_);
  nand (_02890_, _02585_, _02563_);
  not (_02891_, _02570_);
  nand (_02892_, _30214_, _02891_);
  nor (_30254_, _02892_, _02890_);
  nand (_02893_, _02515_, _04636_);
  nor (_02894_, _02695_, _25682_);
  nand (_02895_, _02894_, _30303_);
  nand (_30352_, _02895_, _02893_);
  nor (_02896_, _25926_, _25746_);
  nor (_02897_, _25805_, _25690_);
  nand (_02898_, _02897_, _02896_);
  not (_02899_, _26110_);
  nor (_02900_, _25710_, _23698_);
  nand (_02901_, _02900_, _02899_);
  nor (_02902_, _02901_, _25990_);
  nor (_02903_, _26049_, _25862_);
  nand (_02904_, _02903_, _02902_);
  nor (_30398_, _02904_, _02898_);
  nor (_30443_, _01721_, _23698_);
  nor (_02905_, _02147_, _25611_);
  nor (_02906_, _02499_, _02495_);
  nor (_02907_, _02906_, _25611_);
  not (_02908_, _02907_);
  nor (_02909_, _02908_, _04417_);
  nor (_02910_, _02907_, _25639_);
  nor (_02911_, _02910_, _02909_);
  nor (_02913_, _02911_, _02905_);
  not (_02914_, _02905_);
  nand (_02915_, _25655_, _04417_);
  nor (_02916_, _02915_, _02914_);
  nand (_02917_, _02916_, _01477_);
  nand (_02918_, _02917_, _25603_);
  nor (_02919_, _02918_, _02913_);
  nor (_30493_, _02919_, _23698_);
  nand (_02920_, _00350_, _29344_);
  nor (_02921_, _01699_, _23698_);
  nand (_02922_, _02921_, _02597_);
  nand (_30539_, _02922_, _02920_);
  nand (_02923_, _02596_, _29344_);
  nor (_02924_, _25682_, _04344_);
  nand (_02925_, _02924_, _25609_);
  nor (_30646_, _25680_, _23698_);
  nand (_02926_, _30646_, _02925_);
  nand (_30600_, _02926_, _02923_);
  nand (_02927_, _04442_, _25680_);
  nor (_30695_, _02927_, _23698_);
  nand (_02928_, _01316_, _04388_);
  nand (_02929_, _02783_, _01583_);
  nand (_02930_, _02929_, _02785_);
  nand (_02931_, _02930_, _01318_);
  nor (_02932_, _01318_, _03080_);
  nor (_02933_, _02932_, _01591_);
  nand (_02934_, _02933_, _02931_);
  nand (_30738_, _02934_, _02928_);
  nand (_02935_, _01316_, _04458_);
  nor (_02936_, _02811_, _04458_);
  nand (_02937_, _02811_, _04458_);
  not (_02938_, _02937_);
  nor (_02939_, _02938_, _02936_);
  nand (_02940_, _02939_, _02815_);
  nor (_02941_, _02939_, _02815_);
  nor (_02942_, _02941_, _01663_);
  nand (_02943_, _02942_, _02940_);
  nor (_02944_, _01318_, _03047_);
  nor (_02945_, _02944_, _01591_);
  nand (_02946_, _02945_, _02943_);
  nand (_30787_, _02946_, _02935_);
  not (_02948_, _04458_);
  nand (_02949_, _02176_, _02948_);
  nand (_02950_, _02175_, _04458_);
  nand (_02951_, _02950_, _02949_);
  nand (_02952_, _02951_, _02109_);
  nand (_02953_, _02952_, _29344_);
  nor (_02954_, _01994_, _03085_);
  nor (_02955_, _01996_, _28411_);
  nor (_02956_, _02955_, _02954_);
  nand (_02957_, _02956_, _02182_);
  nor (_02958_, _02957_, _28271_);
  nand (_02959_, _02957_, _28271_);
  nand (_02960_, _02959_, _02029_);
  nor (_02961_, _02960_, _02958_);
  nand (_02962_, _31253_, _26472_);
  nand (_02963_, _02111_, _31352_);
  nor (_02964_, _02133_, _02948_);
  nor (_02965_, _01691_, _28683_);
  nor (_02966_, _02965_, _02964_);
  nand (_02967_, _02966_, _02963_);
  nor (_02968_, _02967_, _02109_);
  nand (_02969_, _02968_, _02962_);
  nor (_02970_, _02969_, _02961_);
  nor (_30835_, _02970_, _02953_);
  not (_02971_, _30894_);
  nor (_30883_, _02971_, _23698_);
  not (_02972_, _02468_);
  nor (_30925_, _02972_, _23698_);
  nor (_30970_, _28714_, _23698_);
  nor (_31021_, _27590_, _23698_);
  nor (_31068_, _28718_, _23698_);
  nor (_02973_, _02505_, _05924_);
  nand (_02974_, _02505_, _25835_);
  nand (_02975_, _02974_, _29344_);
  nor (_31111_, _02975_, _02973_);
  nor (_02976_, _02505_, _05461_);
  not (_02977_, _04740_);
  nand (_02978_, _02505_, _02977_);
  nand (_02979_, _02978_, _29344_);
  nor (_31155_, _02979_, _02976_);
  nor (_02981_, _26209_, _03332_);
  not (_02982_, _02981_);
  not (_02983_, _01683_);
  nor (_02984_, _02983_, _26274_);
  nor (_02985_, _29169_, _26260_);
  not (_02986_, _02985_);
  nor (_02987_, _02986_, _02984_);
  nand (_02988_, _02987_, _26280_);
  nor (_02989_, _26205_, _01186_);
  nor (_02990_, _02989_, _02988_);
  not (_02991_, _02990_);
  not (_02992_, _26381_);
  nor (_02993_, _26329_, _26069_);
  nor (_02994_, _02993_, _02992_);
  nor (_02995_, _02994_, _26499_);
  nor (_02996_, _26205_, _02992_);
  nor (_02997_, _02011_, _26302_);
  nor (_02998_, _02997_, _02996_);
  nand (_02999_, _02998_, _02995_);
  nand (_03000_, _29193_, _26185_);
  nand (_03001_, _03000_, _26233_);
  not (_03002_, _26318_);
  nand (_03003_, _03002_, _26533_);
  nand (_03004_, _29167_, _26246_);
  nand (_03005_, _03004_, _03003_);
  nor (_03006_, _03005_, _03001_);
  nand (_03007_, _03006_, _26254_);
  nor (_03008_, _03007_, _02999_);
  nor (_03009_, _26286_, _29171_);
  not (_03010_, _03009_);
  nor (_03011_, _29166_, _26286_);
  not (_03012_, _03011_);
  nand (_03013_, _03012_, _03010_);
  nor (_03014_, _03013_, _26136_);
  nor (_03015_, _26195_, _26134_);
  nor (_03016_, _03015_, _02018_);
  nand (_03017_, _03016_, _03014_);
  nor (_03018_, _26292_, _26134_);
  not (_03019_, _03018_);
  nor (_03021_, _03019_, _25706_);
  nor (_03022_, _03021_, _03017_);
  nand (_03023_, _03022_, _03008_);
  nor (_03024_, _03023_, _02991_);
  nor (_03025_, _03024_, _25597_);
  nor (_03026_, _03025_, _02982_);
  nand (_03027_, _26915_, _03332_);
  nand (_03028_, _03027_, _29344_);
  nor (_31199_, _03028_, _03026_);
  nor (_03029_, _25592_, _23698_);
  nand (_03030_, _03029_, _03313_);
  nor (_03031_, _02994_, _29174_);
  not (_03032_, _03031_);
  not (_03033_, _26294_);
  nor (_03034_, _26205_, _03033_);
  not (_03035_, _26136_);
  nand (_03036_, _03035_, _29184_);
  nor (_03037_, _03036_, _03034_);
  nor (_03038_, _26381_, _26294_);
  nor (_03039_, _03038_, _26493_);
  nor (_03040_, _02022_, _26130_);
  nor (_03041_, _03040_, _03039_);
  nand (_03042_, _03041_, _03037_);
  nor (_03043_, _03042_, _03032_);
  nand (_03044_, _26302_, _26266_);
  nand (_03045_, _03044_, _26132_);
  nor (_03046_, _01147_, _01145_);
  nand (_03048_, _03046_, _03045_);
  nand (_03050_, _29172_, _26430_);
  nor (_03051_, _29173_, _26195_);
  not (_03052_, _03051_);
  nand (_03053_, _03052_, _03050_);
  nor (_03054_, _29168_, _26152_);
  nor (_03055_, _03054_, _03053_);
  nor (_03056_, _26205_, _02022_);
  not (_03057_, _03056_);
  nand (_03058_, _03018_, _25708_);
  nand (_03059_, _03058_, _03057_);
  nand (_03060_, _26203_, _26300_);
  nor (_03061_, _26523_, _26237_);
  nand (_03063_, _03061_, _03060_);
  nor (_03064_, _03063_, _03059_);
  nand (_03065_, _03064_, _03055_);
  nor (_03066_, _03065_, _03048_);
  nand (_03067_, _03066_, _03043_);
  nor (_03068_, _25611_, _23698_);
  nand (_03069_, _03068_, _03067_);
  nand (_31248_, _03069_, _03030_);
  nor (_03070_, _26059_, _25597_);
  not (_03071_, _03793_);
  nand (_03072_, _25597_, _03071_);
  nand (_03073_, _03072_, _29344_);
  nor (_31297_, _03073_, _03070_);
  nor (_03075_, _01410_, _25597_);
  not (_03077_, _03796_);
  nand (_03079_, _25597_, _03077_);
  nand (_03081_, _03079_, _29344_);
  nor (_31338_, _03081_, _03075_);
  nor (_03084_, _25872_, _25597_);
  not (_03086_, _03799_);
  nand (_03087_, _25597_, _03086_);
  nand (_03088_, _03087_, _29344_);
  nor (_31379_, _03088_, _03084_);
  nor (_03091_, _26001_, _25597_);
  not (_03092_, _03791_);
  nand (_03093_, _25597_, _03092_);
  nand (_03094_, _03093_, _29344_);
  nor (_00002_, _03094_, _03091_);
  nor (_03095_, _26331_, _25706_);
  not (_03096_, _03095_);
  nor (_03097_, _03096_, _26130_);
  nor (_03098_, _03096_, _26181_);
  nor (_03099_, _03098_, _03097_);
  not (_03100_, _03099_);
  not (_03101_, _26333_);
  not (_03102_, _26130_);
  nor (_03103_, _26179_, _03102_);
  nor (_03104_, _03103_, _03101_);
  nor (_03105_, _03104_, _03100_);
  not (_03106_, _03105_);
  nor (_03108_, _03106_, _03015_);
  nor (_03109_, _03108_, _03100_);
  nand (_00045_, _03109_, _03068_);
  not (_03110_, _03108_);
  nor (_03111_, _03101_, _26130_);
  not (_03112_, _03097_);
  nand (_03114_, _03112_, _03068_);
  nor (_03115_, _03114_, _03111_);
  nand (_00086_, _03115_, _03110_);
  nor (_03117_, _01517_, _01392_);
  nand (_03118_, _01420_, _25870_);
  nor (_03120_, _01438_, _03118_);
  nor (_03121_, _03120_, _03117_);
  nand (_03123_, _01490_, _01486_);
  not (_03124_, _03123_);
  nor (_03125_, _03124_, _03330_);
  nand (_03126_, _03125_, _03121_);
  nor (_03127_, _25607_, _03332_);
  not (_03129_, _03127_);
  nor (_03130_, _03129_, _03783_);
  nand (_03132_, _03130_, _03126_);
  nor (_03133_, _03127_, _26165_);
  nor (_03134_, _03133_, _23698_);
  nand (_00127_, _03134_, _03132_);
  nor (_03136_, _25938_, _25597_);
  not (_03137_, _03785_);
  nand (_03139_, _25597_, _03137_);
  nand (_03140_, _03139_, _29344_);
  nor (_00171_, _03140_, _03136_);
  nor (_03141_, _01400_, _25597_);
  not (_03142_, _03788_);
  nand (_03143_, _25597_, _03142_);
  nand (_03144_, _03143_, _29344_);
  nor (_00215_, _03144_, _03141_);
  nor (_00262_, _26478_, _23698_);
  not (_03145_, _26549_);
  nor (_00304_, _03145_, _23698_);
  nor (_03146_, _25817_, _25597_);
  not (_03147_, _03802_);
  nand (_03148_, _25597_, _03147_);
  nand (_03150_, _03148_, _29344_);
  nor (_00353_, _03150_, _03146_);
  nor (_03151_, _03096_, _26205_);
  not (_03152_, _03151_);
  nand (_03153_, _03152_, _03057_);
  not (_03154_, _26406_);
  nor (_03155_, _03154_, _26333_);
  nor (_03156_, _03155_, _26205_);
  nor (_03157_, _03156_, _03153_);
  not (_03158_, _26539_);
  nor (_03159_, _26205_, _26248_);
  not (_03160_, _26284_);
  nor (_03161_, _03160_, _26134_);
  nor (_03162_, _03161_, _03159_);
  nor (_03163_, _29168_, _29164_);
  nor (_03164_, _26205_, _02009_);
  nor (_03165_, _03164_, _03163_);
  nand (_03166_, _03165_, _03162_);
  nor (_03168_, _03166_, _03158_);
  nand (_03170_, _03168_, _03157_);
  nand (_03171_, _26154_, _26179_);
  nand (_03173_, _03171_, _03035_);
  nor (_03175_, _03054_, _03009_);
  nand (_03176_, _03175_, _26525_);
  nor (_03178_, _03176_, _03173_);
  nor (_03179_, _29169_, _26513_);
  nor (_03180_, _03051_, _03034_);
  nand (_03182_, _03180_, _03179_);
  not (_03184_, _26142_);
  nor (_03186_, _29192_, _03184_);
  nand (_03187_, _29167_, _26430_);
  nand (_03189_, _03187_, _29175_);
  nor (_03190_, _03189_, _03186_);
  not (_03191_, _26335_);
  nor (_03192_, _29188_, _03191_);
  nand (_03193_, _03192_, _03190_);
  nor (_03195_, _03193_, _03182_);
  nand (_03196_, _03195_, _03178_);
  nor (_03197_, _03196_, _03170_);
  nor (_03198_, _03197_, _25611_);
  nand (_03200_, _03815_, _03332_);
  nor (_03201_, _26466_, _03330_);
  nand (_03202_, _03109_, _03201_);
  nand (_03203_, _03202_, _03200_);
  nor (_03204_, _03203_, _03198_);
  nor (_00395_, _03204_, _23698_);
  nand (_03205_, _03029_, _03089_);
  nor (_03206_, _26177_, _26069_);
  nand (_03207_, _03206_, _26154_);
  nor (_03208_, _02983_, _26266_);
  nor (_03209_, _26205_, _26266_);
  nor (_03210_, _03209_, _03208_);
  nand (_03211_, _03210_, _03207_);
  nor (_03212_, _26205_, _03101_);
  not (_03213_, _03212_);
  nand (_03214_, _03015_, _25706_);
  nand (_03215_, _03214_, _03213_);
  not (_03216_, _03215_);
  not (_03217_, _26144_);
  nor (_03218_, _26185_, _03217_);
  nor (_03219_, _03218_, _29192_);
  not (_03220_, _03163_);
  nand (_03221_, _03220_, _03003_);
  nor (_03222_, _03221_, _03219_);
  nand (_03223_, _03222_, _03216_);
  nor (_03224_, _03223_, _03211_);
  not (_03225_, _03159_);
  not (_03226_, _26205_);
  nand (_03227_, _26442_, _26511_);
  nand (_03228_, _03227_, _03226_);
  nand (_03229_, _03228_, _03225_);
  not (_03230_, _26349_);
  nor (_03231_, _26499_, _03230_);
  not (_03232_, _26250_);
  not (_03233_, _26521_);
  nand (_03234_, _03233_, _03232_);
  nor (_03235_, _03234_, _26395_);
  nand (_03236_, _03235_, _03231_);
  nor (_03237_, _03236_, _03229_);
  nand (_03238_, _03237_, _03224_);
  nand (_03240_, _03238_, _03068_);
  nand (_00441_, _03240_, _03205_);
  nor (_03241_, _26171_, _26296_);
  nand (_03242_, _26213_, _03201_);
  not (_03243_, _03242_);
  nor (_03244_, _02006_, _25706_);
  not (_03245_, _03244_);
  nor (_03246_, _03245_, _26171_);
  nor (_03247_, _03246_, _03243_);
  not (_03248_, _03247_);
  nor (_03249_, _03248_, _03241_);
  not (_03250_, _03249_);
  nand (_03251_, _03821_, _03332_);
  nand (_03252_, _26446_, _26391_);
  nand (_03253_, _26420_, _26231_);
  nand (_03254_, _03253_, _26371_);
  nor (_03255_, _03254_, _03252_);
  nand (_03256_, _03255_, _26254_);
  nor (_03257_, _26199_, _29171_);
  nor (_03258_, _03096_, _26327_);
  nor (_03259_, _03258_, _03257_);
  not (_03260_, _26436_);
  nor (_03261_, _26509_, _03260_);
  nand (_03262_, _03261_, _03259_);
  not (_03263_, _03262_);
  nand (_03264_, _03263_, _03245_);
  nor (_03265_, _03264_, _03256_);
  nor (_03266_, _26414_, _26144_);
  nor (_03267_, _03266_, _01182_);
  nand (_03269_, _03267_, _26280_);
  nor (_03271_, _03269_, _26353_);
  not (_03273_, _03271_);
  nor (_03275_, _03273_, _26428_);
  nand (_03277_, _03275_, _03265_);
  nand (_03279_, _03277_, _25609_);
  nand (_03281_, _03279_, _03251_);
  nor (_03283_, _03281_, _03250_);
  nor (_00485_, _03283_, _23698_);
  nor (_03286_, _03096_, _26493_);
  nor (_03288_, _03286_, _26320_);
  nand (_03292_, _03288_, _03245_);
  nor (_03294_, _26493_, _02009_);
  nor (_03296_, _03294_, _26499_);
  not (_03298_, _26446_);
  nor (_03300_, _26503_, _03298_);
  nand (_03302_, _03300_, _03296_);
  nor (_03303_, _03302_, _03292_);
  nor (_03304_, _03303_, _25611_);
  nand (_03305_, _03823_, _03332_);
  nand (_03306_, _03305_, _03247_);
  nor (_03307_, _03306_, _03304_);
  nor (_00530_, _03307_, _23698_);
  nand (_03309_, _03813_, _03332_);
  nand (_03310_, _26207_, _25592_);
  nand (_03311_, _03310_, _03309_);
  nand (_03312_, _03311_, _29344_);
  nor (_03314_, _02993_, _25708_);
  nor (_03315_, _03314_, _03226_);
  nor (_03316_, _03315_, _26292_);
  not (_03317_, _29174_);
  nor (_03318_, _26503_, _26424_);
  nand (_03319_, _03318_, _03317_);
  nor (_03320_, _03319_, _03316_);
  not (_03321_, _03320_);
  not (_03322_, _02995_);
  nor (_03323_, _03018_, _26268_);
  not (_03324_, _03323_);
  nor (_03325_, _03324_, _03322_);
  nor (_03326_, _26266_, _26130_);
  nor (_03327_, _03326_, _03151_);
  nand (_03328_, _03327_, _03325_);
  nor (_03329_, _03328_, _03321_);
  nand (_03331_, _03329_, _02990_);
  nand (_03333_, _03331_, _03068_);
  nand (_00579_, _03333_, _03312_);
  nand (_03334_, _03029_, _30689_);
  nor (_03335_, _26300_, _01682_);
  nor (_03336_, _03335_, _26134_);
  not (_03337_, _26357_);
  nand (_03338_, _03337_, _26239_);
  nor (_03340_, _03338_, _03336_);
  nor (_03342_, _02983_, _26152_);
  nor (_03343_, _03342_, _03011_);
  nand (_03344_, _03343_, _03175_);
  nor (_03345_, _03021_, _03056_);
  nand (_03346_, _26420_, _26132_);
  nand (_03347_, _03346_, _01735_);
  nor (_03348_, _03347_, _01145_);
  nand (_03349_, _03348_, _03345_);
  nor (_03350_, _03349_, _03344_);
  nand (_03351_, _03350_, _03340_);
  nand (_03352_, _03351_, _03068_);
  nand (_00620_, _03352_, _03334_);
  nor (_03353_, _03811_, _25592_);
  nor (_03354_, _03353_, _02981_);
  nor (_03356_, _03212_, _03054_);
  nor (_03357_, _03342_, _01736_);
  nand (_03359_, _03357_, _03356_);
  nand (_03361_, _26288_, _26132_);
  nand (_03363_, _03361_, _01141_);
  nor (_03365_, _03363_, _03359_);
  nand (_03367_, _03365_, _03327_);
  nor (_03368_, _02999_, _02988_);
  nand (_03369_, _03368_, _03320_);
  nor (_03370_, _03369_, _03367_);
  nor (_03371_, _03370_, _25611_);
  nor (_03372_, _03371_, _03354_);
  nor (_00663_, _03372_, _23698_);
  nand (_03373_, _03154_, _26069_);
  not (_03374_, _26341_);
  not (_03375_, _26371_);
  nor (_03376_, _03375_, _03374_);
  nand (_03377_, _03376_, _03373_);
  nor (_03378_, _03377_, _03032_);
  nand (_03379_, _03378_, _03263_);
  nand (_03380_, _26426_, _26383_);
  nor (_03381_, _29173_, _03184_);
  nor (_03382_, _03381_, _26503_);
  nand (_03383_, _03382_, _26410_);
  nor (_03384_, _03383_, _26450_);
  not (_03386_, _03296_);
  nor (_03387_, _03386_, _26256_);
  nand (_03388_, _03387_, _03384_);
  nor (_03389_, _03388_, _03380_);
  nor (_03390_, _03292_, _03273_);
  nand (_03391_, _03390_, _03389_);
  nor (_03392_, _03391_, _03379_);
  nor (_03393_, _03392_, _25611_);
  nand (_03394_, _03366_, _03332_);
  nand (_03395_, _03394_, _03249_);
  nor (_03396_, _03395_, _03393_);
  nor (_00704_, _03396_, _23698_);
  nand (_03397_, _03344_, _03068_);
  nand (_03398_, _26213_, _25592_);
  nand (_03399_, _03332_, _30685_);
  nand (_03400_, _03399_, _03398_);
  nand (_03401_, _03400_, _29344_);
  nand (_00745_, _03401_, _03397_);
  nand (_03402_, _03029_, _03358_);
  nand (_03403_, _29191_, _03217_);
  nand (_03404_, _03403_, _03233_);
  nor (_03405_, _03404_, _03163_);
  nand (_03406_, _03323_, _29200_);
  nor (_03407_, _03406_, _03363_);
  nand (_03408_, _03407_, _03405_);
  nor (_03409_, _03408_, _03321_);
  nand (_03410_, _03409_, _03008_);
  nand (_03411_, _03410_, _03068_);
  nand (_00787_, _03411_, _03402_);
  nand (_03412_, _03029_, _03308_);
  nand (_03413_, _03043_, _26355_);
  nand (_03414_, _03413_, _03068_);
  nand (_00830_, _03414_, _03412_);
  not (_03415_, _03202_);
  nand (_03416_, _03245_, _03214_);
  nand (_03417_, _03416_, _25599_);
  nor (_03418_, _03246_, _03332_);
  nand (_03419_, _03418_, _03417_);
  nor (_03420_, _03419_, _03415_);
  nand (_03421_, _03332_, _26949_);
  nand (_03423_, _03421_, _29344_);
  nor (_00872_, _03423_, _03420_);
  nand (_03424_, _03375_, _25595_);
  nand (_03425_, _03424_, _25592_);
  nor (_03426_, _03425_, _03243_);
  nand (_03427_, _26578_, _03332_);
  nand (_03428_, _03427_, _29344_);
  nor (_00910_, _03428_, _03426_);
  nand (_03429_, _03029_, _03090_);
  nor (_03430_, _03211_, _26136_);
  nand (_03431_, _03430_, _03320_);
  nand (_03432_, _03431_, _03068_);
  nand (_00945_, _03432_, _03429_);
  not (_03433_, _02994_);
  nor (_03434_, _02996_, _26499_);
  nand (_03435_, _03434_, _03433_);
  nor (_03436_, _03173_, _03435_);
  nor (_03437_, _03436_, _25611_);
  nand (_03438_, _03360_, _03332_);
  nand (_03439_, _03438_, _03242_);
  nor (_03440_, _03439_, _03437_);
  nor (_00987_, _03440_, _23698_);
  nand (_03441_, _03029_, _03049_);
  nor (_03442_, _03346_, _25708_);
  not (_03443_, _03040_);
  nand (_03444_, _03443_, _26306_);
  nor (_03445_, _03444_, _03442_);
  nor (_03446_, _02021_, _29181_);
  nor (_03447_, _02019_, _01737_);
  nand (_03448_, _03447_, _03446_);
  nor (_03449_, _03448_, _03215_);
  nand (_03450_, _03449_, _03445_);
  nand (_03451_, _03450_, _03068_);
  nand (_01038_, _03451_, _03441_);
  nor (_03452_, _25759_, _25597_);
  not (_03453_, _03341_);
  nand (_03454_, _25597_, _03453_);
  nand (_03455_, _03454_, _29344_);
  nor (_01071_, _03455_, _03452_);
  not (_03456_, _01497_);
  nor (_03458_, _03456_, _25872_);
  not (_03459_, _01514_);
  nand (_03460_, _03459_, _01463_);
  nor (_03461_, _03460_, _03458_);
  not (_03462_, _01431_);
  not (_03463_, _01503_);
  nor (_03464_, _03463_, _01390_);
  nor (_03465_, _03464_, _01428_);
  nand (_03466_, _03465_, _03462_);
  nand (_03467_, _01467_, _01437_);
  not (_03468_, _01466_);
  nand (_03469_, _01528_, _03468_);
  nand (_03470_, _03469_, _01403_);
  nand (_03471_, _03470_, _03467_);
  nor (_03472_, _03471_, _03466_);
  nand (_03473_, _03472_, _01418_);
  nor (_03474_, _03473_, _03126_);
  nand (_03475_, _03474_, _03461_);
  nand (_03476_, _03475_, _25613_);
  nor (_03477_, _03130_, _26167_);
  nor (_03478_, _03477_, _23698_);
  nand (_01105_, _03478_, _03476_);
  not (_03479_, _03068_);
  nor (_03480_, _03479_, _03015_);
  nand (_01142_, _03480_, _03106_);
  nor (_01181_, _26219_, _23698_);
  nor (_03481_, _03151_, _03056_);
  nand (_03482_, _26406_, _03101_);
  nand (_03483_, _03482_, _03226_);
  nand (_03484_, _03483_, _03481_);
  nand (_03485_, _26284_, _26132_);
  not (_03486_, _26331_);
  nand (_03487_, _26385_, _03486_);
  nand (_03488_, _03487_, _03485_);
  nand (_03489_, _03095_, _26316_);
  nand (_03490_, _03011_, _26128_);
  nand (_03491_, _03490_, _03489_);
  nor (_03492_, _03491_, _03488_);
  nand (_03493_, _03492_, _03055_);
  nor (_03494_, _03493_, _03484_);
  nand (_03496_, _26302_, _26274_);
  nand (_03497_, _03496_, _26329_);
  nor (_03498_, _26213_, _26158_);
  nand (_03499_, _03498_, _03497_);
  not (_03500_, _01686_);
  not (_03501_, _02996_);
  nand (_03502_, _03501_, _03500_);
  not (_03503_, _02984_);
  not (_03504_, _03034_);
  nand (_03505_, _03504_, _03503_);
  nor (_03506_, _03505_, _03502_);
  not (_03507_, _26276_);
  nor (_03508_, _29192_, _26286_);
  nor (_03509_, _29173_, _26331_);
  nor (_03510_, _03509_, _03508_);
  nand (_03511_, _03510_, _03507_);
  not (_03512_, _26523_);
  nand (_03513_, _03512_, _26363_);
  nor (_03514_, _03513_, _03511_);
  nand (_03515_, _03514_, _03506_);
  nor (_03516_, _03515_, _03499_);
  nand (_03517_, _03516_, _03494_);
  not (_03518_, _26351_);
  nor (_03519_, _03518_, _26278_);
  not (_03520_, _26252_);
  nand (_03521_, _03171_, _03520_);
  nor (_03522_, _03521_, _03266_);
  nand (_03523_, _03522_, _03519_);
  nor (_03524_, _03523_, _03517_);
  nor (_03525_, _03524_, _25611_);
  nand (_03526_, _03332_, _03181_);
  nor (_03527_, _03398_, _25599_);
  nor (_03528_, _03527_, _03415_);
  nand (_03529_, _03528_, _03526_);
  nor (_03530_, _03529_, _03525_);
  nor (_01232_, _03530_, _23698_);
  not (_03531_, _03416_);
  not (_03532_, _03294_);
  nand (_03533_, _29173_, _26205_);
  nand (_03534_, _03533_, _03217_);
  nand (_03536_, _03534_, _03532_);
  nor (_03537_, _03536_, _03229_);
  nand (_03538_, _03537_, _03531_);
  nor (_03539_, _03538_, _03517_);
  nor (_03540_, _03539_, _25611_);
  nand (_03541_, _03332_, _03174_);
  nand (_03542_, _03541_, _03528_);
  nor (_03543_, _03542_, _03540_);
  nor (_01282_, _03543_, _23698_);
  nor (_01328_, _01764_, _23698_);
  nor (_01371_, _01795_, _23698_);
  nor (_01419_, _01826_, _23698_);
  nor (_01471_, _01855_, _23698_);
  nor (_01518_, _01884_, _23698_);
  nor (_01559_, _01914_, _23698_);
  nor (_01602_, _01941_, _23698_);
  nor (_01643_, _28838_, _23698_);
  nor (_01680_, _28891_, _23698_);
  nor (_01727_, _28736_, _23698_);
  nor (_01770_, _28966_, _23698_);
  nor (_01811_, _29027_, _23698_);
  nor (_01852_, _28060_, _23698_);
  nor (_01895_, _27940_, _23698_);
  nor (_01937_, _25815_, _23698_);
  nor (_01979_, _25870_, _23698_);
  nor (_02032_, _25698_, _23698_);
  nor (_02073_, _26057_, _23698_);
  nor (_02117_, _25998_, _23698_);
  nor (_02160_, _26118_, _23698_);
  nor (_02200_, _25936_, _23698_);
  nor (_02246_, _28683_, _23698_);
  nor (_02286_, _25757_, _23698_);
  nor (_02326_, _31337_, _23698_);
  nor (_02366_, _29651_, _23698_);
  not (_03544_, _30213_);
  nor (_02404_, _03544_, _23698_);
  nor (_02443_, _30357_, _23698_);
  nor (_02481_, _00159_, _23698_);
  not (_03545_, _30649_);
  nor (_02509_, _03545_, _23698_);
  not (_03547_, _30778_);
  nor (_02542_, _03547_, _23698_);
  nor (_02575_, _30840_, _23698_);
  nor (_02611_, _31052_, _23698_);
  nor (_02644_, _00138_, _23698_);
  nor (_02677_, _00079_, _23698_);
  nor (_02711_, _29502_, _23698_);
  nor (_02743_, _29649_, _23698_);
  nor (_03548_, _29346_, _29351_);
  nand (_03549_, _29346_, _29351_);
  nand (_03550_, _03549_, _29344_);
  nor (_02774_, _03550_, _03548_);
  nor (_03551_, _03548_, _29349_);
  not (_03552_, _03548_);
  nor (_03553_, _03552_, _02093_);
  nor (_03554_, _03553_, _03551_);
  nor (_02814_, _03554_, _23698_);
  nor (_02846_, _31107_, _23698_);
  nor (_02879_, _30199_, _23698_);
  not (_03555_, _30362_);
  nor (_02912_, _03555_, _23698_);
  not (_03556_, _30485_);
  nor (_02947_, _03556_, _23698_);
  nor (_02980_, _30653_, _23698_);
  nor (_03020_, _30788_, _23698_);
  nor (_03062_, _30844_, _23698_);
  nor (_03107_, _31284_, _23698_);
  nor (_03149_, _31157_, _23698_);
  nor (_03199_, _31104_, _23698_);
  nor (_03239_, _31043_, _23698_);
  nor (_03290_, _00132_, _23698_);
  nor (_03339_, _00062_, _23698_);
  nor (_03385_, _31385_, _23698_);
  nor (_03422_, _29786_, _23698_);
  nor (_03557_, _29653_, _29661_);
  nor (_03558_, _30195_, _01904_);
  nor (_03559_, _03558_, _03557_);
  nor (_03457_, _03559_, _23698_);
  nor (_03560_, _29653_, _29664_);
  nor (_03561_, _30195_, _29668_);
  nor (_03563_, _03561_, _03560_);
  nor (_03495_, _03563_, _23698_);
  nor (_03535_, _31332_, _23698_);
  nor (_03546_, _31126_, _23698_);
  nor (_03562_, _31062_, _23698_);
  nor (_03592_, _00167_, _23698_);
  nor (_03631_, _00102_, _23698_);
  nor (_03669_, _31415_, _23698_);
  nor (_03708_, _00044_, _23698_);
  nor (_03744_, _31322_, _23698_);
  nand (_03564_, _00783_, _30948_);
  nor (_03565_, _03564_, _26895_);
  not (_03566_, _03565_);
  nor (_03567_, _03566_, _31419_);
  nor (_03568_, _03565_, _01589_);
  not (_03569_, _03568_);
  nand (_03570_, _03569_, _26787_);
  nor (_03571_, _03570_, _03567_);
  nand (_03572_, _29294_, _01589_);
  nand (_03573_, _03565_, _30943_);
  nor (_03574_, _03568_, _29297_);
  nand (_03575_, _03574_, _03573_);
  nand (_03576_, _03575_, _03572_);
  nor (_03577_, _03576_, _03571_);
  nor (_03782_, _03577_, _23698_);
  nor (_03578_, _03566_, _30828_);
  not (_03579_, _01597_);
  nand (_03580_, _03566_, _03579_);
  nand (_03581_, _03580_, _26787_);
  nor (_03582_, _03581_, _03578_);
  nand (_03583_, _29294_, _01597_);
  nor (_03584_, _03564_, _31399_);
  nand (_03585_, _03584_, _30943_);
  nor (_03586_, _03584_, _01597_);
  nor (_03587_, _03586_, _29297_);
  nand (_03588_, _03587_, _03585_);
  nand (_03589_, _03588_, _03583_);
  nor (_03590_, _03589_, _03582_);
  nor (_03836_, _03590_, _23698_);
  nor (_03591_, _03566_, _30692_);
  nand (_03593_, _03566_, _30569_);
  nand (_03594_, _03593_, _26787_);
  nor (_03595_, _03594_, _03591_);
  nand (_03596_, _29294_, _01606_);
  nor (_03597_, _03564_, _00092_);
  nand (_03598_, _03597_, _30943_);
  nor (_03599_, _03597_, _01606_);
  nor (_03600_, _03599_, _29297_);
  nand (_03601_, _03600_, _03598_);
  nand (_03602_, _03601_, _03596_);
  nor (_03603_, _03602_, _03595_);
  nor (_03873_, _03603_, _23698_);
  nor (_03604_, _03566_, _00164_);
  nand (_03605_, _03566_, _00678_);
  nand (_03606_, _03605_, _26787_);
  nor (_03607_, _03606_, _03604_);
  nand (_03608_, _29294_, _01620_);
  nor (_03609_, _03564_, _00105_);
  nand (_03610_, _03609_, _30943_);
  nor (_03611_, _03609_, _01620_);
  nor (_03612_, _03611_, _29297_);
  nand (_03613_, _03612_, _03610_);
  nand (_03614_, _03613_, _03608_);
  nor (_03615_, _03614_, _03607_);
  nor (_03910_, _03615_, _23698_);
  nor (_03616_, _03566_, _02217_);
  nand (_03617_, _03566_, _30272_);
  nand (_03618_, _03617_, _26787_);
  nor (_03619_, _03618_, _03616_);
  nand (_03620_, _29294_, _01627_);
  nor (_03621_, _03564_, _30954_);
  nand (_03622_, _03621_, _30943_);
  nor (_03623_, _03621_, _01627_);
  nor (_03624_, _03623_, _29297_);
  nand (_03625_, _03624_, _03622_);
  nand (_03626_, _03625_, _03620_);
  nor (_03627_, _03626_, _03619_);
  nor (_03951_, _03627_, _23698_);
  nor (_03628_, _03566_, _31067_);
  not (_03629_, _01585_);
  nand (_03632_, _03566_, _03629_);
  nand (_03633_, _03632_, _26787_);
  nor (_03634_, _03633_, _03628_);
  nand (_03635_, _29294_, _01585_);
  nor (_03636_, _03564_, _31071_);
  nand (_03637_, _03636_, _30943_);
  nor (_03638_, _03636_, _01585_);
  nor (_03639_, _03638_, _29297_);
  nand (_03640_, _03639_, _03637_);
  nand (_03641_, _03640_, _03635_);
  nor (_03642_, _03641_, _03634_);
  nor (_03990_, _03642_, _23698_);
  nor (_03643_, _03566_, _31328_);
  nand (_03644_, _03566_, _00687_);
  nand (_03645_, _03644_, _26787_);
  nor (_03646_, _03645_, _03643_);
  nand (_03647_, _29294_, _01609_);
  nor (_03648_, _03564_, _31182_);
  nand (_03649_, _03648_, _30943_);
  nor (_03650_, _03648_, _01609_);
  nor (_03651_, _03650_, _29297_);
  nand (_03652_, _03651_, _03649_);
  nand (_03653_, _03652_, _03647_);
  nor (_03654_, _03653_, _03646_);
  nor (_04030_, _03654_, _23698_);
  nor (_03655_, _03566_, _31253_);
  nand (_03656_, _03566_, _00676_);
  nand (_03657_, _03656_, _26787_);
  nor (_03658_, _03657_, _03655_);
  nand (_03659_, _29294_, _01617_);
  nor (_03660_, _03564_, _31259_);
  nand (_03661_, _03660_, _30943_);
  nor (_03662_, _03660_, _01617_);
  nor (_03663_, _03662_, _29297_);
  nand (_03664_, _03663_, _03661_);
  nand (_03665_, _03664_, _03659_);
  nor (_03666_, _03665_, _03658_);
  nor (_04068_, _03666_, _23698_);
  nor (_03667_, _30882_, _00792_);
  not (_03668_, _03667_);
  nor (_03670_, _26789_, _27726_);
  not (_03671_, _03670_);
  nor (_03672_, _03671_, _00105_);
  not (_03673_, _03672_);
  nor (_03674_, _03673_, _03668_);
  not (_03675_, _03674_);
  nor (_03676_, _03675_, _00828_);
  not (_03677_, _01488_);
  nand (_03678_, _01226_, _01224_);
  nor (_03679_, _00888_, _00841_);
  not (_03680_, _03679_);
  nor (_03681_, _03680_, _00243_);
  not (_03682_, _03681_);
  nor (_03683_, _03682_, _03678_);
  not (_03684_, _03683_);
  nor (_03685_, _03671_, _00092_);
  not (_03686_, _03685_);
  nor (_03687_, _03686_, _03668_);
  nor (_03688_, _03687_, _03684_);
  nor (_03689_, _03688_, _03677_);
  not (_03690_, _01265_);
  not (_03691_, _03688_);
  nor (_03692_, _03691_, _03690_);
  nor (_03693_, _03692_, _03689_);
  nand (_03694_, _03693_, _03675_);
  nand (_03695_, _03694_, _29344_);
  nor (_04107_, _03695_, _03676_);
  nor (_03696_, _03675_, _00750_);
  not (_03697_, _01485_);
  nor (_03698_, _03688_, _03697_);
  not (_03699_, _01432_);
  nor (_03700_, _03691_, _03699_);
  nor (_03701_, _03700_, _03698_);
  nand (_03702_, _03701_, _03675_);
  nand (_03703_, _03702_, _29344_);
  nor (_04145_, _03703_, _03696_);
  nor (_03704_, _03675_, _00800_);
  not (_03705_, _01482_);
  nor (_03706_, _03688_, _03705_);
  nor (_03707_, _03691_, _30300_);
  nor (_03709_, _03707_, _03706_);
  nand (_03710_, _03709_, _03675_);
  nand (_03711_, _03710_, _29344_);
  nor (_04184_, _03711_, _03704_);
  nor (_03712_, _03675_, _27742_);
  not (_03713_, _01479_);
  nor (_03714_, _03688_, _03713_);
  not (_03715_, _01405_);
  nor (_03716_, _03691_, _03715_);
  nor (_03717_, _03716_, _03714_);
  nand (_03718_, _03717_, _03675_);
  nand (_03719_, _03718_, _29344_);
  nor (_04222_, _03719_, _03712_);
  nor (_03720_, _03675_, _00811_);
  not (_03721_, _01476_);
  nor (_03722_, _03688_, _03721_);
  nor (_03723_, _03691_, _30584_);
  nor (_03724_, _03723_, _03722_);
  nand (_03725_, _03724_, _03675_);
  nand (_03726_, _03725_, _29344_);
  nor (_04255_, _03726_, _03720_);
  nor (_03727_, _03675_, _28244_);
  not (_03728_, _01473_);
  nor (_03729_, _03688_, _03728_);
  not (_03730_, _01412_);
  nor (_03731_, _03691_, _03730_);
  nor (_03732_, _03731_, _03729_);
  nand (_03733_, _03732_, _03675_);
  nand (_03734_, _03733_, _29344_);
  nor (_04294_, _03734_, _03727_);
  nor (_03735_, _03688_, _01469_);
  nor (_03736_, _03691_, _01295_);
  nor (_03737_, _03736_, _03735_);
  nor (_03738_, _03737_, _03674_);
  nand (_03739_, _03674_, _27888_);
  nand (_03740_, _03739_, _29344_);
  nor (_04331_, _03740_, _03738_);
  not (_03741_, _01459_);
  nor (_03742_, _03683_, _03741_);
  not (_03743_, _01369_);
  nor (_03745_, _03684_, _03743_);
  nor (_03746_, _03745_, _03742_);
  nor (_03747_, _03746_, _03687_);
  not (_03748_, _03687_);
  nor (_03749_, _03748_, _28639_);
  nor (_03750_, _03749_, _03747_);
  nor (_03751_, _03750_, _03674_);
  nor (_03752_, _03675_, _03741_);
  nor (_03753_, _03752_, _03751_);
  nor (_04374_, _03753_, _23698_);
  not (_03754_, _01456_);
  nor (_03755_, _03683_, _03754_);
  not (_03756_, _01389_);
  nor (_03757_, _03684_, _03756_);
  nor (_03758_, _03757_, _03755_);
  nor (_03759_, _03758_, _03687_);
  nor (_03760_, _03748_, _28598_);
  nor (_03761_, _03760_, _03759_);
  nor (_03762_, _03761_, _03674_);
  nor (_03763_, _03675_, _03754_);
  nor (_03764_, _03763_, _03762_);
  nor (_04420_, _03764_, _23698_);
  nor (_03765_, _00105_, _27726_);
  nand (_03766_, _03765_, _03667_);
  nor (_03767_, _03766_, _26789_);
  nand (_03768_, _03687_, _27584_);
  nor (_03769_, _03683_, _30298_);
  nor (_03770_, _03684_, _30311_);
  nor (_03771_, _03770_, _03769_);
  nand (_03772_, _03771_, _03748_);
  nand (_03773_, _03772_, _03768_);
  nor (_03774_, _03773_, _03767_);
  nor (_03775_, _03675_, _30298_);
  nor (_03776_, _03775_, _03774_);
  nor (_04460_, _03776_, _23698_);
  nor (_03777_, _03748_, _27742_);
  not (_03778_, _01450_);
  nor (_03779_, _03683_, _03778_);
  not (_03780_, _01415_);
  nor (_03781_, _03684_, _03780_);
  nor (_03784_, _03781_, _03779_);
  nand (_03786_, _03784_, _03748_);
  nand (_03787_, _03786_, _03675_);
  nor (_03789_, _03787_, _03777_);
  nor (_03790_, _03675_, _03778_);
  nor (_03792_, _03790_, _03789_);
  nor (_04499_, _03792_, _23698_);
  nor (_03794_, _27726_, _26640_);
  not (_03795_, _03794_);
  nor (_03797_, _03795_, _02097_);
  nand (_03798_, _03797_, _29298_);
  not (_03800_, _03798_);
  not (_03801_, _01259_);
  not (_03803_, _03678_);
  nand (_03804_, _03803_, _03801_);
  nand (_03805_, _03804_, _00421_);
  nor (_03806_, _03805_, _03800_);
  nor (_03807_, _31182_, _30943_);
  nand (_03808_, _31182_, _01249_);
  nand (_03810_, _03808_, _03800_);
  nor (_03812_, _03810_, _03807_);
  nor (_03814_, _03812_, _03806_);
  nor (_03816_, _03671_, _26895_);
  not (_03818_, _03816_);
  nor (_03820_, _03818_, _03668_);
  nor (_03822_, _03820_, _03814_);
  nand (_03824_, _03820_, _28639_);
  nand (_03825_, _03824_, _29344_);
  nor (_04538_, _03825_, _03822_);
  nor (_03826_, _03798_, _31071_);
  not (_03827_, _03826_);
  nor (_03828_, _03827_, _30944_);
  nor (_03829_, _03826_, _00841_);
  nor (_03830_, _03829_, _03828_);
  nor (_03831_, _03830_, _03820_);
  nand (_03832_, _03820_, _28598_);
  nand (_03833_, _03832_, _29344_);
  nor (_04575_, _03833_, _03831_);
  nand (_03834_, _03800_, _30953_);
  nor (_03835_, _03834_, _30944_);
  not (_03837_, _03820_);
  nand (_03838_, _03834_, _30307_);
  nand (_03839_, _03838_, _03837_);
  nor (_03840_, _03839_, _03835_);
  nor (_03841_, _03837_, _27584_);
  nor (_03842_, _03841_, _03840_);
  nor (_04610_, _03842_, _23698_);
  nand (_03843_, _03800_, _00104_);
  nor (_03844_, _03843_, _30944_);
  nand (_03845_, _03843_, _00442_);
  nand (_03846_, _03845_, _03837_);
  nor (_03847_, _03846_, _03844_);
  nor (_03848_, _03837_, _27718_);
  nor (_03849_, _03848_, _03847_);
  nor (_04651_, _03849_, _23698_);
  nor (_03850_, _03798_, _00092_);
  not (_03851_, _03850_);
  nor (_03852_, _03851_, _30944_);
  nor (_03853_, _03850_, _01238_);
  nor (_03854_, _03853_, _03852_);
  nor (_03855_, _03854_, _03820_);
  nand (_03856_, _03820_, _28540_);
  nand (_03857_, _03856_, _29344_);
  nor (_04691_, _03857_, _03855_);
  nor (_03858_, _03798_, _31399_);
  not (_03859_, _03858_);
  nor (_03860_, _03859_, _30944_);
  nor (_03861_, _03858_, _01229_);
  nor (_03862_, _03861_, _03860_);
  nor (_03863_, _03862_, _03820_);
  nand (_03864_, _03820_, _28157_);
  nand (_03865_, _03864_, _29344_);
  nor (_04735_, _03865_, _03863_);
  nand (_03866_, _03687_, _28540_);
  nor (_03867_, _03683_, _30581_);
  nor (_03868_, _03684_, _30595_);
  nor (_03869_, _03868_, _03867_);
  nand (_03870_, _03869_, _03748_);
  nand (_03871_, _03870_, _03866_);
  nor (_03872_, _03871_, _03767_);
  nor (_03874_, _03675_, _30581_);
  nor (_03875_, _03874_, _03872_);
  nor (_04784_, _03875_, _23698_);
  nand (_03876_, _03800_, _26893_);
  nor (_03877_, _03876_, _30944_);
  nand (_03878_, _03876_, _00243_);
  nand (_03879_, _03878_, _03837_);
  nor (_03880_, _03879_, _03877_);
  nor (_03881_, _03837_, _27888_);
  nor (_03882_, _03881_, _03880_);
  nor (_04831_, _03882_, _23698_);
  nor (_03883_, _03748_, _28244_);
  nand (_03884_, _03684_, _01444_);
  nand (_03885_, _03683_, _01421_);
  nand (_03886_, _03885_, _03884_);
  nor (_03887_, _03886_, _03687_);
  nor (_03888_, _03887_, _03883_);
  nor (_03889_, _03888_, _03674_);
  not (_03890_, _01444_);
  nand (_03891_, _03674_, _03890_);
  nand (_03892_, _03891_, _29344_);
  nor (_04874_, _03892_, _03889_);
  nor (_03893_, _03683_, _01441_);
  nor (_03894_, _03684_, _01423_);
  nor (_03895_, _03894_, _03893_);
  nor (_03896_, _03895_, _03687_);
  nor (_03897_, _03748_, _27886_);
  nor (_03898_, _03897_, _03896_);
  nor (_03899_, _03898_, _03674_);
  nand (_03900_, _03674_, _00235_);
  nand (_03901_, _03900_, _29344_);
  nor (_04922_, _03901_, _03899_);
  nor (_03902_, _03678_, _01252_);
  nand (_03903_, _03902_, _03679_);
  not (_03904_, _03903_);
  nand (_03905_, _01234_, _01229_);
  not (_03906_, _03905_);
  not (_03907_, _30964_);
  nor (_03908_, _01229_, _03907_);
  nor (_03909_, _03908_, _03906_);
  nor (_03911_, _03909_, _30592_);
  not (_03912_, _03911_);
  not (_03913_, _01268_);
  not (_03914_, _01421_);
  nor (_03915_, _00245_, _03914_);
  nand (_03916_, _03915_, _01383_);
  nor (_03917_, _03916_, _03780_);
  not (_03918_, _03917_);
  nor (_03919_, _03918_, _30311_);
  not (_03920_, _03919_);
  nor (_03921_, _03920_, _03756_);
  not (_03922_, _03921_);
  nor (_03923_, _03922_, _03743_);
  not (_03924_, _03923_);
  nor (_03925_, _03924_, _03913_);
  not (_03926_, _03925_);
  nor (_03927_, _03926_, _00238_);
  nor (_03928_, _30584_, _03715_);
  nor (_03929_, _03730_, _30300_);
  nand (_03930_, _03929_, _03928_);
  nor (_03931_, _03930_, _03699_);
  nand (_03932_, _03931_, _03927_);
  nor (_03933_, _03932_, _03912_);
  not (_03934_, _03933_);
  nor (_03935_, _03934_, _03690_);
  nor (_03936_, _03933_, _01265_);
  nor (_03937_, _03936_, _03935_);
  not (_03938_, _01263_);
  nor (_03939_, _03690_, _03938_);
  not (_03940_, _03939_);
  nor (_03941_, _03940_, _03932_);
  not (_03942_, _03941_);
  nor (_03943_, _03912_, _03681_);
  nand (_03944_, _03943_, _01488_);
  nor (_03945_, _03944_, _03942_);
  nor (_03946_, _03945_, _03937_);
  nor (_03947_, _03946_, _03904_);
  nand (_03948_, _03904_, _01488_);
  nor (_03949_, _03671_, _30954_);
  not (_03950_, _03949_);
  nor (_03952_, _03950_, _03668_);
  not (_03953_, _03952_);
  nand (_03954_, _03953_, _03948_);
  nor (_03955_, _03954_, _03947_);
  nor (_03956_, _31071_, _27726_);
  not (_03957_, _03956_);
  nor (_03958_, _03957_, _26789_);
  not (_03959_, _03958_);
  nor (_03960_, _03959_, _03668_);
  not (_03961_, _03960_);
  nand (_03962_, _03952_, _03690_);
  nand (_03963_, _03962_, _03961_);
  nor (_03964_, _03963_, _03955_);
  nor (_03965_, _03961_, _28639_);
  nor (_03966_, _03965_, _03964_);
  nor (_04962_, _03966_, _23698_);
  nor (_03967_, _03903_, _01485_);
  not (_03968_, _03927_);
  nor (_03969_, _03968_, _03912_);
  not (_03970_, _03969_);
  nor (_03971_, _03970_, _03930_);
  not (_03972_, _03971_);
  nand (_03973_, _03972_, _01432_);
  nand (_03974_, _03971_, _03699_);
  nand (_03975_, _03974_, _03973_);
  not (_03976_, _03943_);
  nor (_03977_, _03976_, _03697_);
  nand (_03978_, _03977_, _03941_);
  nand (_03979_, _03978_, _03903_);
  nor (_03980_, _03979_, _03975_);
  nor (_03981_, _03980_, _03967_);
  nor (_03982_, _03960_, _03952_);
  nand (_03983_, _03982_, _03981_);
  nand (_03984_, _03952_, _01432_);
  nand (_03985_, _03984_, _03983_);
  nor (_03986_, _03961_, _28598_);
  nor (_03987_, _03986_, _03985_);
  nor (_04998_, _03987_, _23698_);
  nor (_03988_, _03953_, _30300_);
  nor (_03989_, _03970_, _03730_);
  not (_03991_, _03989_);
  nor (_03992_, _03991_, _30584_);
  not (_03993_, _03992_);
  nor (_03994_, _03993_, _03715_);
  nor (_03995_, _03994_, _01291_);
  nor (_03996_, _03995_, _03971_);
  nor (_03997_, _03976_, _03705_);
  nand (_03998_, _03997_, _03941_);
  nand (_03999_, _03998_, _03903_);
  nor (_04000_, _03999_, _03996_);
  nor (_04001_, _03903_, _01482_);
  nor (_04002_, _04001_, _04000_);
  nand (_04003_, _04002_, _03982_);
  nand (_04004_, _03960_, _00800_);
  nand (_04005_, _04004_, _04003_);
  nor (_04006_, _04005_, _03988_);
  nor (_05038_, _04006_, _23698_);
  nor (_04007_, _03953_, _03715_);
  nor (_04008_, _03992_, _01405_);
  nor (_04009_, _04008_, _03994_);
  nor (_04010_, _03976_, _03713_);
  nand (_04011_, _04010_, _03941_);
  nand (_04012_, _04011_, _03903_);
  nor (_04013_, _04012_, _04009_);
  nor (_04014_, _03903_, _01479_);
  nor (_04015_, _04014_, _04013_);
  nand (_04016_, _04015_, _03982_);
  nand (_04017_, _03960_, _27742_);
  nand (_04018_, _04017_, _04016_);
  nor (_04019_, _04018_, _04007_);
  nor (_05103_, _04019_, _23698_);
  not (_04020_, _03982_);
  nand (_04021_, _03904_, _03721_);
  nand (_04022_, _03991_, _30584_);
  nand (_04023_, _04022_, _03993_);
  nand (_04024_, _03943_, _01476_);
  nor (_04025_, _04024_, _03942_);
  nor (_04026_, _04025_, _03904_);
  nand (_04027_, _04026_, _04023_);
  nand (_04028_, _04027_, _04021_);
  nor (_04031_, _04028_, _04020_);
  nand (_04032_, _03960_, _00811_);
  nand (_04033_, _03952_, _01409_);
  nand (_04034_, _04033_, _04032_);
  nor (_04035_, _04034_, _04031_);
  nor (_05169_, _04035_, _23698_);
  nor (_04036_, _03969_, _01412_);
  nor (_04037_, _04036_, _03989_);
  nor (_04038_, _04037_, _03904_);
  nor (_04039_, _03976_, _03728_);
  nand (_04040_, _04039_, _03941_);
  nand (_04041_, _04040_, _04038_);
  nand (_04042_, _03904_, _03728_);
  nand (_04043_, _04042_, _04041_);
  nor (_04044_, _04043_, _04020_);
  nand (_04045_, _03960_, _28244_);
  nand (_04046_, _03952_, _01412_);
  nand (_04047_, _04046_, _04045_);
  nor (_04048_, _04047_, _04044_);
  nor (_05210_, _04048_, _23698_);
  not (_04049_, _01469_);
  nor (_04050_, _03976_, _04049_);
  nand (_04051_, _04050_, _03941_);
  nor (_04052_, _03926_, _03912_);
  nor (_04053_, _04052_, _01295_);
  nor (_04054_, _04053_, _03969_);
  nor (_04055_, _04054_, _03904_);
  nand (_04056_, _04055_, _04051_);
  nand (_04057_, _03904_, _04049_);
  nand (_04058_, _04057_, _04056_);
  nor (_04059_, _04058_, _03952_);
  nand (_04060_, _03952_, _01295_);
  nand (_04061_, _04060_, _03961_);
  nor (_04062_, _04061_, _04059_);
  nand (_04063_, _03960_, _27888_);
  nand (_04064_, _04063_, _29344_);
  nor (_05250_, _04064_, _04062_);
  nor (_04065_, _03953_, _28639_);
  nor (_04066_, _03976_, _03741_);
  nand (_04067_, _04066_, _03941_);
  nand (_04069_, _03921_, _03911_);
  nor (_04070_, _04069_, _01369_);
  nand (_04071_, _04069_, _01369_);
  nand (_04072_, _04071_, _03903_);
  nor (_04073_, _04072_, _04070_);
  nand (_04074_, _04073_, _04067_);
  nor (_04075_, _03903_, _01459_);
  nor (_04076_, _04075_, _03952_);
  nand (_04077_, _04076_, _04074_);
  nand (_04078_, _04077_, _03961_);
  nor (_04079_, _04078_, _04065_);
  nand (_04080_, _03960_, _03743_);
  nand (_04081_, _04080_, _29344_);
  nor (_05288_, _04081_, _04079_);
  nor (_04082_, _03953_, _28598_);
  nor (_04083_, _03903_, _01456_);
  nand (_04084_, _03943_, _01456_);
  nor (_04085_, _04084_, _03942_);
  nand (_04086_, _03919_, _03911_);
  nand (_04087_, _04086_, _03756_);
  nand (_04088_, _04087_, _04069_);
  nand (_04089_, _04088_, _03903_);
  nor (_04090_, _04089_, _04085_);
  nor (_04091_, _04090_, _04083_);
  nand (_04092_, _04091_, _03953_);
  nand (_04093_, _04092_, _03961_);
  nor (_04094_, _04093_, _04082_);
  nand (_04095_, _03960_, _03756_);
  nand (_04096_, _04095_, _29344_);
  nor (_05328_, _04096_, _04094_);
  nand (_04097_, _03943_, _01453_);
  nor (_04098_, _04097_, _03942_);
  nand (_04099_, _03917_, _03911_);
  nand (_04100_, _04099_, _30311_);
  nand (_04101_, _04100_, _04086_);
  nand (_04102_, _04101_, _03903_);
  nor (_04103_, _04102_, _04098_);
  nand (_04104_, _03904_, _30298_);
  nand (_04105_, _04104_, _03953_);
  nor (_04106_, _04105_, _04103_);
  nor (_04108_, _03953_, _27584_);
  nor (_04109_, _04108_, _04106_);
  nor (_04110_, _04109_, _03960_);
  nor (_04111_, _03961_, _30311_);
  nor (_04112_, _04111_, _04110_);
  nor (_05378_, _04112_, _23698_);
  nor (_04113_, _03953_, _27718_);
  nor (_04114_, _03903_, _01450_);
  nand (_04115_, _03943_, _01450_);
  nor (_04116_, _04115_, _03942_);
  not (_04117_, _03916_);
  nand (_04118_, _04117_, _03911_);
  nand (_04119_, _04118_, _03780_);
  nand (_04120_, _04119_, _04099_);
  nand (_04121_, _04120_, _03903_);
  nor (_04122_, _04121_, _04116_);
  nor (_04123_, _04122_, _04114_);
  nand (_04124_, _04123_, _03953_);
  nand (_04125_, _04124_, _03961_);
  nor (_04126_, _04125_, _04113_);
  nand (_04127_, _03960_, _03780_);
  nand (_04128_, _04127_, _29344_);
  nor (_05434_, _04128_, _04126_);
  nand (_04129_, _03943_, _01447_);
  nor (_04130_, _04129_, _03942_);
  nand (_04131_, _03915_, _03911_);
  nand (_04132_, _04131_, _30595_);
  nand (_04133_, _04132_, _04118_);
  nand (_04134_, _04133_, _03903_);
  nor (_04135_, _04134_, _04130_);
  nand (_04136_, _03904_, _30581_);
  nand (_04137_, _04136_, _03953_);
  nor (_04138_, _04137_, _04135_);
  nor (_04139_, _03953_, _28540_);
  nor (_04140_, _04139_, _04138_);
  nor (_04141_, _04140_, _03960_);
  nor (_04142_, _03961_, _30595_);
  nor (_04143_, _04142_, _04141_);
  nor (_05488_, _04143_, _23698_);
  nand (_04144_, _03943_, _01444_);
  nor (_04146_, _04144_, _03942_);
  nand (_04147_, _03911_, _01423_);
  nand (_04148_, _04147_, _03914_);
  nand (_04149_, _04148_, _04131_);
  nand (_04150_, _04149_, _03903_);
  nor (_04151_, _04150_, _04146_);
  nand (_04152_, _03904_, _03890_);
  nand (_04153_, _04152_, _03953_);
  nor (_04154_, _04153_, _04151_);
  nand (_04155_, _03952_, _28244_);
  nand (_04156_, _04155_, _03961_);
  nor (_04157_, _04156_, _04154_);
  nand (_04158_, _03960_, _03914_);
  nand (_04159_, _04158_, _29344_);
  nor (_05522_, _04159_, _04157_);
  nor (_04160_, _03911_, _01423_);
  nand (_04161_, _03682_, _01441_);
  nor (_04162_, _04161_, _03942_);
  nor (_04163_, _04162_, _04147_);
  nor (_04164_, _04163_, _04160_);
  nor (_04165_, _04164_, _03904_);
  nand (_04166_, _03904_, _00235_);
  nand (_04167_, _04166_, _03953_);
  nor (_04168_, _04167_, _04165_);
  nand (_04169_, _03952_, _27886_);
  nand (_04170_, _04169_, _03961_);
  nor (_04171_, _04170_, _04168_);
  nand (_04172_, _03960_, _00245_);
  nand (_04173_, _04172_, _29344_);
  nor (_05559_, _04173_, _04171_);
  nand (_04174_, _31258_, _30944_);
  nand (_04175_, _31259_, _01345_);
  nand (_04176_, _04175_, _04174_);
  nor (_04177_, _04176_, _03798_);
  nand (_04178_, _00438_, _03801_);
  nor (_04179_, _04178_, _03800_);
  nor (_04180_, _04179_, _04177_);
  nor (_04181_, _04180_, _03820_);
  nand (_04182_, _03820_, _28481_);
  nand (_04183_, _04182_, _29344_);
  nor (_05600_, _04183_, _04181_);
  nor (_04185_, _03902_, _03680_);
  nand (_04186_, _04185_, _03911_);
  nor (_04187_, _04186_, _03942_);
  nor (_04188_, _04187_, _04020_);
  nand (_04189_, _04020_, _03801_);
  nand (_04190_, _04189_, _29344_);
  nor (_05647_, _04190_, _04188_);
  nor (_04191_, _03961_, _28482_);
  nor (_04192_, _03935_, _01263_);
  nand (_04193_, _03682_, _01307_);
  nand (_04194_, _04193_, _03911_);
  nor (_04195_, _04194_, _03942_);
  nor (_04196_, _04195_, _04192_);
  nor (_04197_, _04196_, _03904_);
  not (_04198_, _01307_);
  nand (_04199_, _03904_, _04198_);
  nand (_04200_, _04199_, _03953_);
  nor (_04201_, _04200_, _04197_);
  nor (_04202_, _03953_, _03938_);
  nor (_04203_, _04202_, _04201_);
  nand (_04204_, _04203_, _03961_);
  nand (_04205_, _04204_, _29344_);
  nor (_05686_, _04205_, _04191_);
  nor (_04206_, _03953_, _28481_);
  not (_04207_, _01303_);
  nor (_04208_, _03976_, _04207_);
  nand (_04209_, _04208_, _03941_);
  nor (_04210_, _03924_, _03912_);
  nor (_04211_, _04210_, _01268_);
  nor (_04212_, _04211_, _04052_);
  nor (_04213_, _04212_, _03904_);
  nand (_04214_, _04213_, _04209_);
  nor (_04215_, _03903_, _01303_);
  nor (_04216_, _04215_, _03952_);
  nand (_04217_, _04216_, _04214_);
  nand (_04218_, _04217_, _03961_);
  nor (_04219_, _04218_, _04206_);
  nand (_04220_, _03960_, _03913_);
  nand (_04221_, _04220_, _29344_);
  nor (_05726_, _04221_, _04219_);
  not (_04223_, _06028_);
  nand (_04224_, _01299_, _04223_);
  nor (_05766_, _04224_, _23698_);
  nor (_04225_, _03912_, _03679_);
  nand (_04226_, _04225_, _03982_);
  nor (_04227_, _04226_, _03941_);
  not (_04228_, _00839_);
  nand (_04229_, _04226_, _04228_);
  nand (_04230_, _04229_, _29344_);
  nor (_05804_, _04230_, _04227_);
  nor (_04231_, _03675_, _28482_);
  nand (_04232_, _03688_, _03938_);
  nand (_04233_, _03691_, _04198_);
  nand (_04234_, _04233_, _04232_);
  nand (_04235_, _04234_, _03675_);
  nand (_04236_, _04235_, _29344_);
  nor (_05842_, _04236_, _04231_);
  nor (_04237_, _03748_, _28482_);
  nor (_04238_, _03683_, _04207_);
  nor (_04239_, _03684_, _03913_);
  nor (_04240_, _04239_, _04238_);
  nand (_04241_, _04240_, _03748_);
  nand (_04242_, _04241_, _03675_);
  nor (_04243_, _04242_, _04237_);
  nor (_04244_, _03675_, _04207_);
  nor (_04245_, _04244_, _04243_);
  nor (_05881_, _04245_, _23698_);
  not (_04246_, _01284_);
  nand (_04247_, _01287_, _04246_);
  nor (_05929_, _04247_, _23698_);
  nor (_05980_, _04246_, _23698_);
  nor (_06018_, _04223_, _23698_);
  not (_04248_, _00961_);
  not (_04249_, _00963_);
  nor (_04250_, _04249_, _04248_);
  not (_04251_, _04250_);
  not (_04252_, _00847_);
  not (_04253_, _00806_);
  nor (_04254_, _00916_, _00801_);
  nor (_04256_, _04254_, _04253_);
  nand (_04257_, _04256_, _00810_);
  nor (_04258_, _04257_, _04252_);
  not (_04259_, _04258_);
  nor (_04260_, _04259_, _04251_);
  nor (_04261_, _04260_, _00953_);
  not (_04262_, _00953_);
  nor (_04263_, _04251_, _04262_);
  nor (_04264_, _04263_, _04257_);
  not (_04265_, _04257_);
  nand (_04266_, _00810_, _00784_);
  nor (_04267_, _04266_, _04254_);
  nor (_04268_, _04267_, _04265_);
  nor (_04269_, _04268_, _04252_);
  not (_04270_, _04269_);
  nor (_04271_, _04270_, _04264_);
  nor (_04272_, _04271_, _23698_);
  not (_04273_, _04272_);
  nor (_06070_, _04273_, _04261_);
  not (_04274_, _27953_);
  nor (_04275_, _26683_, _04274_);
  nor (_04276_, _00795_, _26789_);
  nand (_04277_, _04276_, _04275_);
  not (_04278_, _04277_);
  not (_04279_, _00947_);
  not (_04280_, _00776_);
  not (_04281_, _04254_);
  nand (_04282_, _04281_, _00791_);
  nor (_04283_, _04282_, _04280_);
  not (_04284_, _00971_);
  not (_04285_, _00973_);
  nor (_04286_, _04285_, _04284_);
  nand (_04287_, _04286_, _04283_);
  nand (_04288_, _04287_, _04279_);
  nor (_04289_, _04287_, _04279_);
  nor (_04290_, _04289_, _23698_);
  nand (_04291_, _04290_, _04288_);
  nor (_06112_, _04291_, _04278_);
  nor (_04292_, _27610_, _26679_);
  not (_04293_, _04292_);
  nor (_04295_, _29299_, _04293_);
  not (_04296_, _04295_);
  nor (_04297_, _04296_, _00768_);
  not (_04298_, _04297_);
  nor (_04299_, _04298_, _31182_);
  not (_04300_, _04299_);
  nor (_04301_, _04300_, _30944_);
  nor (_04302_, _04299_, _00801_);
  nor (_04303_, _04302_, _04301_);
  not (_04304_, _04275_);
  nor (_04305_, _04304_, _03818_);
  nor (_04306_, _04305_, _04303_);
  nand (_04307_, _04305_, _28639_);
  nand (_04308_, _04307_, _29344_);
  nor (_06161_, _04308_, _04306_);
  nand (_04309_, _04283_, _00973_);
  nand (_04310_, _04309_, _04284_);
  not (_04311_, _04287_);
  nor (_04312_, _04311_, _23698_);
  nand (_04313_, _04312_, _04310_);
  nor (_06206_, _04313_, _04278_);
  nand (_04314_, _04297_, _31070_);
  nor (_04315_, _04314_, _30944_);
  not (_04316_, _04305_);
  nand (_04317_, _04314_, _00506_);
  nand (_04318_, _04317_, _04316_);
  nor (_04319_, _04318_, _04315_);
  nor (_04320_, _04316_, _28598_);
  nor (_04321_, _04320_, _04319_);
  nor (_06246_, _04321_, _23698_);
  nand (_04322_, _04297_, _30953_);
  nor (_04323_, _04322_, _30944_);
  nand (_04324_, _04322_, _00514_);
  nand (_04325_, _04324_, _04316_);
  nor (_04326_, _04325_, _04323_);
  nor (_04327_, _04316_, _27584_);
  nor (_04328_, _04327_, _04326_);
  nor (_06283_, _04328_, _23698_);
  nor (_04329_, _00847_, _23698_);
  nand (_04330_, _04329_, _01016_);
  nor (_04332_, _04252_, _23698_);
  nand (_04333_, _04332_, _01018_);
  nand (_06324_, _04333_, _04330_);
  nand (_04334_, _04329_, _01013_);
  nand (_04335_, _04332_, _01015_);
  nand (_06366_, _04335_, _04334_);
  nor (_04336_, _04283_, _00973_);
  nor (_04337_, _04336_, _23698_);
  nand (_04338_, _04337_, _04309_);
  nor (_06417_, _04338_, _04278_);
  nor (_04339_, _04270_, _04249_);
  nand (_04341_, _04259_, _04249_);
  nand (_04343_, _04341_, _29344_);
  nor (_06463_, _04343_, _04339_);
  nand (_04345_, _04297_, _00104_);
  nor (_04346_, _04345_, _30944_);
  not (_04347_, _00941_);
  nand (_04348_, _04345_, _04347_);
  nand (_04350_, _04348_, _04316_);
  nor (_04351_, _04350_, _04346_);
  nor (_04352_, _04316_, _27718_);
  nor (_04353_, _04352_, _04351_);
  nor (_06514_, _04353_, _23698_);
  nor (_04354_, _00092_, _30943_);
  nand (_04355_, _00092_, _00929_);
  nand (_04356_, _04355_, _04297_);
  nor (_04357_, _04356_, _04354_);
  nor (_04359_, _00894_, _00847_);
  nand (_04360_, _04359_, _04281_);
  not (_04362_, _04360_);
  nand (_04363_, _04362_, _00765_);
  nand (_04364_, _04360_, _00929_);
  nand (_04365_, _04364_, _04363_);
  nor (_04366_, _04365_, _04297_);
  nor (_04367_, _04366_, _04357_);
  nor (_04369_, _04367_, _04305_);
  nand (_04370_, _04305_, _28540_);
  nand (_04372_, _04370_, _29344_);
  nor (_06575_, _04372_, _04369_);
  nor (_04373_, _04269_, _04248_);
  nand (_04375_, _04249_, _04248_);
  nand (_04377_, _04375_, _04251_);
  nor (_04378_, _04377_, _04259_);
  nor (_04379_, _04378_, _04373_);
  nor (_06635_, _04379_, _23698_);
  not (_04380_, _00869_);
  nand (_04381_, _04263_, _04380_);
  nor (_04382_, _04381_, _04259_);
  nor (_04383_, _04382_, _00859_);
  not (_04384_, _00813_);
  nand (_04385_, _04382_, _04384_);
  nand (_04387_, _04385_, _29344_);
  nor (_06676_, _04387_, _04383_);
  nor (_04389_, _00818_, _00514_);
  nand (_04391_, _04389_, _04253_);
  nor (_04392_, _04391_, _04281_);
  nor (_04393_, _04392_, _04267_);
  nor (_04394_, _04393_, _04265_);
  not (_04395_, _01042_);
  nor (_04396_, _04281_, _04253_);
  not (_04397_, _04396_);
  nor (_04398_, _04397_, _03907_);
  nor (_04399_, _04249_, _00961_);
  nor (_04400_, _00953_, _04380_);
  nand (_04401_, _04400_, _04399_);
  nor (_04402_, _04401_, _04257_);
  nor (_04403_, _04402_, _04398_);
  nand (_04404_, _04403_, _04395_);
  nor (_04405_, _04404_, _04394_);
  not (_04406_, _04329_);
  nor (_04407_, _04406_, _04395_);
  not (_04408_, _04332_);
  nor (_04409_, _04403_, _01013_);
  nor (_04410_, _04409_, _04408_);
  nor (_04411_, _04410_, _04407_);
  nor (_06718_, _04411_, _04405_);
  nand (_04413_, _04329_, _00877_);
  not (_04415_, _04403_);
  nand (_04416_, _04415_, _00765_);
  not (_04418_, _04394_);
  not (_04421_, _00877_);
  nor (_04422_, _04415_, _04421_);
  nand (_04423_, _04422_, _04418_);
  nand (_04424_, _04423_, _04416_);
  nand (_04425_, _04424_, _04332_);
  nand (_06759_, _04425_, _04413_);
  nand (_04426_, _04329_, _01034_);
  nand (_04427_, _04415_, _00877_);
  not (_04428_, _01034_);
  nor (_04429_, _04415_, _04428_);
  nand (_04430_, _04429_, _04418_);
  nand (_04431_, _04430_, _04427_);
  nand (_04432_, _04431_, _04332_);
  nand (_06800_, _04432_, _04426_);
  not (_04433_, _00894_);
  nand (_04434_, _00509_, _04433_);
  nor (_04435_, _04434_, _04297_);
  nand (_04436_, _31399_, _00920_);
  nand (_04437_, _04436_, _04297_);
  nor (_04438_, _04437_, _31400_);
  nor (_04439_, _04438_, _04435_);
  nor (_04440_, _04439_, _04305_);
  nand (_04441_, _04305_, _28157_);
  nand (_04443_, _04441_, _29344_);
  nor (_06841_, _04443_, _04440_);
  nor (_04444_, _30944_, _26895_);
  nand (_04445_, _26895_, _00516_);
  nand (_04446_, _04445_, _04297_);
  nor (_04447_, _04446_, _04444_);
  nor (_04448_, _00765_, _00506_);
  nand (_04450_, _04448_, _04281_);
  nand (_04451_, _04450_, _04359_);
  nand (_04452_, _04451_, _00516_);
  nand (_04453_, _04452_, _04298_);
  nand (_04454_, _04453_, _04316_);
  nor (_04455_, _04454_, _04447_);
  nand (_04456_, _04305_, _27888_);
  nand (_04457_, _04456_, _29344_);
  nor (_06882_, _04457_, _04455_);
  nand (_04459_, _00778_, _27977_);
  nor (_04461_, _04459_, _00828_);
  not (_04462_, _01197_);
  nand (_04463_, _04459_, _04462_);
  nand (_04464_, _04463_, _29344_);
  nor (_06923_, _04464_, _04461_);
  nor (_04465_, _04459_, _00750_);
  not (_04467_, _01195_);
  nand (_04468_, _04459_, _04467_);
  nand (_04470_, _04468_, _29344_);
  nor (_06966_, _04470_, _04465_);
  nor (_04472_, _04459_, _00800_);
  not (_04474_, _01193_);
  nand (_04475_, _04459_, _04474_);
  nand (_04476_, _04475_, _29344_);
  nor (_07008_, _04476_, _04472_);
  nand (_04477_, _04329_, _01030_);
  nand (_04478_, _04415_, _01034_);
  not (_04479_, _01030_);
  nor (_04480_, _04392_, _04265_);
  nand (_04481_, _04480_, _04267_);
  nand (_04482_, _04481_, _04479_);
  not (_04483_, _04401_);
  nor (_04484_, _04483_, _04257_);
  nor (_04485_, _04484_, _04480_);
  nor (_04486_, _04485_, _04398_);
  nand (_04487_, _04486_, _04482_);
  nand (_04488_, _04487_, _04478_);
  nand (_04489_, _04488_, _04332_);
  nand (_07050_, _04489_, _04477_);
  nor (_04490_, _04459_, _27742_);
  not (_04491_, _01191_);
  nand (_04492_, _04459_, _04491_);
  nand (_04493_, _04492_, _29344_);
  nor (_07091_, _04493_, _04490_);
  nor (_04494_, _04459_, _00811_);
  nand (_04495_, _04459_, _30630_);
  nand (_04496_, _04495_, _29344_);
  nor (_07132_, _04496_, _04494_);
  nand (_04497_, _04329_, _01027_);
  not (_04498_, _01027_);
  nand (_04500_, _04418_, _04498_);
  nand (_04501_, _04500_, _04403_);
  nand (_04502_, _04415_, _01030_);
  nand (_04503_, _04502_, _04501_);
  nand (_04504_, _04503_, _04332_);
  nand (_07161_, _04504_, _04497_);
  nand (_04505_, _04329_, _01023_);
  nor (_04506_, _04394_, _01023_);
  nand (_04507_, _04506_, _04403_);
  nor (_04508_, _04403_, _01027_);
  nor (_04509_, _04508_, _04408_);
  nand (_04511_, _04509_, _04507_);
  nand (_07196_, _04511_, _04505_);
  nor (_04512_, _04459_, _28244_);
  not (_04513_, _01187_);
  nand (_04515_, _04459_, _04513_);
  nand (_04516_, _04515_, _29344_);
  nor (_07230_, _04516_, _04512_);
  nor (_04517_, _04459_, _27886_);
  nand (_04518_, _04459_, _00273_);
  nand (_04519_, _04518_, _29344_);
  nor (_07269_, _04519_, _04517_);
  not (_04520_, _00904_);
  nor (_04521_, _04280_, _03907_);
  nand (_04522_, _04521_, _04254_);
  not (_04523_, _04522_);
  not (_04524_, _04283_);
  nor (_04525_, _00973_, _00971_);
  nor (_04526_, _00947_, _00900_);
  nand (_04527_, _04526_, _04525_);
  nor (_04528_, _04527_, _04524_);
  nor (_04529_, _04528_, _04523_);
  nor (_04530_, _04529_, _04520_);
  not (_04531_, _00978_);
  not (_04532_, _04529_);
  nor (_04533_, _04532_, _04531_);
  nor (_04534_, _04533_, _04530_);
  nor (_04535_, _04534_, _04278_);
  nand (_04536_, _04347_, _00916_);
  nand (_04537_, _04536_, _04281_);
  nor (_04539_, _04537_, _04277_);
  nor (_04540_, _04539_, _04535_);
  nor (_07307_, _04540_, _23698_);
  nor (_04541_, _04277_, _04254_);
  not (_04542_, _04541_);
  nor (_04543_, _04542_, _28482_);
  not (_04544_, _00981_);
  nand (_04545_, _04529_, _04544_);
  nand (_04546_, _04532_, _04531_);
  nand (_04547_, _04546_, _04545_);
  nand (_04548_, _04547_, _04277_);
  nand (_04549_, _04548_, _29344_);
  nor (_07346_, _04549_, _04543_);
  nor (_04550_, _04277_, _00916_);
  nand (_04551_, _04550_, _00521_);
  nor (_04552_, _04551_, _28481_);
  nand (_04553_, _04532_, _00981_);
  nand (_04554_, _04529_, _00983_);
  nand (_04555_, _04554_, _04553_);
  nand (_04556_, _04555_, _04277_);
  nand (_04557_, _04541_, _00828_);
  nand (_04558_, _04557_, _04556_);
  nor (_04559_, _04558_, _04552_);
  nor (_07383_, _04559_, _23698_);
  nor (_04560_, _04277_, _04281_);
  not (_04561_, _04560_);
  nor (_04562_, _04561_, _28639_);
  nand (_04563_, _04541_, _00750_);
  nand (_04564_, _04532_, _00983_);
  nand (_04565_, _04529_, _00985_);
  nand (_04566_, _04565_, _04564_);
  nand (_04567_, _04566_, _04277_);
  nand (_04568_, _04567_, _04563_);
  nor (_04569_, _04568_, _04562_);
  nor (_07423_, _04569_, _23698_);
  nor (_04570_, _04551_, _28598_);
  nand (_04571_, _04532_, _00985_);
  nand (_04572_, _04529_, _00988_);
  nand (_04573_, _04572_, _04571_);
  nand (_04574_, _04573_, _04277_);
  nand (_04576_, _04541_, _00800_);
  nand (_04577_, _04576_, _04574_);
  nor (_04578_, _04577_, _04570_);
  nor (_07461_, _04578_, _23698_);
  not (_04579_, _01039_);
  nand (_04580_, _04403_, _04579_);
  nor (_04581_, _04580_, _04394_);
  nor (_04582_, _04406_, _04579_);
  nor (_04583_, _04403_, _01042_);
  nor (_04584_, _04583_, _04408_);
  nor (_04585_, _04584_, _04582_);
  nor (_07498_, _04585_, _04581_);
  nand (_04586_, _04329_, _01020_);
  nor (_04587_, _04394_, _01020_);
  nand (_04588_, _04587_, _04403_);
  nor (_04589_, _04403_, _01023_);
  nor (_04590_, _04589_, _04408_);
  nand (_04591_, _04590_, _04588_);
  nand (_07537_, _04591_, _04586_);
  nor (_04592_, _04394_, _01016_);
  nand (_04593_, _04592_, _04403_);
  nor (_04594_, _04403_, _01020_);
  nor (_04595_, _04594_, _04408_);
  nand (_04596_, _04595_, _04593_);
  nand (_07583_, _04596_, _04330_);
  nor (_04597_, _04394_, _01013_);
  nand (_04598_, _04597_, _04403_);
  nor (_04599_, _04403_, _01016_);
  nor (_04600_, _04599_, _04408_);
  nand (_04601_, _04600_, _04598_);
  nand (_07623_, _04601_, _04334_);
  nor (_04602_, _04551_, _27584_);
  nand (_04603_, _04532_, _00988_);
  nand (_04604_, _04529_, _00990_);
  nand (_04605_, _04604_, _04603_);
  nand (_04606_, _04605_, _04277_);
  nand (_04607_, _04541_, _27742_);
  nand (_04608_, _04607_, _04606_);
  nor (_04609_, _04608_, _04602_);
  nor (_07664_, _04609_, _23698_);
  nor (_04611_, _04551_, _27718_);
  nand (_04612_, _04532_, _00990_);
  nand (_04613_, _04529_, _00992_);
  nand (_04614_, _04613_, _04612_);
  nand (_04615_, _04614_, _04277_);
  nand (_04616_, _04541_, _00811_);
  nand (_04618_, _04616_, _04615_);
  nor (_04619_, _04618_, _04611_);
  nor (_07707_, _04619_, _23698_);
  nor (_04620_, _04551_, _28540_);
  nand (_04621_, _04532_, _00992_);
  nand (_04622_, _04529_, _00995_);
  nand (_04623_, _04622_, _04621_);
  nand (_04624_, _04623_, _04277_);
  nand (_04625_, _04541_, _28244_);
  nand (_04626_, _04625_, _04624_);
  nor (_04627_, _04626_, _04620_);
  nor (_07752_, _04627_, _23698_);
  nand (_04628_, _04532_, _00995_);
  nand (_04629_, _04529_, _00996_);
  nand (_04630_, _04629_, _04628_);
  nand (_04631_, _04630_, _04277_);
  nand (_04632_, _04541_, _27886_);
  nand (_04633_, _04632_, _04631_);
  nor (_04634_, _04561_, _28157_);
  nor (_04635_, _04634_, _04633_);
  nor (_07795_, _04635_, _23698_);
  nor (_04638_, _30997_, _30995_);
  nor (_04639_, _04638_, _00264_);
  not (_04640_, _04639_);
  nor (_04641_, _04640_, _00841_);
  not (_04642_, _00916_);
  nor (_04643_, _04642_, _00801_);
  nor (_04644_, _00431_, _04228_);
  nor (_04645_, _04644_, _04643_);
  not (_04646_, _04645_);
  nor (_04647_, _04646_, _04641_);
  not (_04648_, _00831_);
  not (_04649_, _00834_);
  nand (_04650_, _04649_, _04648_);
  nand (_04652_, _04650_, _29344_);
  nor (_07841_, _04652_, _04647_);
  nand (_04653_, _04382_, _29344_);
  nand (_04654_, _04272_, _00869_);
  nand (_07887_, _04654_, _04653_);
  nand (_04655_, _04332_, _01025_);
  nand (_07933_, _04655_, _04505_);
  nand (_04656_, _04332_, _01029_);
  nand (_07974_, _04656_, _04497_);
  nand (_04657_, _04332_, _01032_);
  nand (_08024_, _04657_, _04477_);
  nand (_04659_, _04297_, _31258_);
  nor (_04661_, _04659_, _30944_);
  nand (_04662_, _04659_, _04642_);
  nand (_04663_, _04662_, _04316_);
  nor (_04664_, _04663_, _04661_);
  nor (_04665_, _04316_, _28481_);
  nor (_04667_, _04665_, _04664_);
  nor (_08072_, _04667_, _23698_);
  nor (_04668_, _04459_, _28482_);
  nand (_04669_, _04459_, _04649_);
  nand (_04670_, _04669_, _29344_);
  nor (_08114_, _04670_, _04668_);
  nor (_04671_, _04532_, _04520_);
  nor (_04672_, _04671_, _04278_);
  not (_04673_, _04550_);
  nand (_04674_, _04673_, _29344_);
  nor (_08156_, _04674_, _04672_);
  nor (_04675_, _04375_, _04259_);
  nand (_04676_, _04675_, _04400_);
  nor (_04677_, _04676_, _00813_);
  not (_04679_, _00814_);
  nand (_04681_, _04676_, _04679_);
  nand (_04683_, _04681_, _29344_);
  nor (_08199_, _04683_, _04677_);
  nand (_04685_, _04332_, _01036_);
  nand (_08243_, _04685_, _04426_);
  nand (_04687_, _04289_, _00900_);
  nor (_04688_, _04289_, _00900_);
  nor (_04690_, _04688_, _23698_);
  nand (_04692_, _04690_, _04687_);
  nor (_08288_, _04692_, _04278_);
  not (_04694_, _00848_);
  nand (_04695_, _04403_, _04694_);
  nor (_04697_, _04695_, _04394_);
  nor (_04698_, _04406_, _04694_);
  nor (_04699_, _04403_, _01039_);
  nor (_04700_, _04699_, _04408_);
  nor (_04701_, _04700_, _04698_);
  nor (_08332_, _04701_, _04697_);
  nand (_04702_, _04332_, _01022_);
  nand (_08378_, _04702_, _04586_);
  nand (_04703_, _04523_, _00996_);
  nor (_04704_, _00996_, _00995_);
  nor (_04705_, _00978_, _00904_);
  nor (_04706_, _00983_, _00981_);
  nand (_04707_, _04706_, _04705_);
  nor (_04708_, _00992_, _00990_);
  nor (_04709_, _00988_, _00985_);
  nand (_04710_, _04709_, _04708_);
  nor (_04711_, _04710_, _04707_);
  nand (_04712_, _04711_, _04704_);
  nor (_04713_, _04712_, _04522_);
  nand (_04714_, _04713_, _01000_);
  nand (_04715_, _04714_, _04703_);
  nand (_04716_, _04528_, _00996_);
  not (_04718_, _04528_);
  not (_04719_, _01000_);
  nor (_04721_, _04523_, _04719_);
  nand (_04722_, _04721_, _04718_);
  nand (_04723_, _04722_, _04716_);
  nor (_04725_, _04723_, _04715_);
  nor (_04726_, _04725_, _04278_);
  nor (_04727_, _04561_, _27888_);
  nor (_04729_, _04727_, _04726_);
  nor (_08444_, _04729_, _23698_);
  nor (_04730_, _04527_, _01000_);
  not (_04732_, _04730_);
  nor (_04733_, _04732_, _04712_);
  not (_04734_, _04527_);
  nor (_04737_, _04734_, _04433_);
  nor (_04738_, _04737_, _04733_);
  nor (_04739_, _04738_, _04524_);
  nand (_04741_, _04282_, _00776_);
  nor (_04742_, _04741_, _04433_);
  nor (_04743_, _04742_, _04739_);
  nor (_04745_, _04743_, _04523_);
  nor (_04746_, _04745_, _04713_);
  nand (_04747_, _04277_, _29344_);
  nor (_08508_, _04747_, _04746_);
  nor (_04749_, _04647_, _00834_);
  nor (_04750_, _04749_, _00831_);
  nand (_04752_, _04749_, _00831_);
  nand (_04753_, _04752_, _29344_);
  nor (_08572_, _04753_, _04750_);
  nand (_04755_, _04332_, _00878_);
  nand (_08616_, _04755_, _04413_);
  not (_04756_, _04282_);
  nand (_04758_, _04733_, _04756_);
  nand (_04759_, _04758_, _00776_);
  nor (_04760_, _04759_, _04713_);
  nor (_04762_, _04760_, _04278_);
  nor (_08657_, _04762_, _23698_);
  not (_04763_, _00824_);
  nor (_04765_, _04763_, _00813_);
  nor (_04766_, _04765_, _04266_);
  nor (_04767_, _04267_, _04256_);
  nor (_04769_, _04767_, _04766_);
  nand (_04770_, _04480_, _04397_);
  nor (_04771_, _04770_, _04769_);
  nor (_08698_, _04771_, _04408_);
  nor (_04773_, _04408_, _00848_);
  nand (_08750_, _04773_, _04415_);
  nor (_04775_, _00810_, _00514_);
  nand (_04776_, _04281_, _00847_);
  nor (_04777_, _04776_, _04775_);
  nand (_04779_, _04777_, _04257_);
  nand (_04780_, _04779_, _00824_);
  nor (_04781_, _04779_, _04384_);
  nor (_04783_, _04781_, _23698_);
  nand (_08792_, _04783_, _04780_);
  nor (_04785_, _04640_, _00888_);
  nor (_04787_, _30307_, _04228_);
  nor (_04788_, _04787_, _04643_);
  not (_04789_, _04788_);
  nor (_04791_, _04789_, _04785_);
  nor (_04792_, _00834_, _00803_);
  nor (_04793_, _04792_, _04791_);
  nor (_04795_, _04793_, _04791_);
  nor (_04796_, _04795_, _00803_);
  nand (_04797_, _04793_, _04649_);
  nand (_04799_, _04797_, _29344_);
  nor (_08845_, _04799_, _04796_);
  not (_04800_, _04793_);
  nor (_08897_, _04800_, _23698_);
  not (_04802_, _00765_);
  nand (_04803_, _04252_, _04802_);
  nand (_04804_, _04803_, _29344_);
  nand (_04805_, _04398_, _00813_);
  nand (_04806_, _00859_, _00813_);
  not (_04807_, _00859_);
  nand (_04808_, _04807_, _04384_);
  nand (_04809_, _04808_, _00814_);
  nand (_04810_, _04809_, _04806_);
  nand (_04812_, _04810_, _04402_);
  nand (_04813_, _04812_, _04805_);
  nor (_04815_, _04415_, _04394_);
  nor (_04816_, _04815_, _04252_);
  nor (_04818_, _04816_, _04802_);
  nor (_04819_, _04818_, _04813_);
  nor (_08959_, _04819_, _04804_);
  not (_04821_, _00417_);
  nand (_04822_, _00318_, _00201_);
  not (_04823_, _04822_);
  nor (_04824_, _04823_, _04821_);
  not (_04825_, _04824_);
  not (_04826_, _00201_);
  not (_04827_, _00627_);
  nor (_04828_, _04827_, _04821_);
  not (_04829_, _00641_);
  nor (_04832_, _04829_, _00417_);
  nor (_04833_, _04832_, _00624_);
  not (_04834_, _04833_);
  nor (_04835_, _04834_, _04828_);
  nor (_04836_, _04835_, _04826_);
  not (_04837_, _04836_);
  not (_04838_, _00204_);
  not (_04839_, _00207_);
  nor (_04840_, _01345_, _01249_);
  nor (_04841_, _04840_, _04839_);
  not (_04842_, _04841_);
  nor (_04843_, _04842_, _04838_);
  nor (_04844_, _00920_, _00818_);
  nor (_04845_, _04844_, _30287_);
  not (_04846_, _04845_);
  nor (_04847_, _04846_, _30291_);
  nor (_04848_, _04847_, _04843_);
  nor (_04849_, _00598_, _00226_);
  not (_04850_, _04849_);
  nor (_04851_, _04850_, _00228_);
  not (_04852_, _04851_);
  not (_04853_, _00435_);
  not (_04854_, _00250_);
  nor (_04855_, _00596_, _04854_);
  not (_04856_, _04855_);
  nor (_04857_, _04856_, _04853_);
  not (_04858_, _04857_);
  nand (_04859_, _04858_, _04852_);
  nand (_04860_, _00382_, _00224_);
  nor (_04862_, _04860_, _00480_);
  not (_04863_, _04862_);
  not (_04864_, _00512_);
  nor (_04865_, _04864_, _30605_);
  not (_04866_, _04865_);
  nor (_04867_, _04866_, _30608_);
  not (_04869_, _04867_);
  nand (_04870_, _04869_, _04863_);
  nor (_04871_, _04870_, _04859_);
  nand (_04872_, _04871_, _04848_);
  nand (_04873_, _04872_, _04837_);
  not (_04875_, _04873_);
  nor (_04876_, _00624_, _00201_);
  not (_04878_, _04876_);
  nor (_04880_, _04842_, _00204_);
  nor (_04881_, _04846_, _00230_);
  nor (_04882_, _04881_, _04880_);
  not (_04883_, _04882_);
  nor (_04884_, _04860_, _00246_);
  nor (_04885_, _04884_, _04883_);
  nor (_04886_, _04885_, _04878_);
  nor (_04887_, _04850_, _00464_);
  nor (_04888_, _04856_, _00435_);
  nor (_04890_, _04866_, _00495_);
  nor (_04891_, _04890_, _04888_);
  not (_04892_, _04891_);
  nor (_04894_, _04892_, _04887_);
  nor (_04895_, _04894_, _04878_);
  nor (_04896_, _04895_, _04886_);
  nor (_04898_, _04896_, _04875_);
  not (_04899_, _04898_);
  nor (_04900_, _04899_, _04825_);
  nand (_04902_, _04875_, _04824_);
  nand (_04903_, _04902_, _04829_);
  nand (_04904_, _04903_, _29344_);
  nor (_09014_, _04904_, _04900_);
  nor (_04906_, _04296_, _03795_);
  nand (_04907_, _04906_, _26893_);
  nand (_04909_, _04907_, _00610_);
  nor (_04910_, _03818_, _27955_);
  not (_04911_, _04910_);
  nand (_04913_, _04911_, _04909_);
  nor (_04914_, _04907_, _30944_);
  nor (_04915_, _04914_, _04913_);
  nor (_04916_, _04911_, _27888_);
  nor (_04917_, _04916_, _04915_);
  nor (_09071_, _04917_, _23698_);
  nand (_04918_, _04906_, _00091_);
  nand (_04919_, _04918_, _00604_);
  nand (_04920_, _04919_, _04911_);
  nor (_04921_, _04918_, _30944_);
  nor (_04923_, _04921_, _04920_);
  nor (_04924_, _04911_, _28540_);
  nor (_04925_, _04924_, _04923_);
  nor (_09112_, _04925_, _23698_);
  nand (_04926_, _04906_, _30953_);
  nand (_04927_, _04926_, _00608_);
  nand (_04928_, _04927_, _04911_);
  nor (_04929_, _04926_, _30944_);
  nor (_04930_, _04929_, _04928_);
  nor (_04931_, _04911_, _27584_);
  nor (_04932_, _04931_, _04930_);
  nor (_09158_, _04932_, _23698_);
  nor (_04933_, _03795_, _00770_);
  nand (_04934_, _04933_, _26893_);
  nor (_04935_, _04934_, _30944_);
  nand (_04936_, _04934_, _00226_);
  nor (_04937_, _30885_, _04274_);
  nand (_04938_, _04937_, _03816_);
  nand (_04939_, _04938_, _04936_);
  nor (_04940_, _04939_, _04935_);
  nor (_04941_, _04938_, _27888_);
  nor (_04942_, _04941_, _04940_);
  nor (_09208_, _04942_, _23698_);
  nand (_04943_, _04933_, _27961_);
  nor (_04944_, _04943_, _30944_);
  nand (_04946_, _04943_, _04854_);
  nand (_04947_, _04946_, _04938_);
  nor (_04948_, _04947_, _04944_);
  nor (_04949_, _04938_, _28157_);
  nor (_04951_, _04949_, _04948_);
  nor (_09259_, _04951_, _23698_);
  nand (_04952_, _04933_, _00091_);
  nor (_04953_, _04952_, _30944_);
  nand (_04954_, _04952_, _30605_);
  nand (_04955_, _04954_, _04938_);
  nor (_04957_, _04955_, _04953_);
  nor (_04958_, _04938_, _28540_);
  nor (_04959_, _04958_, _04957_);
  nor (_09312_, _04959_, _23698_);
  nand (_04961_, _04933_, _00104_);
  nor (_04963_, _04961_, _30944_);
  nand (_04964_, _04961_, _00626_);
  nand (_04965_, _04964_, _04938_);
  nor (_04966_, _04965_, _04963_);
  nor (_04967_, _04938_, _27718_);
  nor (_04968_, _04967_, _04966_);
  nor (_09361_, _04968_, _23698_);
  nand (_04969_, _04933_, _30953_);
  nor (_04970_, _04969_, _30944_);
  nand (_04971_, _04969_, _30287_);
  nand (_04972_, _04971_, _04938_);
  nor (_04973_, _04972_, _04970_);
  nor (_04974_, _04938_, _27584_);
  nor (_04975_, _04974_, _04973_);
  nor (_09415_, _04975_, _23698_);
  nand (_04976_, _04933_, _31070_);
  nor (_04977_, _04976_, _30944_);
  nand (_04978_, _04976_, _04839_);
  nand (_04979_, _04978_, _04938_);
  nor (_04980_, _04979_, _04977_);
  nor (_04981_, _04938_, _28598_);
  nor (_04982_, _04981_, _04980_);
  nor (_09463_, _04982_, _23698_);
  nand (_04983_, _04933_, _31181_);
  nor (_04984_, _04983_, _30944_);
  nand (_04985_, _04983_, _00631_);
  nand (_04986_, _04985_, _04938_);
  nor (_04987_, _04986_, _04984_);
  nor (_04988_, _04938_, _28639_);
  nor (_04989_, _04988_, _04987_);
  nor (_09516_, _04989_, _23698_);
  nand (_04990_, _00771_, _26893_);
  nor (_04991_, _04990_, _30944_);
  nand (_04992_, _04990_, _00228_);
  nand (_04993_, _04992_, _00779_);
  nor (_04994_, _04993_, _04991_);
  nor (_04995_, _00788_, _27888_);
  nor (_04996_, _04995_, _04994_);
  nor (_09566_, _04996_, _23698_);
  nand (_04997_, _00771_, _00091_);
  nor (_04999_, _04997_, _30944_);
  nand (_05000_, _04997_, _30608_);
  nand (_05001_, _05000_, _00779_);
  nor (_05002_, _05001_, _04999_);
  nor (_05003_, _00788_, _28540_);
  nor (_05004_, _05003_, _05002_);
  nor (_09617_, _05004_, _23698_);
  nand (_05005_, _00771_, _27961_);
  nor (_05006_, _05005_, _30944_);
  nand (_05007_, _05005_, _04853_);
  nand (_05008_, _05007_, _00779_);
  nor (_05009_, _05008_, _05006_);
  nor (_05010_, _00788_, _28157_);
  nor (_05011_, _05010_, _05009_);
  nor (_09672_, _05011_, _23698_);
  nand (_05012_, _00771_, _00104_);
  nor (_05013_, _05012_, _30944_);
  nand (_05014_, _05012_, _00480_);
  nand (_05015_, _05014_, _00779_);
  nor (_05016_, _05015_, _05013_);
  nor (_05017_, _00788_, _27718_);
  nor (_05018_, _05017_, _05016_);
  nor (_09719_, _05018_, _23698_);
  nand (_05019_, _00771_, _30953_);
  nor (_05020_, _05019_, _30944_);
  nand (_05021_, _05019_, _30291_);
  nand (_05022_, _05021_, _00779_);
  nor (_05023_, _05022_, _05020_);
  nor (_05024_, _00788_, _27584_);
  nor (_05025_, _05024_, _05023_);
  nor (_09760_, _05025_, _23698_);
  nand (_05026_, _00771_, _31070_);
  nor (_05027_, _05026_, _30944_);
  nand (_05029_, _05026_, _04838_);
  nand (_05030_, _05029_, _00779_);
  nor (_05032_, _05030_, _05027_);
  nor (_05033_, _00788_, _28598_);
  nor (_05035_, _05033_, _05032_);
  nor (_09802_, _05035_, _23698_);
  nand (_05037_, _00771_, _31181_);
  nor (_05039_, _05037_, _30944_);
  nand (_05041_, _05037_, _00489_);
  nand (_05042_, _05041_, _00779_);
  nor (_05044_, _05042_, _05039_);
  nor (_05045_, _00788_, _28639_);
  nor (_05047_, _05045_, _05044_);
  nor (_09843_, _05047_, _23698_);
  not (_05049_, _04887_);
  not (_05050_, _04888_);
  nand (_05052_, _05050_, _05049_);
  not (_05053_, _04884_);
  not (_05055_, _04890_);
  nand (_05056_, _05055_, _05053_);
  nor (_05058_, _04883_, _02588_);
  nor (_05059_, _05058_, _05056_);
  nor (_05061_, _05059_, _05052_);
  nand (_05062_, _05061_, _04898_);
  not (_05064_, _04848_);
  nor (_05065_, _05064_, _02588_);
  nor (_05067_, _05065_, _04870_);
  nor (_05068_, _05067_, _04859_);
  nand (_05070_, _05068_, _04875_);
  nand (_05071_, _05070_, _05062_);
  nor (_05073_, _05071_, _04823_);
  nand (_05075_, _04823_, _02588_);
  nand (_05077_, _05075_, _29344_);
  nor (_09884_, _05077_, _05073_);
  nand (_05080_, _04894_, _05053_);
  nor (_05082_, _04883_, _00549_);
  nor (_05084_, _05082_, _05080_);
  nand (_05086_, _05084_, _04898_);
  nor (_05088_, _04848_, _04836_);
  nand (_05090_, _05088_, _04871_);
  nand (_05092_, _05090_, _05086_);
  nor (_05094_, _05092_, _04823_);
  not (_05096_, _00549_);
  nand (_05098_, _04823_, _05096_);
  nand (_05100_, _05098_, _29344_);
  nor (_09925_, _05100_, _05094_);
  nor (_05102_, _04823_, _00417_);
  not (_05105_, _05102_);
  nor (_05106_, _05105_, _04899_);
  nand (_05108_, _05102_, _04875_);
  nand (_05109_, _05108_, _04827_);
  nand (_05111_, _05109_, _29344_);
  nor (_09966_, _05111_, _05106_);
  not (_05113_, _04843_);
  nor (_05114_, _05113_, _04821_);
  nor (_05116_, _05114_, _00408_);
  not (_05117_, _04847_);
  nor (_05119_, _05117_, _04821_);
  nor (_05120_, _05119_, _04862_);
  not (_05122_, _05120_);
  nor (_05123_, _05122_, _05116_);
  nor (_05125_, _04867_, _04857_);
  not (_05126_, _00408_);
  nor (_05128_, _00417_, _05126_);
  nand (_05129_, _05128_, _04862_);
  nand (_05131_, _05129_, _05125_);
  nor (_05132_, _05131_, _05123_);
  not (_05134_, _05125_);
  nor (_05135_, _05134_, _04851_);
  nor (_05137_, _00417_, _00408_);
  nor (_05138_, _05137_, _04851_);
  nor (_05140_, _05138_, _05135_);
  nor (_05141_, _05140_, _05132_);
  nor (_05143_, _04873_, _04851_);
  nor (_05144_, _05128_, _04873_);
  nor (_05146_, _05144_, _05143_);
  nor (_05148_, _05146_, _05141_);
  not (_05150_, _04896_);
  nor (_05152_, _05150_, _04875_);
  nand (_05154_, _05152_, _05126_);
  not (_05156_, _04881_);
  nor (_05158_, _05156_, _04821_);
  nor (_05160_, _05158_, _04884_);
  not (_05162_, _04880_);
  nor (_05164_, _05162_, _04821_);
  nor (_05166_, _05164_, _00408_);
  nor (_05168_, _05166_, _04892_);
  nand (_05171_, _05168_, _05160_);
  not (_05173_, _05137_);
  nand (_05175_, _05173_, _04892_);
  nand (_05176_, _05175_, _05171_);
  nand (_05177_, _05176_, _05049_);
  not (_05178_, _05128_);
  nor (_05179_, _04892_, _05053_);
  nor (_05180_, _05179_, _04887_);
  nor (_05181_, _05180_, _05178_);
  nor (_05182_, _05181_, _04899_);
  nand (_05183_, _05182_, _05177_);
  nand (_05184_, _05183_, _05154_);
  nor (_05185_, _05184_, _05148_);
  nor (_05186_, _05185_, _04823_);
  nand (_05187_, _04823_, _05126_);
  nand (_05188_, _05187_, _29344_);
  nor (_10007_, _05188_, _05186_);
  nor (_10048_, _04822_, _02587_);
  not (_05189_, _00554_);
  nand (_05190_, _05162_, _05189_);
  nand (_05191_, _05190_, _05156_);
  nand (_05192_, _05191_, _05053_);
  nand (_05193_, _05192_, _05055_);
  nand (_05194_, _05193_, _05050_);
  nand (_05195_, _05194_, _04898_);
  nor (_05196_, _05195_, _04887_);
  nand (_05197_, _05113_, _05189_);
  nand (_05198_, _05197_, _05117_);
  nand (_05199_, _05198_, _04863_);
  nand (_05200_, _05199_, _04869_);
  nand (_05201_, _05200_, _04858_);
  nand (_05202_, _05201_, _05143_);
  nand (_05203_, _05202_, _04822_);
  nor (_05204_, _05203_, _05196_);
  nand (_05205_, _04823_, _05189_);
  nand (_05206_, _05205_, _29344_);
  nor (_10089_, _05206_, _05204_);
  nor (_05207_, _04875_, _04823_);
  nor (_05208_, _05207_, _04821_);
  nand (_05209_, _05152_, _05102_);
  nand (_05211_, _05209_, _29344_);
  nor (_10130_, _05211_, _05208_);
  not (_05212_, _00473_);
  nor (_05213_, _05212_, _04821_);
  not (_05214_, _05213_);
  nor (_05215_, _05214_, _04858_);
  nor (_05216_, _05113_, _00417_);
  nor (_05217_, _05216_, _05212_);
  nand (_05218_, _04847_, _04821_);
  nand (_05219_, _05218_, _04863_);
  nor (_05220_, _05219_, _05217_);
  nand (_05221_, _04858_, _04863_);
  nand (_05222_, _05221_, _05214_);
  nand (_05223_, _05222_, _04869_);
  nor (_05224_, _05223_, _05220_);
  nor (_05225_, _05224_, _05215_);
  nor (_05226_, _05225_, _04851_);
  nand (_05227_, _05212_, _00417_);
  nand (_05228_, _04867_, _04858_);
  nand (_05229_, _05228_, _04852_);
  nand (_05230_, _05229_, _05227_);
  nand (_05231_, _05230_, _04875_);
  nor (_05232_, _05231_, _05226_);
  nor (_05233_, _05214_, _05050_);
  nor (_05234_, _05162_, _00417_);
  nor (_05235_, _05234_, _05212_);
  nor (_05236_, _05156_, _00417_);
  nor (_05237_, _05236_, _04884_);
  not (_05238_, _05237_);
  nor (_05239_, _05238_, _05235_);
  nand (_05240_, _05050_, _05053_);
  nand (_05241_, _05240_, _05214_);
  nand (_05242_, _05241_, _05055_);
  nor (_05243_, _05242_, _05239_);
  nor (_05244_, _05243_, _05233_);
  nor (_05245_, _05244_, _04887_);
  nor (_05246_, _00473_, _04821_);
  nor (_05247_, _05055_, _04888_);
  nor (_05248_, _05247_, _04887_);
  nor (_05249_, _05248_, _05246_);
  nor (_05251_, _05249_, _04875_);
  nand (_05252_, _05251_, _05150_);
  nor (_05253_, _05252_, _05245_);
  nor (_05254_, _05253_, _05232_);
  nor (_05255_, _05254_, _04823_);
  nor (_05256_, _05152_, _04823_);
  not (_05257_, _05256_);
  nand (_05258_, _05257_, _05212_);
  nand (_05259_, _05258_, _29344_);
  nor (_10171_, _05259_, _05255_);
  nor (_05260_, _04822_, _02589_);
  nor (_05261_, _05260_, _05256_);
  nor (_10213_, _05261_, _23698_);
  nor (_10255_, _04822_, _02829_);
  not (_05262_, _00559_);
  nor (_05263_, _04822_, _05262_);
  nor (_05264_, _05263_, _05256_);
  nor (_10298_, _05264_, _23698_);
  nor (_05265_, _05216_, _00340_);
  nor (_05266_, _05265_, _05219_);
  not (_05267_, _00340_);
  nor (_05268_, _04821_, _05267_);
  not (_05269_, _05268_);
  nor (_05270_, _05269_, _04863_);
  nor (_05271_, _05270_, _05266_);
  nor (_05272_, _05271_, _05134_);
  nor (_05273_, _04821_, _00340_);
  nor (_05274_, _05273_, _05125_);
  nor (_05275_, _05274_, _05272_);
  nor (_05276_, _05275_, _04851_);
  nor (_05277_, _05268_, _04873_);
  nor (_05278_, _05277_, _05143_);
  nor (_05279_, _05278_, _05276_);
  nand (_05280_, _05152_, _05267_);
  not (_05281_, _05273_);
  nor (_05282_, _05281_, _04891_);
  nor (_05283_, _05282_, _04887_);
  not (_05284_, _05234_);
  nand (_05285_, _05284_, _05267_);
  nand (_05286_, _05285_, _05237_);
  nand (_05289_, _05286_, _04891_);
  nand (_05290_, _05289_, _05283_);
  nor (_05291_, _05269_, _05180_);
  nor (_05292_, _05291_, _04899_);
  nand (_05293_, _05292_, _05290_);
  nand (_05294_, _05293_, _05280_);
  nor (_05295_, _05294_, _05279_);
  nor (_05296_, _05295_, _04823_);
  nand (_05297_, _04823_, _05267_);
  nand (_05298_, _05297_, _29344_);
  nor (_10339_, _05298_, _05296_);
  not (_05299_, _00565_);
  nor (_05300_, _05299_, _00417_);
  not (_05301_, _05300_);
  nor (_05302_, _05301_, _04858_);
  nor (_05303_, _05114_, _05299_);
  nor (_05304_, _05303_, _05122_);
  nand (_05305_, _05301_, _05221_);
  nand (_05306_, _05305_, _04869_);
  nor (_05307_, _05306_, _05304_);
  nor (_05308_, _05307_, _05302_);
  nor (_05309_, _05308_, _04851_);
  nor (_05310_, _00565_, _00417_);
  not (_05311_, _05310_);
  nand (_05312_, _05311_, _05229_);
  nand (_05313_, _05312_, _04875_);
  nor (_05314_, _05313_, _05309_);
  nor (_05315_, _05301_, _05050_);
  not (_05316_, _05160_);
  nor (_05317_, _05164_, _05299_);
  nor (_05318_, _05317_, _05316_);
  nand (_05319_, _05301_, _05240_);
  nand (_05320_, _05319_, _05055_);
  nor (_05321_, _05320_, _05318_);
  nor (_05322_, _05321_, _05315_);
  nor (_05323_, _05322_, _04887_);
  nor (_05324_, _05310_, _05248_);
  nor (_05325_, _05324_, _04875_);
  nand (_05326_, _05325_, _05150_);
  nor (_05327_, _05326_, _05323_);
  nor (_05329_, _05327_, _05314_);
  nor (_05330_, _05329_, _04823_);
  nand (_05331_, _05257_, _05299_);
  nand (_05332_, _05331_, _29344_);
  nor (_10380_, _05332_, _05330_);
  nand (_05333_, _04933_, _31258_);
  nor (_05334_, _05333_, _30944_);
  nand (_05335_, _05333_, _00624_);
  nand (_05336_, _05335_, _04938_);
  nor (_05337_, _05336_, _05334_);
  nor (_05338_, _04938_, _28481_);
  nor (_05340_, _05338_, _05337_);
  nor (_10421_, _05340_, _23698_);
  nand (_05343_, _04906_, _31181_);
  nand (_05345_, _05343_, _00602_);
  nand (_05347_, _05345_, _04911_);
  nor (_05349_, _05343_, _30944_);
  nor (_05351_, _05349_, _05347_);
  nor (_05352_, _04911_, _28639_);
  nor (_05353_, _05352_, _05351_);
  nor (_10461_, _05353_, _23698_);
  nor (_05354_, _29297_, _27726_);
  nand (_05356_, _05354_, _31258_);
  nor (_05357_, _05356_, _27955_);
  not (_05358_, _05357_);
  nor (_05360_, _05358_, _30944_);
  not (_05361_, _00270_);
  nor (_05363_, _05300_, _05213_);
  nor (_05364_, _05363_, _04826_);
  nor (_05365_, _05364_, _05361_);
  nor (_05366_, _04821_, _00345_);
  not (_05368_, _05366_);
  nor (_05369_, _00417_, _00347_);
  nor (_05370_, _05369_, _04826_);
  nand (_05371_, _05370_, _05368_);
  nor (_05372_, _05268_, _05128_);
  not (_05373_, _05372_);
  nor (_05374_, _05373_, _05371_);
  nand (_05376_, _05374_, _05365_);
  nand (_05377_, _05376_, _00382_);
  nand (_05380_, _05377_, _04640_);
  nor (_05381_, _05380_, _05357_);
  nor (_05383_, _05381_, _05360_);
  nor (_05384_, _05383_, _04910_);
  nand (_05385_, _04910_, _28481_);
  nand (_05386_, _05385_, _29344_);
  nor (_10502_, _05386_, _05384_);
  not (_05387_, _10762_);
  nor (_05389_, _00277_, _05387_);
  not (_05391_, _05365_);
  nor (_05393_, _05372_, _04826_);
  nand (_05395_, _05393_, _05371_);
  nor (_05396_, _05395_, _05391_);
  nor (_05397_, _05396_, _00596_);
  nor (_05399_, _05397_, _05389_);
  nor (_05400_, _03957_, _27955_);
  nand (_05401_, _05400_, _29295_);
  nand (_05402_, _05401_, _05399_);
  nand (_05404_, _05402_, _04911_);
  nor (_05406_, _05401_, _30944_);
  nor (_05408_, _05406_, _05404_);
  nor (_05410_, _04911_, _28598_);
  nor (_05411_, _05410_, _05408_);
  nor (_10543_, _05411_, _23698_);
  nand (_05412_, _25952_, _00289_);
  nand (_05414_, _05364_, _00270_);
  not (_05416_, _05393_);
  nand (_05417_, _05416_, _05371_);
  nor (_05418_, _05417_, _05414_);
  nor (_05419_, _05418_, _00598_);
  nor (_05421_, _05419_, _05412_);
  nor (_05423_, _00795_, _27955_);
  nand (_05424_, _05423_, _29295_);
  nand (_05425_, _05424_, _05421_);
  nand (_05426_, _05425_, _04911_);
  nor (_05428_, _05424_, _30944_);
  nor (_05430_, _05428_, _05426_);
  nor (_05431_, _04911_, _28157_);
  nor (_05432_, _05431_, _05430_);
  nor (_10584_, _05432_, _23698_);
  not (_05435_, _03765_);
  nor (_05436_, _05435_, _27955_);
  nand (_05437_, _05436_, _29295_);
  nor (_05438_, _05437_, _30944_);
  nor (_05440_, _05414_, _05395_);
  nor (_05441_, _05440_, _04864_);
  nand (_05442_, _05441_, _00315_);
  nand (_05444_, _05437_, _05442_);
  nand (_05445_, _05444_, _04911_);
  nor (_05447_, _05445_, _05438_);
  nor (_05449_, _04911_, _27718_);
  nor (_05451_, _05449_, _05447_);
  nor (_10628_, _05451_, _23698_);
  not (_05454_, _00347_);
  nor (_05456_, _04822_, _05454_);
  nor (_05458_, _04862_, _05064_);
  nor (_05460_, _05135_, _04836_);
  nand (_05462_, _05460_, _05458_);
  nand (_05463_, _05462_, _00417_);
  nor (_05465_, _04886_, _04875_);
  nor (_05466_, _05465_, _05463_);
  nor (_05467_, _05466_, _00347_);
  nor (_05469_, _04894_, _04821_);
  nand (_05470_, _05469_, _04898_);
  not (_05471_, _05460_);
  nand (_05473_, _05471_, _04822_);
  nand (_05474_, _05473_, _05105_);
  nand (_05475_, _05474_, _05470_);
  nor (_05476_, _05475_, _05467_);
  nor (_05477_, _05476_, _05456_);
  nor (_10669_, _05477_, _23698_);
  not (_05479_, _00345_);
  nor (_05480_, _04822_, _05479_);
  nand (_05481_, _04895_, _04821_);
  nor (_05482_, _05481_, _04875_);
  nand (_05483_, _05473_, _04825_);
  nand (_05484_, _05483_, _05368_);
  nor (_05485_, _05484_, _05482_);
  nor (_05486_, _05485_, _05480_);
  not (_05487_, _05465_);
  nand (_05489_, _05487_, _05462_);
  nand (_05490_, _05489_, _05479_);
  nand (_05492_, _05490_, _29344_);
  nor (_10710_, _05492_, _05486_);
  nor (_10751_, _05387_, _23698_);
  nand (_05494_, _04896_, _04826_);
  nor (_05495_, _05494_, _04875_);
  nor (_05496_, _04821_, _00374_);
  nand (_05498_, _05496_, _04823_);
  nand (_05499_, _05498_, _29344_);
  nor (_10793_, _05499_, _05495_);
  nand (_05500_, _04896_, _00374_);
  nor (_05501_, _05500_, _04875_);
  not (_05502_, _05496_);
  nand (_05503_, _04821_, _00374_);
  nand (_05504_, _05503_, _05502_);
  nand (_05505_, _05504_, _04875_);
  nand (_05506_, _05505_, _04822_);
  nor (_05507_, _05506_, _05501_);
  nand (_05508_, _05504_, _04823_);
  nand (_05509_, _05508_, _29344_);
  nor (_10834_, _05509_, _05507_);
  nor (_10875_, _04822_, _02920_);
  nor (_10916_, _04638_, _23698_);
  nand (_05510_, _04276_, _27977_);
  nor (_05511_, _05510_, _00828_);
  not (_05512_, _30984_);
  nand (_05513_, _05510_, _05512_);
  nand (_05514_, _05513_, _29344_);
  nor (_10988_, _05514_, _05511_);
  nor (_05515_, _05510_, _00750_);
  not (_05516_, _00018_);
  nand (_05517_, _05510_, _05516_);
  nand (_05518_, _05517_, _29344_);
  nor (_11029_, _05518_, _05515_);
  nor (_05519_, _05510_, _00800_);
  nand (_05520_, _05510_, _30281_);
  nand (_05521_, _05520_, _29344_);
  nor (_11071_, _05521_, _05519_);
  nor (_05523_, _05510_, _27742_);
  not (_05524_, _00162_);
  nand (_05525_, _05510_, _05524_);
  nand (_05526_, _05525_, _29344_);
  nor (_11112_, _05526_, _05523_);
  nor (_05527_, _05510_, _00811_);
  not (_05528_, _30961_);
  nand (_05529_, _05510_, _05528_);
  nand (_05530_, _05529_, _29344_);
  nor (_11153_, _05530_, _05527_);
  nor (_05531_, _05510_, _28244_);
  not (_05532_, _00155_);
  nand (_05533_, _05510_, _05532_);
  nand (_05534_, _05533_, _29344_);
  nor (_11194_, _05534_, _05531_);
  nor (_05535_, _05510_, _27886_);
  nand (_05536_, _05510_, _00222_);
  nand (_05537_, _05536_, _29344_);
  nor (_11235_, _05537_, _05535_);
  nor (_05538_, _03950_, _27955_);
  not (_05539_, _05538_);
  nor (_05540_, _05539_, _28639_);
  nor (_05541_, _03686_, _27955_);
  nand (_05542_, _05541_, _31018_);
  not (_05543_, _31064_);
  not (_05544_, _31066_);
  nor (_05545_, _05544_, _05543_);
  not (_05546_, _31176_);
  not (_05547_, _31178_);
  not (_05548_, _31216_);
  nor (_05549_, _05548_, _00275_);
  not (_05550_, _05549_);
  nor (_05551_, _05550_, _05547_);
  not (_05552_, _05551_);
  nor (_05553_, _05552_, _05546_);
  nand (_05554_, _05553_, _05545_);
  not (_05555_, _12684_);
  nand (_05556_, _30971_, _05555_);
  nand (_05557_, _05556_, _30961_);
  nor (_05558_, _30964_, _30961_);
  nor (_05560_, _05558_, _00608_);
  nand (_05561_, _05560_, _05557_);
  not (_05562_, _31135_);
  not (_05563_, _31246_);
  not (_05564_, _31202_);
  nor (_05565_, _00268_, _05564_);
  nand (_05566_, _05565_, _31243_);
  nor (_05567_, _05566_, _05563_);
  not (_05568_, _05567_);
  nor (_05569_, _05568_, _05562_);
  not (_05570_, _05569_);
  nor (_05571_, _05570_, _05561_);
  not (_05572_, _05571_);
  nor (_05573_, _05572_, _05554_);
  nand (_05574_, _05573_, _31018_);
  nor (_05575_, _00158_, _00155_);
  not (_05576_, _05575_);
  nor (_05577_, _05573_, _31018_);
  nor (_05578_, _05577_, _05576_);
  nand (_05579_, _05578_, _05574_);
  nor (_05580_, _00222_, _00155_);
  not (_05581_, _31018_);
  not (_05582_, _31150_);
  not (_05583_, _31251_);
  not (_05584_, _31254_);
  nor (_05585_, _05584_, _05583_);
  nand (_05586_, _05585_, _05569_);
  nor (_05587_, _05586_, _05561_);
  not (_05588_, _05587_);
  nor (_05589_, _05588_, _05582_);
  not (_05590_, _05554_);
  nand (_05591_, _05590_, _05589_);
  nand (_05592_, _05591_, _05581_);
  nand (_05593_, _05592_, _05580_);
  not (_05594_, _05589_);
  nor (_05595_, _05554_, _05581_);
  not (_05596_, _05595_);
  nor (_05597_, _05596_, _05594_);
  nor (_05598_, _05597_, _05593_);
  nor (_05599_, _00602_, _03907_);
  nand (_05601_, _05599_, _05551_);
  nor (_05602_, _05601_, _05546_);
  nand (_05603_, _05602_, _31066_);
  nor (_05604_, _05603_, _05543_);
  nand (_05605_, _05604_, _00158_);
  nor (_05606_, _05605_, _05581_);
  nand (_05607_, _05605_, _05581_);
  nand (_05609_, _05607_, _00155_);
  nor (_05610_, _05609_, _05606_);
  nor (_05611_, _05610_, _05598_);
  nand (_05612_, _05611_, _05579_);
  nor (_05613_, _05541_, _05538_);
  nand (_05615_, _05613_, _05612_);
  nand (_05616_, _05615_, _05542_);
  nor (_05617_, _05616_, _05540_);
  nor (_11275_, _05617_, _23698_);
  nor (_05619_, _05539_, _00750_);
  not (_05620_, _05541_);
  nor (_05621_, _00158_, _05532_);
  nor (_05622_, _05621_, _05580_);
  not (_05624_, _05622_);
  not (_05625_, _05553_);
  nor (_05626_, _05625_, _05594_);
  nand (_05628_, _05626_, _31066_);
  nor (_05629_, _05628_, _00155_);
  nor (_05630_, _05629_, _31064_);
  not (_05632_, _05629_);
  nor (_05633_, _05632_, _05543_);
  nor (_05634_, _05633_, _05630_);
  nand (_05635_, _05634_, _05624_);
  nor (_05637_, _05572_, _05625_);
  nand (_05638_, _05637_, _31066_);
  nor (_05639_, _05638_, _05543_);
  nand (_05640_, _05638_, _05543_);
  nand (_05641_, _05640_, _05575_);
  nor (_05642_, _05641_, _05639_);
  nand (_05643_, _05603_, _05543_);
  nor (_05644_, _00222_, _05532_);
  not (_05645_, _05644_);
  nor (_05646_, _05645_, _05604_);
  nand (_05648_, _05646_, _05643_);
  nand (_05649_, _05648_, _05539_);
  nor (_05650_, _05649_, _05642_);
  nand (_05651_, _05650_, _05635_);
  nand (_05652_, _05651_, _05620_);
  nor (_05653_, _05652_, _05619_);
  nor (_05654_, _05620_, _05543_);
  nor (_05655_, _05654_, _05653_);
  nor (_11316_, _05655_, _23698_);
  nor (_05656_, _05620_, _05544_);
  nor (_05657_, _05539_, _00800_);
  nor (_05658_, _05626_, _31066_);
  nand (_05659_, _05628_, _05580_);
  nor (_05660_, _05659_, _05658_);
  nor (_05661_, _05637_, _31066_);
  nor (_05662_, _05661_, _05576_);
  nand (_05663_, _05662_, _05638_);
  nor (_05664_, _05602_, _31066_);
  nand (_05665_, _05644_, _05603_);
  nor (_05666_, _05665_, _05664_);
  not (_05667_, _05621_);
  nor (_05668_, _05667_, _05544_);
  nor (_05669_, _05668_, _05666_);
  nand (_05670_, _05669_, _05663_);
  nor (_05671_, _05670_, _05660_);
  nand (_05672_, _05671_, _05539_);
  nand (_05673_, _05672_, _05620_);
  nor (_05674_, _05673_, _05657_);
  nor (_05675_, _05674_, _05656_);
  nor (_11357_, _05675_, _23698_);
  nor (_05676_, _05539_, _27718_);
  nand (_05677_, _05541_, _31176_);
  nand (_05678_, _05601_, _05546_);
  nor (_05679_, _05645_, _05602_);
  nand (_05680_, _05679_, _05678_);
  nand (_05681_, _05551_, _05589_);
  nor (_05682_, _05681_, _00155_);
  nor (_05683_, _05682_, _31176_);
  not (_05684_, _05580_);
  nor (_05685_, _05626_, _05684_);
  nor (_05687_, _05685_, _05621_);
  nor (_05688_, _05687_, _05683_);
  nor (_05689_, _05572_, _05552_);
  nor (_05690_, _05689_, _31176_);
  not (_05691_, _05637_);
  nand (_05692_, _05691_, _05575_);
  nor (_05693_, _05692_, _05690_);
  nor (_05694_, _05693_, _05688_);
  nand (_05695_, _05694_, _05680_);
  nand (_05696_, _05695_, _05613_);
  nand (_05697_, _05696_, _05677_);
  nor (_05698_, _05697_, _05676_);
  nor (_11398_, _05698_, _23698_);
  nor (_05699_, _05620_, _05547_);
  nor (_05700_, _05539_, _00811_);
  nor (_05701_, _05572_, _05550_);
  nor (_05702_, _05701_, _31178_);
  nand (_05703_, _05701_, _31178_);
  nand (_05704_, _05703_, _05575_);
  nor (_05705_, _05704_, _05702_);
  nor (_05706_, _05550_, _05594_);
  nor (_05707_, _05706_, _31178_);
  nor (_05708_, _05707_, _05684_);
  nand (_05709_, _05708_, _05681_);
  not (_05710_, _05599_);
  nor (_05711_, _05710_, _05550_);
  nor (_05712_, _05711_, _31178_);
  nand (_05713_, _05644_, _05601_);
  nor (_05714_, _05713_, _05712_);
  nor (_05715_, _05667_, _05547_);
  nor (_05716_, _05715_, _05714_);
  nand (_05717_, _05716_, _05709_);
  nor (_05718_, _05717_, _05705_);
  nand (_05719_, _05718_, _05539_);
  nand (_05720_, _05719_, _05620_);
  nor (_05721_, _05720_, _05700_);
  nor (_05722_, _05721_, _05699_);
  nor (_11439_, _05722_, _23698_);
  nor (_05723_, _05539_, _28157_);
  nand (_05724_, _05541_, _31216_);
  nor (_05727_, _05710_, _00275_);
  not (_05728_, _05727_);
  nand (_05729_, _05728_, _05548_);
  nor (_05730_, _05645_, _05711_);
  nand (_05731_, _05730_, _05729_);
  nor (_05732_, _05594_, _00155_);
  nand (_05733_, _05732_, _31037_);
  not (_05734_, _05733_);
  nor (_05735_, _05734_, _31216_);
  nor (_05736_, _05706_, _05684_);
  nor (_05737_, _05736_, _05621_);
  nor (_05738_, _05737_, _05735_);
  nor (_05739_, _05561_, _00275_);
  nand (_05740_, _05739_, _05569_);
  nor (_05741_, _05740_, _05548_);
  nand (_05742_, _05740_, _05548_);
  nand (_05743_, _05742_, _05575_);
  nor (_05744_, _05743_, _05741_);
  nor (_05745_, _05744_, _05738_);
  nand (_05746_, _05745_, _05731_);
  nand (_05747_, _05746_, _05613_);
  nand (_05748_, _05747_, _05724_);
  nor (_05749_, _05748_, _05723_);
  nor (_11481_, _05749_, _23698_);
  nor (_05750_, _05539_, _27888_);
  nand (_05751_, _05541_, _31037_);
  nand (_05752_, _05572_, _31037_);
  nand (_05753_, _05571_, _00275_);
  nand (_05754_, _05753_, _05752_);
  nand (_05755_, _05754_, _05575_);
  nand (_05756_, _05710_, _00275_);
  nand (_05757_, _05756_, _05644_);
  nor (_05758_, _05757_, _05727_);
  nor (_05759_, _05732_, _31037_);
  nand (_05760_, _05733_, _05624_);
  nor (_05761_, _05760_, _05759_);
  nor (_05762_, _05761_, _05758_);
  nand (_05763_, _05762_, _05755_);
  nand (_05764_, _05763_, _05613_);
  nand (_05765_, _05764_, _05751_);
  nor (_05767_, _05765_, _05750_);
  nor (_11522_, _05767_, _23698_);
  nor (_05768_, _05572_, _05583_);
  nor (_05769_, _05768_, _31254_);
  nand (_05770_, _05576_, _05588_);
  nor (_05771_, _05770_, _05769_);
  nor (_05772_, _05667_, _05594_);
  not (_05773_, _05772_);
  nor (_05774_, _05773_, _05581_);
  nor (_05775_, _05774_, _05771_);
  nor (_05776_, _05775_, _05538_);
  nor (_05777_, _05575_, _05538_);
  nor (_05778_, _05777_, _05584_);
  nor (_05779_, _05778_, _05776_);
  nor (_05780_, _05779_, _05541_);
  nor (_05781_, _05620_, _28639_);
  nor (_05782_, _05781_, _05780_);
  nor (_11563_, _05782_, _23698_);
  nor (_05783_, _05620_, _00750_);
  not (_05784_, _05777_);
  nor (_05785_, _05784_, _05572_);
  nand (_05786_, _05785_, _31251_);
  not (_05787_, _05785_);
  nand (_05788_, _05787_, _05583_);
  nand (_05789_, _05788_, _05786_);
  nand (_05790_, _05772_, _31064_);
  nor (_05791_, _05790_, _05538_);
  nor (_05792_, _05791_, _05541_);
  nand (_05793_, _05792_, _05789_);
  nand (_05794_, _05793_, _29344_);
  nor (_11604_, _05794_, _05783_);
  nor (_05795_, _05620_, _00800_);
  not (_05796_, _31243_);
  nor (_05797_, _05561_, _00268_);
  not (_05798_, _05797_);
  nor (_05799_, _05798_, _05564_);
  not (_05800_, _05799_);
  nor (_05801_, _05800_, _05796_);
  not (_05802_, _05801_);
  nor (_05803_, _05802_, _05563_);
  nor (_05805_, _05803_, _31135_);
  nor (_05806_, _05805_, _05571_);
  not (_05807_, _05668_);
  nor (_05808_, _05807_, _05594_);
  nor (_05809_, _05808_, _05806_);
  nand (_05810_, _05809_, _05613_);
  nor (_05811_, _05539_, _31135_);
  nor (_05812_, _05811_, _23698_);
  nand (_05813_, _05812_, _05810_);
  nor (_11645_, _05813_, _05795_);
  nand (_05814_, _05538_, _31246_);
  not (_05815_, _05803_);
  nand (_05816_, _05802_, _05563_);
  nand (_05817_, _05816_, _05815_);
  nand (_05818_, _05772_, _31176_);
  nand (_05819_, _05818_, _05817_);
  nand (_05820_, _05819_, _05613_);
  nand (_05821_, _05820_, _05814_);
  nor (_05822_, _05620_, _27718_);
  nor (_05823_, _05822_, _05821_);
  nor (_11686_, _05823_, _23698_);
  nand (_05824_, _05538_, _31243_);
  nand (_05825_, _05800_, _05796_);
  nand (_05826_, _05825_, _05802_);
  nand (_05827_, _05715_, _05589_);
  nand (_05828_, _05827_, _05826_);
  nand (_05829_, _05828_, _05613_);
  nand (_05830_, _05829_, _05824_);
  nor (_05831_, _05620_, _28540_);
  nor (_05832_, _05831_, _05830_);
  nor (_11727_, _05832_, _23698_);
  nand (_05833_, _05538_, _31202_);
  nand (_05834_, _05798_, _05564_);
  nand (_05835_, _05834_, _05800_);
  nand (_05836_, _05772_, _31216_);
  nand (_05837_, _05836_, _05835_);
  nand (_05838_, _05837_, _05613_);
  nand (_05839_, _05838_, _05833_);
  nor (_05840_, _05620_, _28157_);
  nor (_05841_, _05840_, _05839_);
  nor (_11768_, _05841_, _23698_);
  nor (_05843_, _05539_, _00268_);
  nand (_05844_, _05541_, _27886_);
  nand (_05845_, _05561_, _00268_);
  nand (_05846_, _05845_, _05798_);
  nor (_05847_, _05594_, _00275_);
  nand (_05848_, _05621_, _05847_);
  nand (_05849_, _05848_, _05846_);
  nand (_05850_, _05849_, _05613_);
  nand (_05851_, _05850_, _05844_);
  nor (_05852_, _05851_, _05843_);
  nor (_11809_, _05852_, _23698_);
  not (_05853_, _31268_);
  nor (_05854_, _03673_, _27955_);
  not (_05855_, _05854_);
  nor (_05856_, _05855_, _05853_);
  nor (_05857_, _03959_, _27955_);
  not (_05858_, _05857_);
  nor (_05859_, _05858_, _00828_);
  not (_05860_, _31271_);
  not (_05861_, _12641_);
  nand (_05862_, _30990_, _05861_);
  nand (_05863_, _05862_, _30984_);
  nor (_05864_, _00602_, _30978_);
  not (_05865_, _05864_);
  nor (_05866_, _30984_, _30964_);
  nor (_05867_, _05866_, _05865_);
  nand (_05868_, _05867_, _05863_);
  not (_05869_, _31022_);
  not (_05870_, _31158_);
  not (_05871_, _31285_);
  nor (_05872_, _05871_, _05870_);
  not (_05873_, _05872_);
  nor (_05874_, _05873_, _05869_);
  not (_05875_, _31275_);
  nor (_05876_, _00265_, _05875_);
  not (_05877_, _05876_);
  not (_05878_, _31232_);
  not (_05879_, _31208_);
  not (_05880_, _31210_);
  nor (_05882_, _05880_, _05879_);
  nand (_05883_, _05882_, _31144_);
  nor (_05884_, _05883_, _05878_);
  nand (_05885_, _05884_, _31031_);
  nor (_05886_, _05885_, _05877_);
  not (_05887_, _05886_);
  not (_05888_, _31029_);
  not (_05889_, _31082_);
  nor (_05890_, _05889_, _05888_);
  nand (_05891_, _05890_, _31290_);
  nor (_05892_, _05891_, _05887_);
  nand (_05893_, _05892_, _05874_);
  nor (_05894_, _05893_, _05868_);
  not (_05895_, _05894_);
  nor (_05896_, _05895_, _05860_);
  nor (_05898_, _05896_, _31268_);
  nor (_05899_, _30281_, _00018_);
  nor (_05901_, _05860_, _05853_);
  not (_05902_, _05901_);
  nor (_05903_, _05902_, _05895_);
  not (_05904_, _05903_);
  nand (_05905_, _05904_, _05899_);
  nor (_05906_, _05905_, _05898_);
  nand (_05907_, _05886_, _05874_);
  nor (_05908_, _05868_, _05860_);
  not (_05909_, _05908_);
  nor (_05910_, _05909_, _05907_);
  nor (_05911_, _05910_, _31268_);
  nor (_05912_, _05516_, _05853_);
  nor (_05913_, _00022_, _00018_);
  not (_05914_, _05913_);
  nand (_05916_, _05910_, _31268_);
  not (_05917_, _05916_);
  nor (_05919_, _05917_, _05914_);
  nor (_05920_, _05919_, _05912_);
  nor (_05922_, _05920_, _05911_);
  nor (_05923_, _05922_, _05906_);
  nand (_05925_, _05923_, _05858_);
  nand (_05926_, _05925_, _05855_);
  nor (_05928_, _05926_, _05859_);
  nor (_05930_, _05928_, _05856_);
  nor (_11850_, _05930_, _23698_);
  nor (_05932_, _05858_, _28598_);
  nand (_05933_, _05854_, _31271_);
  nor (_05934_, _05854_, _05857_);
  nand (_05936_, _05895_, _05860_);
  not (_05938_, _05899_);
  nor (_05939_, _05938_, _05896_);
  nand (_05940_, _05939_, _05936_);
  not (_05941_, _05868_);
  not (_05943_, _05885_);
  nor (_05944_, _05877_, _05873_);
  nand (_05945_, _05944_, _05943_);
  nor (_05947_, _05945_, _05869_);
  nand (_05948_, _05947_, _05941_);
  nand (_05950_, _05948_, _05860_);
  nand (_05951_, _00018_, _31271_);
  not (_05952_, _05910_);
  nand (_05953_, _05913_, _05952_);
  nand (_05955_, _05953_, _05951_);
  nand (_05956_, _05955_, _05950_);
  nand (_05958_, _05956_, _05940_);
  nand (_05960_, _05958_, _05934_);
  nand (_05961_, _05960_, _05933_);
  nor (_05962_, _05961_, _05932_);
  nor (_11892_, _05962_, _23698_);
  nor (_05965_, _05858_, _27584_);
  nand (_05966_, _05854_, _31022_);
  nor (_05968_, _05885_, _05868_);
  not (_05969_, _05891_);
  nor (_05970_, _05969_, _30281_);
  nor (_05971_, _05877_, _00018_);
  nand (_05972_, _05971_, _05872_);
  nor (_05973_, _05972_, _05970_);
  nand (_05974_, _05973_, _05968_);
  nor (_05975_, _05974_, _05869_);
  not (_05976_, _05974_);
  nor (_05977_, _05976_, _31022_);
  nor (_05978_, _05977_, _05975_);
  nand (_05979_, _05978_, _05934_);
  nand (_05981_, _05979_, _05966_);
  nor (_05982_, _05981_, _05965_);
  nor (_11933_, _05982_, _23698_);
  nor (_05983_, _05858_, _27718_);
  nand (_05984_, _05854_, _31158_);
  nor (_05985_, _00018_, _05871_);
  nand (_05986_, _05985_, _05941_);
  nor (_05987_, _05986_, _05970_);
  nand (_05988_, _05987_, _05886_);
  not (_05989_, _05988_);
  nor (_05990_, _05989_, _31158_);
  nor (_05991_, _05988_, _05870_);
  nor (_05992_, _05991_, _05990_);
  nand (_05993_, _05992_, _05934_);
  nand (_05994_, _05993_, _05984_);
  nor (_05995_, _05994_, _05983_);
  nor (_11974_, _05995_, _23698_);
  nor (_05996_, _05858_, _28540_);
  nand (_05997_, _05854_, _31285_);
  nor (_05998_, _05914_, _05887_);
  not (_05999_, _05892_);
  nor (_06000_, _05938_, _05999_);
  nor (_06001_, _06000_, _05998_);
  nor (_06002_, _06001_, _05868_);
  nor (_06003_, _06002_, _31285_);
  nor (_06004_, _06003_, _05989_);
  nand (_06005_, _06004_, _05934_);
  nand (_06006_, _06005_, _05997_);
  nor (_06007_, _06006_, _05996_);
  nor (_12015_, _06007_, _23698_);
  nor (_06008_, _05858_, _28157_);
  nand (_06009_, _05854_, _31275_);
  not (_06010_, _05968_);
  nor (_06011_, _06010_, _00265_);
  nor (_06012_, _05970_, _00018_);
  nand (_06013_, _06012_, _06011_);
  nor (_06014_, _06013_, _05875_);
  not (_06015_, _06013_);
  nor (_06016_, _06015_, _31275_);
  nor (_06017_, _06016_, _06014_);
  nand (_06019_, _06017_, _05934_);
  nand (_06020_, _06019_, _06009_);
  nor (_06021_, _06020_, _06008_);
  nor (_12055_, _06021_, _23698_);
  not (_06022_, _05934_);
  nand (_06023_, _06010_, _00265_);
  nor (_06024_, _06011_, _05914_);
  nand (_06025_, _06024_, _06023_);
  nor (_06026_, _05516_, _00265_);
  nand (_06027_, _06011_, _05969_);
  nor (_06029_, _06010_, _05891_);
  not (_06030_, _06029_);
  nand (_06031_, _06030_, _00265_);
  nand (_06032_, _06031_, _06027_);
  nor (_06033_, _06032_, _05938_);
  nor (_06034_, _06033_, _06026_);
  nand (_06035_, _06034_, _06025_);
  nor (_06036_, _06035_, _06022_);
  nand (_06037_, _05857_, _27888_);
  nor (_06038_, _05855_, _31277_);
  nor (_06039_, _06038_, _23698_);
  nand (_06041_, _06039_, _06037_);
  nor (_12096_, _06041_, _06036_);
  nor (_06044_, _05855_, _00828_);
  not (_06046_, _31290_);
  nor (_06048_, _06010_, _05888_);
  nor (_06050_, _00022_, _05516_);
  nor (_06052_, _06050_, _05899_);
  nor (_06053_, _06052_, _05857_);
  nand (_06054_, _06053_, _06048_);
  nand (_06055_, _06054_, _06046_);
  nand (_06056_, _06048_, _31290_);
  not (_06057_, _06056_);
  nand (_06058_, _06053_, _06057_);
  nand (_06060_, _06058_, _06055_);
  not (_06062_, _06050_);
  nor (_06064_, _06062_, _06030_);
  nand (_06066_, _06064_, _31268_);
  nand (_06068_, _06066_, _05855_);
  nand (_06069_, _06068_, _05858_);
  nand (_06071_, _06069_, _06060_);
  nand (_06073_, _06071_, _29344_);
  nor (_12137_, _06073_, _06044_);
  nor (_06074_, _05855_, _00750_);
  nand (_06075_, _06053_, _05968_);
  nand (_06076_, _06075_, _31029_);
  not (_06077_, _06064_);
  nor (_06078_, _06077_, _05860_);
  nor (_06079_, _06078_, _05854_);
  nor (_06080_, _06079_, _05857_);
  nor (_06081_, _06075_, _31029_);
  nor (_06082_, _06081_, _06080_);
  nand (_06083_, _06082_, _06076_);
  nand (_06084_, _06083_, _29344_);
  nor (_12178_, _06084_, _06074_);
  not (_06085_, _05884_);
  nor (_06086_, _06085_, _05868_);
  nor (_06087_, _30281_, _05516_);
  nor (_06088_, _06087_, _05857_);
  nand (_06089_, _06088_, _06086_);
  nor (_06090_, _06089_, _31031_);
  nand (_06092_, _06050_, _31022_);
  nor (_06093_, _06092_, _05891_);
  nand (_06095_, _06093_, _05943_);
  nor (_06096_, _06095_, _05868_);
  nand (_06097_, _06096_, _05858_);
  nand (_06098_, _06089_, _31031_);
  nand (_06099_, _06098_, _06097_);
  nor (_06100_, _06099_, _06090_);
  nor (_06102_, _06100_, _05854_);
  nor (_06103_, _05855_, _27584_);
  nor (_06104_, _06103_, _06102_);
  nor (_12219_, _06104_, _23698_);
  nor (_06105_, _05855_, _27742_);
  nor (_06106_, _05883_, _05868_);
  nand (_06107_, _06088_, _06106_);
  nand (_06108_, _06107_, _05878_);
  nand (_06109_, _06108_, _06089_);
  nand (_06110_, _06064_, _31158_);
  nand (_06111_, _06110_, _05855_);
  nand (_06113_, _06111_, _05858_);
  nand (_06115_, _06113_, _06109_);
  nand (_06116_, _06115_, _29344_);
  nor (_12260_, _06116_, _06105_);
  nor (_06118_, _05855_, _00811_);
  not (_06120_, _06088_);
  not (_06121_, _05882_);
  nor (_06123_, _06121_, _05868_);
  nor (_06124_, _06123_, _31144_);
  nor (_06126_, _06124_, _06106_);
  nor (_06127_, _06126_, _06120_);
  nor (_06129_, _06088_, _31144_);
  nor (_06130_, _06129_, _06127_);
  nor (_06132_, _06056_, _05889_);
  not (_06134_, _06132_);
  nor (_06136_, _06062_, _06134_);
  nand (_06137_, _06136_, _31285_);
  nor (_06138_, _06137_, _05857_);
  nor (_06139_, _06138_, _06130_);
  nand (_06140_, _06139_, _05855_);
  nand (_06141_, _06140_, _29344_);
  nor (_12302_, _06141_, _06118_);
  nor (_06142_, _05855_, _28244_);
  nor (_06143_, _05868_, _05880_);
  nand (_06144_, _06088_, _06143_);
  nand (_06145_, _06144_, _31208_);
  nor (_06146_, _06144_, _31208_);
  nor (_06147_, _06077_, _05875_);
  nand (_06148_, _06147_, _05858_);
  nand (_06149_, _06148_, _05855_);
  nor (_06150_, _06149_, _06146_);
  nand (_06151_, _06150_, _06145_);
  nand (_06152_, _06151_, _29344_);
  nor (_12343_, _06152_, _06142_);
  nor (_06153_, _06088_, _05880_);
  nor (_06154_, _05941_, _31210_);
  nor (_06155_, _06154_, _06143_);
  nor (_06156_, _06027_, _05516_);
  nor (_06157_, _06156_, _06155_);
  nor (_06158_, _06157_, _06087_);
  nor (_06162_, _06158_, _05854_);
  nor (_06163_, _06162_, _05857_);
  nor (_06164_, _06163_, _06153_);
  nand (_06166_, _05854_, _27888_);
  nand (_06168_, _06166_, _29344_);
  nor (_12384_, _06168_, _06164_);
  nor (_06171_, _05620_, _28482_);
  nor (_06173_, _05784_, _05588_);
  not (_06175_, _06173_);
  nand (_06177_, _06175_, _31150_);
  nor (_06178_, _06175_, _31150_);
  not (_06179_, _30999_);
  nor (_06180_, _05773_, _06179_);
  nor (_06181_, _06180_, _05541_);
  nor (_06182_, _06181_, _05538_);
  nor (_06183_, _06182_, _06178_);
  nand (_06184_, _06183_, _06177_);
  nand (_06185_, _06184_, _29344_);
  nor (_12425_, _06185_, _06171_);
  not (_06186_, _05613_);
  nor (_06187_, _05596_, _06179_);
  not (_06188_, _06187_);
  nand (_06189_, _06188_, _05532_);
  nor (_06190_, _05575_, _05594_);
  nand (_06191_, _06190_, _06189_);
  not (_06192_, _05561_);
  nor (_06193_, _06192_, _05387_);
  not (_06194_, _05574_);
  nand (_06195_, _06194_, _30999_);
  nor (_06196_, _06195_, _05576_);
  nor (_06197_, _06196_, _06193_);
  nand (_06198_, _06197_, _06191_);
  nand (_06199_, _06198_, _29344_);
  nor (_12466_, _06199_, _06186_);
  nand (_06200_, _05868_, _30997_);
  not (_06201_, _05893_);
  not (_06202_, _31078_);
  nor (_06203_, _05902_, _06202_);
  nand (_06204_, _06203_, _05941_);
  not (_06205_, _06204_);
  nand (_06207_, _06205_, _06201_);
  nand (_06208_, _06207_, _06200_);
  nand (_06209_, _06208_, _05899_);
  not (_06210_, _06200_);
  nor (_06211_, _06204_, _05907_);
  nor (_06212_, _06211_, _06210_);
  nor (_06213_, _06212_, _05914_);
  nand (_06214_, _06087_, _30997_);
  nor (_06215_, _06200_, _06062_);
  nor (_06216_, _06215_, _06136_);
  nand (_06217_, _06216_, _06214_);
  nor (_06218_, _06217_, _06213_);
  nand (_06219_, _06218_, _06209_);
  nand (_06220_, _06219_, _29344_);
  nor (_12507_, _06220_, _06022_);
  nor (_06221_, _05858_, _28482_);
  nor (_06222_, _05916_, _05914_);
  nor (_06223_, _05904_, _05938_);
  nor (_06224_, _06223_, _06222_);
  not (_06225_, _06224_);
  nor (_06226_, _06225_, _06202_);
  nor (_06227_, _06224_, _31078_);
  nor (_06228_, _06227_, _06226_);
  nor (_06229_, _06228_, _05854_);
  nor (_06230_, _06229_, _05857_);
  nor (_06231_, _06230_, _06221_);
  nor (_06232_, _05855_, _06202_);
  nor (_06233_, _06232_, _06231_);
  nor (_12548_, _06233_, _23698_);
  not (_06234_, _06052_);
  nand (_06235_, _06056_, _05889_);
  nand (_06236_, _06235_, _06234_);
  nor (_06237_, _06236_, _06132_);
  nor (_06238_, _06077_, _06202_);
  nor (_06239_, _06238_, _06237_);
  nor (_06240_, _06239_, _06022_);
  nor (_06241_, _06053_, _05889_);
  nor (_06242_, _06241_, _05854_);
  nor (_06244_, _05855_, _28482_);
  nor (_06245_, _06244_, _06242_);
  nor (_06247_, _06245_, _06240_);
  nor (_12589_, _06247_, _23698_);
  nor (_12630_, _05861_, _23698_);
  nor (_12672_, _05555_, _23698_);
  nor (_06248_, _05510_, _28482_);
  not (_06249_, _30978_);
  nand (_06250_, _05510_, _06249_);
  nand (_06251_, _06250_, _29344_);
  nor (_12715_, _06251_, _06248_);
  nor (_06252_, _05539_, _28481_);
  nand (_06253_, _05541_, _30999_);
  nand (_06254_, _05599_, _05595_);
  nand (_06255_, _06254_, _06179_);
  nor (_06256_, _06254_, _06179_);
  nor (_06257_, _06256_, _05645_);
  nand (_06258_, _06257_, _06255_);
  not (_06259_, _05597_);
  nor (_06260_, _06259_, _00155_);
  nor (_06261_, _06260_, _30999_);
  nand (_06262_, _06187_, _05732_);
  nand (_06263_, _06262_, _05624_);
  nor (_06265_, _06263_, _06261_);
  nor (_06266_, _06194_, _30999_);
  nand (_06267_, _06195_, _05575_);
  nor (_06268_, _06267_, _06266_);
  nor (_06270_, _06268_, _06265_);
  nand (_06271_, _06270_, _06258_);
  nand (_06272_, _06271_, _05613_);
  nand (_06273_, _06272_, _06253_);
  nor (_06274_, _06273_, _06252_);
  nor (_12756_, _06274_, _23698_);
  nand (_06275_, _06188_, _05599_);
  nor (_06276_, _05599_, _30995_);
  nand (_06277_, _05644_, _29344_);
  nor (_06278_, _06277_, _06276_);
  nand (_06279_, _06278_, _06275_);
  nor (_12797_, _06279_, _06186_);
  not (_06280_, _01315_);
  nand (_06281_, _01290_, _17122_);
  nand (_06282_, _01296_, _17151_);
  nand (_06284_, _06282_, _06281_);
  nand (_06285_, _06284_, _01204_);
  nand (_06286_, _01296_, _17208_);
  nand (_06287_, _01290_, _17179_);
  nand (_06288_, _06287_, _06286_);
  nand (_06289_, _06288_, _01206_);
  nand (_06290_, _06289_, _06285_);
  nand (_06291_, _06290_, _01260_);
  nand (_06292_, _01290_, _17237_);
  nand (_06293_, _01296_, _17265_);
  nand (_06294_, _06293_, _06292_);
  nand (_06295_, _06294_, _01204_);
  nand (_06296_, _01296_, _17323_);
  nand (_06297_, _01290_, _17294_);
  nand (_06298_, _06297_, _06296_);
  nand (_06299_, _06298_, _01206_);
  nand (_06300_, _06299_, _06295_);
  nand (_06301_, _06300_, _01262_);
  nand (_06302_, _06301_, _06291_);
  nand (_06303_, _06302_, _01275_);
  nor (_06304_, _01296_, _17351_);
  nor (_06305_, _01290_, _17380_);
  nor (_06306_, _06305_, _06304_);
  nand (_06307_, _06306_, _01204_);
  nor (_06308_, _01290_, _17439_);
  nor (_06309_, _01296_, _17411_);
  nor (_06310_, _06309_, _06308_);
  nand (_06311_, _06310_, _01206_);
  nand (_06312_, _06311_, _06307_);
  nand (_06313_, _06312_, _01260_);
  nor (_06314_, _01296_, _17468_);
  nor (_06315_, _01290_, _17497_);
  nor (_06316_, _06315_, _06314_);
  nand (_06317_, _06316_, _01204_);
  nor (_06318_, _01290_, _17554_);
  nor (_06319_, _01296_, _17525_);
  nor (_06320_, _06319_, _06318_);
  nand (_06321_, _06320_, _01206_);
  nand (_06322_, _06321_, _06317_);
  nand (_06323_, _06322_, _01262_);
  nand (_06325_, _06323_, _06313_);
  nand (_06326_, _06325_, _01274_);
  nand (_06327_, _06326_, _06303_);
  nand (_06328_, _06327_, _01241_);
  nand (_06329_, _01296_, _16677_);
  nand (_06330_, _01290_, _16648_);
  nand (_06331_, _06330_, _06329_);
  nand (_06332_, _06331_, _01204_);
  nand (_06333_, _01290_, _16705_);
  nand (_06334_, _01296_, _16734_);
  nand (_06335_, _06334_, _06333_);
  nand (_06336_, _06335_, _01206_);
  nand (_06337_, _06336_, _06332_);
  nand (_06338_, _06337_, _01260_);
  nand (_06339_, _01296_, _16791_);
  nand (_06340_, _01290_, _16763_);
  nand (_06341_, _06340_, _06339_);
  nand (_06342_, _06341_, _01204_);
  nand (_06343_, _01290_, _16820_);
  nand (_06344_, _01296_, _16850_);
  nand (_06345_, _06344_, _06343_);
  nand (_06346_, _06345_, _01206_);
  nand (_06347_, _06346_, _06342_);
  nand (_06348_, _06347_, _01262_);
  nand (_06349_, _06348_, _06338_);
  nand (_06350_, _06349_, _01275_);
  nor (_06351_, _01296_, _16936_);
  nor (_06352_, _01290_, _16964_);
  nor (_06353_, _06352_, _06351_);
  nand (_06354_, _06353_, _01206_);
  nand (_06355_, _01290_, _16878_);
  nand (_06356_, _01296_, _16907_);
  nand (_06357_, _06356_, _06355_);
  nand (_06358_, _06357_, _01204_);
  nand (_06360_, _06358_, _06354_);
  nand (_06361_, _06360_, _01260_);
  nor (_06362_, _01296_, _17050_);
  nor (_06363_, _01290_, _17079_);
  nor (_06364_, _06363_, _06362_);
  nand (_06365_, _06364_, _01206_);
  nand (_06367_, _01290_, _16993_);
  nand (_06368_, _01296_, _17022_);
  nand (_06369_, _06368_, _06367_);
  nand (_06370_, _06369_, _01204_);
  nand (_06371_, _06370_, _06365_);
  nand (_06372_, _06371_, _01262_);
  nand (_06373_, _06372_, _06361_);
  nand (_06374_, _06373_, _01274_);
  nand (_06375_, _06374_, _06350_);
  nand (_06377_, _06375_, _01308_);
  nand (_06378_, _06377_, _06328_);
  nand (_06379_, _06378_, _01245_);
  nand (_06381_, _01296_, _15535_);
  nand (_06382_, _01290_, _15473_);
  nand (_06383_, _06382_, _06381_);
  nand (_06385_, _06383_, _01204_);
  nand (_06386_, _01290_, _15591_);
  nand (_06387_, _01296_, _15633_);
  nand (_06389_, _06387_, _06386_);
  nand (_06390_, _06389_, _01206_);
  nand (_06391_, _06390_, _06385_);
  nand (_06393_, _06391_, _01260_);
  nand (_06394_, _01296_, _15724_);
  nand (_06395_, _01290_, _15689_);
  nand (_06396_, _06395_, _06394_);
  nand (_06397_, _06396_, _01204_);
  nand (_06399_, _01290_, _15760_);
  nand (_06400_, _01296_, _15795_);
  nand (_06401_, _06400_, _06399_);
  nand (_06403_, _06401_, _01206_);
  nand (_06404_, _06403_, _06397_);
  nand (_06405_, _06404_, _01262_);
  nand (_06407_, _06405_, _06393_);
  nand (_06408_, _06407_, _01275_);
  nor (_06409_, _01296_, _15921_);
  nor (_06410_, _01290_, _15956_);
  nor (_06412_, _06410_, _06409_);
  nand (_06413_, _06412_, _01206_);
  nand (_06414_, _01290_, _15850_);
  nand (_06416_, _01296_, _15886_);
  nand (_06418_, _06416_, _06414_);
  nand (_06419_, _06418_, _01204_);
  nand (_06420_, _06419_, _06413_);
  nand (_06421_, _06420_, _01260_);
  nor (_06423_, _01296_, _16070_);
  nor (_06424_, _01290_, _16105_);
  nor (_06425_, _06424_, _06423_);
  nand (_06427_, _06425_, _01206_);
  nand (_06428_, _01290_, _15999_);
  nand (_06429_, _01296_, _16035_);
  nand (_06430_, _06429_, _06428_);
  nand (_06431_, _06430_, _01204_);
  nand (_06432_, _06431_, _06427_);
  nand (_06433_, _06432_, _01262_);
  nand (_06434_, _06433_, _06421_);
  nand (_06435_, _06434_, _01274_);
  nand (_06436_, _06435_, _06408_);
  nand (_06437_, _06436_, _01308_);
  nand (_06439_, _01290_, _16161_);
  nand (_06440_, _01296_, _16189_);
  nand (_06442_, _06440_, _06439_);
  nand (_06443_, _06442_, _01204_);
  nand (_06445_, _01296_, _16247_);
  nand (_06446_, _01290_, _16218_);
  nand (_06447_, _06446_, _06445_);
  nand (_06448_, _06447_, _01206_);
  nand (_06449_, _06448_, _06443_);
  nand (_06450_, _06449_, _01260_);
  nand (_06451_, _01290_, _16276_);
  nand (_06452_, _01296_, _16305_);
  nand (_06453_, _06452_, _06451_);
  nand (_06454_, _06453_, _01204_);
  nand (_06455_, _01296_, _16362_);
  nand (_06456_, _01290_, _16334_);
  nand (_06457_, _06456_, _06455_);
  nand (_06458_, _06457_, _01206_);
  nand (_06459_, _06458_, _06454_);
  nand (_06460_, _06459_, _01262_);
  nand (_06461_, _06460_, _06450_);
  nand (_06462_, _06461_, _01275_);
  nor (_06464_, _01296_, _16391_);
  nor (_06465_, _01290_, _16420_);
  nor (_06466_, _06465_, _06464_);
  nand (_06467_, _06466_, _01204_);
  nor (_06468_, _01290_, _16477_);
  nor (_06469_, _01296_, _16448_);
  nor (_06470_, _06469_, _06468_);
  nand (_06471_, _06470_, _01206_);
  nand (_06472_, _06471_, _06467_);
  nand (_06473_, _06472_, _01260_);
  nor (_06474_, _01296_, _16506_);
  nor (_06475_, _01290_, _16534_);
  nor (_06477_, _06475_, _06474_);
  nand (_06478_, _06477_, _01204_);
  nor (_06480_, _01290_, _16593_);
  nor (_06481_, _01296_, _16564_);
  nor (_06483_, _06481_, _06480_);
  nand (_06484_, _06483_, _01206_);
  nand (_06485_, _06484_, _06478_);
  nand (_06486_, _06485_, _01262_);
  nand (_06487_, _06486_, _06473_);
  nand (_06488_, _06487_, _01274_);
  nand (_06490_, _06488_, _06462_);
  nand (_06491_, _06490_, _01241_);
  nand (_06493_, _06491_, _06437_);
  nand (_06494_, _06493_, _01244_);
  nand (_06496_, _06494_, _06379_);
  nor (_06497_, _06496_, _01231_);
  nand (_06498_, _01296_, _18573_);
  nand (_06499_, _01290_, _18543_);
  nand (_06500_, _06499_, _06498_);
  nand (_06501_, _06500_, _01204_);
  nand (_06502_, _01290_, _18599_);
  nand (_06504_, _01296_, _18633_);
  nand (_06505_, _06504_, _06502_);
  nand (_06507_, _06505_, _01206_);
  nand (_06508_, _06507_, _06501_);
  nand (_06510_, _06508_, _01260_);
  nand (_06511_, _01296_, _18701_);
  nand (_06513_, _01290_, _18667_);
  nand (_06515_, _06513_, _06511_);
  nand (_06517_, _06515_, _01204_);
  nand (_06518_, _01290_, _18735_);
  nand (_06520_, _01296_, _18775_);
  nand (_06521_, _06520_, _06518_);
  nand (_06523_, _06521_, _01206_);
  nand (_06524_, _06523_, _06517_);
  nand (_06526_, _06524_, _01262_);
  nand (_06527_, _06526_, _06510_);
  nand (_06529_, _06527_, _01275_);
  nor (_06530_, _01296_, _18900_);
  nor (_06532_, _01290_, _18943_);
  nor (_06533_, _06532_, _06530_);
  nand (_06535_, _06533_, _01206_);
  nand (_06536_, _01290_, _18817_);
  nand (_06538_, _01296_, _18859_);
  nand (_06539_, _06538_, _06536_);
  nand (_06541_, _06539_, _01204_);
  nand (_06542_, _06541_, _06535_);
  nand (_06544_, _06542_, _01260_);
  nor (_06545_, _01296_, _19068_);
  nor (_06547_, _01290_, _19109_);
  nor (_06548_, _06547_, _06545_);
  nand (_06550_, _06548_, _01206_);
  nand (_06551_, _01290_, _18985_);
  nand (_06553_, _01296_, _19026_);
  nand (_06554_, _06553_, _06551_);
  nand (_06556_, _06554_, _01204_);
  nand (_06557_, _06556_, _06550_);
  nand (_06559_, _06557_, _01262_);
  nand (_06560_, _06559_, _06544_);
  nand (_06562_, _06560_, _01274_);
  nand (_06563_, _06562_, _06529_);
  nand (_06565_, _06563_, _01308_);
  nand (_06566_, _01290_, _19161_);
  nand (_06568_, _01296_, _19202_);
  nand (_06569_, _06568_, _06566_);
  nand (_06571_, _06569_, _01204_);
  nand (_06572_, _01296_, _19272_);
  nand (_06574_, _01290_, _19236_);
  nand (_06576_, _06574_, _06572_);
  nand (_06578_, _06576_, _01206_);
  nand (_06579_, _06578_, _06571_);
  nand (_06581_, _06579_, _01260_);
  nand (_06582_, _01290_, _19311_);
  nand (_06584_, _01296_, _19352_);
  nand (_06585_, _06584_, _06582_);
  nand (_06587_, _06585_, _01204_);
  nand (_06588_, _01296_, _19432_);
  nand (_06590_, _01290_, _19392_);
  nand (_06591_, _06590_, _06588_);
  nand (_06593_, _06591_, _01206_);
  nand (_06594_, _06593_, _06587_);
  nand (_06596_, _06594_, _01262_);
  nand (_06597_, _06596_, _06581_);
  nand (_06599_, _06597_, _01275_);
  nor (_06600_, _01296_, _19472_);
  nor (_06602_, _01290_, _19512_);
  nor (_06603_, _06602_, _06600_);
  nand (_06605_, _06603_, _01204_);
  nor (_06606_, _01290_, _19592_);
  nor (_06608_, _01296_, _19552_);
  nor (_06609_, _06608_, _06606_);
  nand (_06611_, _06609_, _01206_);
  nand (_06612_, _06611_, _06605_);
  nand (_06614_, _06612_, _01260_);
  nor (_06615_, _01296_, _19632_);
  nor (_06617_, _01290_, _19672_);
  nor (_06618_, _06617_, _06615_);
  nand (_06620_, _06618_, _01204_);
  nor (_06621_, _01290_, _19754_);
  nor (_06623_, _01296_, _19713_);
  nor (_06624_, _06623_, _06621_);
  nand (_06626_, _06624_, _01206_);
  nand (_06627_, _06626_, _06620_);
  nand (_06629_, _06627_, _01262_);
  nand (_06630_, _06629_, _06614_);
  nand (_06631_, _06630_, _01274_);
  nand (_06632_, _06631_, _06599_);
  nand (_06633_, _06632_, _01241_);
  nand (_06636_, _06633_, _06565_);
  nand (_06637_, _06636_, _01245_);
  nor (_06638_, _01296_, _18422_);
  nor (_06639_, _01290_, _18450_);
  nor (_06640_, _06639_, _06638_);
  nand (_06641_, _06640_, _01204_);
  nor (_06642_, _01290_, _18508_);
  nor (_06643_, _01296_, _18479_);
  nor (_06644_, _06643_, _06642_);
  nand (_06645_, _06644_, _01206_);
  nand (_06646_, _06645_, _06641_);
  nand (_06647_, _06646_, _01262_);
  nor (_06648_, _01296_, _18307_);
  nor (_06649_, _01290_, _18336_);
  nor (_06650_, _06649_, _06648_);
  nand (_06651_, _06650_, _01204_);
  nor (_06652_, _01290_, _18393_);
  nor (_06653_, _01296_, _18364_);
  nor (_06654_, _06653_, _06652_);
  nand (_06655_, _06654_, _01206_);
  nand (_06656_, _06655_, _06651_);
  nand (_06657_, _06656_, _01260_);
  nand (_06658_, _06657_, _06647_);
  nand (_06659_, _06658_, _01274_);
  nand (_06660_, _01290_, _18191_);
  nand (_06661_, _01296_, _18220_);
  nand (_06662_, _06661_, _06660_);
  nand (_06663_, _06662_, _01204_);
  nand (_06664_, _01296_, _18278_);
  nand (_06665_, _01290_, _18249_);
  nand (_06666_, _06665_, _06664_);
  nand (_06667_, _06666_, _01206_);
  nand (_06668_, _06667_, _06663_);
  nand (_06669_, _06668_, _01262_);
  nand (_06670_, _01290_, _18077_);
  nand (_06671_, _01296_, _18105_);
  nand (_06672_, _06671_, _06670_);
  nand (_06673_, _06672_, _01204_);
  nand (_06674_, _01296_, _18163_);
  nand (_06675_, _01290_, _18134_);
  nand (_06677_, _06675_, _06674_);
  nand (_06678_, _06677_, _01206_);
  nand (_06679_, _06678_, _06673_);
  nand (_06680_, _06679_, _01260_);
  nand (_06681_, _06680_, _06669_);
  nand (_06682_, _06681_, _01275_);
  nand (_06683_, _06682_, _06659_);
  nand (_06684_, _06683_, _01241_);
  nor (_06685_, _01296_, _18013_);
  nor (_06686_, _01290_, _18041_);
  nor (_06687_, _06686_, _06685_);
  nand (_06688_, _06687_, _01206_);
  nand (_06689_, _01290_, _17954_);
  nand (_06690_, _01296_, _17984_);
  nand (_06691_, _06690_, _06689_);
  nand (_06692_, _06691_, _01204_);
  nand (_06693_, _06692_, _06688_);
  nand (_06694_, _06693_, _01262_);
  nor (_06695_, _01296_, _17897_);
  nor (_06696_, _01290_, _17926_);
  nor (_06697_, _06696_, _06695_);
  nand (_06698_, _06697_, _01206_);
  nand (_06699_, _01290_, _17840_);
  nand (_06700_, _01296_, _17868_);
  nand (_06701_, _06700_, _06699_);
  nand (_06702_, _06701_, _01204_);
  nand (_06703_, _06702_, _06698_);
  nand (_06704_, _06703_, _01260_);
  nand (_06705_, _06704_, _06694_);
  nand (_06706_, _06705_, _01274_);
  nand (_06707_, _01296_, _17754_);
  nand (_06708_, _01290_, _17725_);
  nand (_06709_, _06708_, _06707_);
  nand (_06710_, _06709_, _01204_);
  nand (_06711_, _01290_, _17782_);
  nand (_06712_, _01296_, _17811_);
  nand (_06714_, _06712_, _06711_);
  nand (_06715_, _06714_, _01206_);
  nand (_06716_, _06715_, _06710_);
  nand (_06717_, _06716_, _01262_);
  nand (_06719_, _01296_, _17638_);
  nand (_06720_, _01290_, _17609_);
  nand (_06721_, _06720_, _06719_);
  nand (_06722_, _06721_, _01204_);
  nand (_06723_, _01290_, _17667_);
  nand (_06724_, _01296_, _17696_);
  nand (_06725_, _06724_, _06723_);
  nand (_06726_, _06725_, _01206_);
  nand (_06727_, _06726_, _06722_);
  nand (_06728_, _06727_, _01260_);
  nand (_06729_, _06728_, _06717_);
  nand (_06730_, _06729_, _01275_);
  nand (_06731_, _06730_, _06706_);
  nand (_06732_, _06731_, _01308_);
  nand (_06733_, _06732_, _06684_);
  nand (_06734_, _06733_, _01244_);
  nand (_06735_, _06734_, _06637_);
  nor (_06736_, _06735_, _01235_);
  nor (_06737_, _06736_, _06497_);
  nor (_06738_, _06737_, _28717_);
  nand (_06739_, _01290_, _21232_);
  nand (_06740_, _01296_, _21271_);
  nand (_06741_, _06740_, _06739_);
  nand (_06742_, _06741_, _01206_);
  nand (_06743_, _01296_, _21193_);
  nand (_06744_, _01290_, _21154_);
  nand (_06745_, _06744_, _06743_);
  nand (_06746_, _06745_, _01204_);
  nand (_06747_, _06746_, _06742_);
  nand (_06748_, _06747_, _01260_);
  nand (_06749_, _01290_, _21388_);
  nand (_06750_, _01296_, _21427_);
  nand (_06751_, _06750_, _06749_);
  nand (_06752_, _06751_, _01206_);
  nand (_06753_, _01296_, _21350_);
  nand (_06754_, _01290_, _21310_);
  nand (_06755_, _06754_, _06753_);
  nand (_06756_, _06755_, _01204_);
  nand (_06757_, _06756_, _06752_);
  nand (_06758_, _06757_, _01262_);
  nand (_06760_, _06758_, _06748_);
  nand (_06761_, _06760_, _01275_);
  nand (_06762_, _01290_, _21466_);
  nand (_06763_, _01296_, _21504_);
  nand (_06764_, _06763_, _06762_);
  nand (_06765_, _06764_, _01204_);
  nor (_06766_, _01296_, _21543_);
  nor (_06767_, _01290_, _21582_);
  nor (_06768_, _06767_, _06766_);
  nand (_06769_, _06768_, _01206_);
  nand (_06770_, _06769_, _06765_);
  nand (_06771_, _06770_, _01260_);
  nand (_06772_, _01290_, _21620_);
  nand (_06773_, _01296_, _21659_);
  nand (_06774_, _06773_, _06772_);
  nand (_06775_, _06774_, _01204_);
  nor (_06776_, _01296_, _21698_);
  nor (_06777_, _01290_, _21737_);
  nor (_06778_, _06777_, _06776_);
  nand (_06779_, _06778_, _01206_);
  nand (_06780_, _06779_, _06775_);
  nand (_06781_, _06780_, _01262_);
  nand (_06782_, _06781_, _06771_);
  nand (_06783_, _06782_, _01274_);
  nand (_06784_, _06783_, _06761_);
  nand (_06785_, _06784_, _01308_);
  nand (_06786_, _01290_, _21786_);
  nand (_06787_, _01296_, _21825_);
  nand (_06788_, _06787_, _06786_);
  nand (_06789_, _06788_, _01204_);
  nand (_06790_, _01296_, _21902_);
  nand (_06791_, _01290_, _21863_);
  nand (_06792_, _06791_, _06790_);
  nand (_06793_, _06792_, _01206_);
  nand (_06794_, _06793_, _06789_);
  nand (_06795_, _06794_, _01260_);
  nand (_06796_, _01290_, _21941_);
  nand (_06797_, _01296_, _21980_);
  nand (_06798_, _06797_, _06796_);
  nand (_06799_, _06798_, _01204_);
  nand (_06801_, _01296_, _22058_);
  nand (_06802_, _01290_, _22018_);
  nand (_06803_, _06802_, _06801_);
  nand (_06804_, _06803_, _01206_);
  nand (_06805_, _06804_, _06799_);
  nand (_06806_, _06805_, _01262_);
  nand (_06807_, _06806_, _06795_);
  nand (_06808_, _06807_, _01275_);
  nor (_06809_, _01296_, _22101_);
  nor (_06810_, _01290_, _22143_);
  nor (_06811_, _06810_, _06809_);
  nand (_06812_, _06811_, _01204_);
  nor (_06813_, _01290_, _22227_);
  nor (_06814_, _01296_, _22185_);
  nor (_06815_, _06814_, _06813_);
  nand (_06816_, _06815_, _01206_);
  nand (_06817_, _06816_, _06812_);
  nand (_06818_, _06817_, _01260_);
  nor (_06819_, _01296_, _22269_);
  nor (_06820_, _01290_, _22311_);
  nor (_06821_, _06820_, _06819_);
  nor (_06822_, _06821_, _01206_);
  nor (_06823_, _01290_, _22395_);
  nor (_06824_, _01296_, _22353_);
  nor (_06825_, _06824_, _06823_);
  nor (_06826_, _06825_, _01204_);
  nor (_06827_, _06826_, _06822_);
  nand (_06828_, _06827_, _01262_);
  nand (_06829_, _06828_, _06818_);
  nand (_06830_, _06829_, _01274_);
  nand (_06831_, _06830_, _06808_);
  nand (_06832_, _06831_, _01241_);
  nand (_06833_, _06832_, _06785_);
  nand (_06834_, _06833_, _01245_);
  nand (_06835_, _01290_, _19844_);
  nand (_06836_, _01296_, _19885_);
  nand (_06837_, _06836_, _06835_);
  nand (_06838_, _06837_, _01204_);
  nand (_06839_, _01296_, _19967_);
  nand (_06840_, _01290_, _19926_);
  nand (_06842_, _06840_, _06839_);
  nand (_06843_, _06842_, _01206_);
  nand (_06844_, _06843_, _06838_);
  nand (_06845_, _06844_, _01260_);
  nand (_06846_, _01290_, _20008_);
  nand (_06847_, _01296_, _20050_);
  nand (_06848_, _06847_, _06846_);
  nand (_06849_, _06848_, _01204_);
  nand (_06850_, _01296_, _20133_);
  nand (_06851_, _01290_, _20091_);
  nand (_06852_, _06851_, _06850_);
  nand (_06853_, _06852_, _01206_);
  nand (_06854_, _06853_, _06849_);
  nand (_06855_, _06854_, _01262_);
  nand (_06856_, _06855_, _06845_);
  nand (_06857_, _06856_, _01275_);
  nor (_06858_, _01296_, _20174_);
  nor (_06859_, _01290_, _20215_);
  nor (_06860_, _06859_, _06858_);
  nand (_06861_, _06860_, _01204_);
  nor (_06862_, _01290_, _20298_);
  nor (_06863_, _01296_, _20256_);
  nor (_06864_, _06863_, _06862_);
  nand (_06865_, _06864_, _01206_);
  nand (_06866_, _06865_, _06861_);
  nand (_06867_, _06866_, _01260_);
  nor (_06868_, _01296_, _20339_);
  nor (_06869_, _01290_, _20380_);
  nor (_06870_, _06869_, _06868_);
  nand (_06871_, _06870_, _01204_);
  nor (_06872_, _01290_, _20462_);
  nor (_06873_, _01296_, _20421_);
  nor (_06874_, _06873_, _06872_);
  nand (_06875_, _06874_, _01206_);
  nand (_06876_, _06875_, _06871_);
  nand (_06877_, _06876_, _01262_);
  nand (_06878_, _06877_, _06867_);
  nand (_06879_, _06878_, _01274_);
  nand (_06880_, _06879_, _06857_);
  nand (_06881_, _06880_, _01308_);
  nand (_06883_, _01290_, _20512_);
  nand (_06884_, _01296_, _20553_);
  nand (_06885_, _06884_, _06883_);
  nand (_06886_, _06885_, _01204_);
  nand (_06887_, _01296_, _20633_);
  nand (_06888_, _01290_, _20593_);
  nand (_06889_, _06888_, _06887_);
  nand (_06890_, _06889_, _01206_);
  nand (_06891_, _06890_, _06886_);
  nand (_06892_, _06891_, _01260_);
  nand (_06893_, _01290_, _20674_);
  nand (_06894_, _01296_, _20714_);
  nand (_06895_, _06894_, _06893_);
  nand (_06896_, _06895_, _01204_);
  nand (_06897_, _01296_, _20793_);
  nand (_06898_, _01290_, _20754_);
  nand (_06899_, _06898_, _06897_);
  nand (_06900_, _06899_, _01206_);
  nand (_06901_, _06900_, _06896_);
  nand (_06902_, _06901_, _01262_);
  nand (_06903_, _06902_, _06892_);
  nand (_06904_, _06903_, _01275_);
  nor (_06905_, _01296_, _20832_);
  nor (_06906_, _01290_, _20871_);
  nor (_06907_, _06906_, _06905_);
  nand (_06908_, _06907_, _01204_);
  nor (_06909_, _01290_, _20950_);
  nor (_06910_, _01296_, _20909_);
  nor (_06911_, _06910_, _06909_);
  nand (_06912_, _06911_, _01206_);
  nand (_06913_, _06912_, _06908_);
  nand (_06914_, _06913_, _01260_);
  nor (_06915_, _01296_, _20989_);
  nor (_06916_, _01290_, _21028_);
  nor (_06917_, _06916_, _06915_);
  nand (_06918_, _06917_, _01204_);
  nor (_06919_, _01290_, _21106_);
  nor (_06920_, _01296_, _21067_);
  nor (_06921_, _06920_, _06919_);
  nand (_06922_, _06921_, _01206_);
  nand (_06924_, _06922_, _06918_);
  nand (_06925_, _06924_, _01262_);
  nand (_06926_, _06925_, _06914_);
  nand (_06927_, _06926_, _01274_);
  nand (_06928_, _06927_, _06904_);
  nand (_06929_, _06928_, _01241_);
  nand (_06930_, _06929_, _06881_);
  nand (_06931_, _06930_, _01244_);
  nand (_06932_, _06931_, _06834_);
  nor (_06933_, _06932_, _01231_);
  nand (_06934_, _01296_, _23288_);
  nand (_06935_, _01290_, _23286_);
  nand (_06936_, _06935_, _06934_);
  nand (_06937_, _06936_, _01204_);
  nand (_06939_, _01290_, _23290_);
  nand (_06941_, _01296_, _23292_);
  nand (_06942_, _06941_, _06939_);
  nand (_06943_, _06942_, _01206_);
  nand (_06944_, _06943_, _06937_);
  nand (_06945_, _06944_, _01260_);
  nand (_06946_, _01296_, _23296_);
  nand (_06947_, _01290_, _23294_);
  nand (_06948_, _06947_, _06946_);
  nand (_06949_, _06948_, _01204_);
  nand (_06950_, _01290_, _23298_);
  nand (_06951_, _01296_, _23300_);
  nand (_06952_, _06951_, _06950_);
  nand (_06953_, _06952_, _01206_);
  nand (_06954_, _06953_, _06949_);
  nand (_06955_, _06954_, _01262_);
  nand (_06956_, _06955_, _06945_);
  nand (_06957_, _06956_, _01275_);
  nor (_06958_, _01296_, _23307_);
  nor (_06959_, _01290_, _23309_);
  nor (_06960_, _06959_, _06958_);
  nand (_06961_, _06960_, _01206_);
  nand (_06962_, _01290_, _23302_);
  nand (_06963_, _01296_, _23305_);
  nand (_06964_, _06963_, _06962_);
  nand (_06965_, _06964_, _01204_);
  nand (_06967_, _06965_, _06961_);
  nand (_06968_, _06967_, _01260_);
  nor (_06969_, _01296_, _23315_);
  nor (_06970_, _01290_, _23317_);
  nor (_06972_, _06970_, _06969_);
  nand (_06973_, _06972_, _01206_);
  nand (_06974_, _01290_, _23311_);
  nand (_06975_, _01296_, _23313_);
  nand (_06976_, _06975_, _06974_);
  nand (_06977_, _06976_, _01204_);
  nand (_06978_, _06977_, _06973_);
  nand (_06979_, _06978_, _01262_);
  nand (_06980_, _06979_, _06968_);
  nand (_06981_, _06980_, _01274_);
  nand (_06982_, _06981_, _06957_);
  nand (_06983_, _06982_, _01308_);
  nand (_06984_, _01290_, _23319_);
  nand (_06985_, _01296_, _23321_);
  nand (_06986_, _06985_, _06984_);
  nand (_06987_, _06986_, _01204_);
  nand (_06988_, _01296_, _23326_);
  nand (_06989_, _01290_, _23323_);
  nand (_06990_, _06989_, _06988_);
  nand (_06991_, _06990_, _01206_);
  nand (_06992_, _06991_, _06987_);
  nand (_06993_, _06992_, _01260_);
  nand (_06994_, _01290_, _23328_);
  nand (_06995_, _01296_, _23330_);
  nand (_06996_, _06995_, _06994_);
  nand (_06997_, _06996_, _01204_);
  nand (_06998_, _01296_, _23334_);
  nand (_06999_, _01290_, _23332_);
  nand (_07000_, _06999_, _06998_);
  nand (_07001_, _07000_, _01206_);
  nand (_07002_, _07001_, _06997_);
  nand (_07003_, _07002_, _01262_);
  nand (_07004_, _07003_, _06993_);
  nand (_07005_, _07004_, _01275_);
  nor (_07006_, _01296_, _23336_);
  nor (_07007_, _01290_, _23338_);
  nor (_07009_, _07007_, _07006_);
  nand (_07010_, _07009_, _01204_);
  nor (_07011_, _01290_, _23342_);
  nor (_07012_, _01296_, _23340_);
  nor (_07013_, _07012_, _07011_);
  nand (_07014_, _07013_, _01206_);
  nand (_07015_, _07014_, _07010_);
  nand (_07016_, _07015_, _01260_);
  nor (_07017_, _01296_, _23344_);
  nor (_07018_, _01290_, _23348_);
  nor (_07019_, _07018_, _07017_);
  nand (_07020_, _07019_, _01204_);
  nor (_07021_, _01290_, _23352_);
  nor (_07022_, _01296_, _23350_);
  nor (_07023_, _07022_, _07021_);
  nand (_07024_, _07023_, _01206_);
  nand (_07025_, _07024_, _07020_);
  nand (_07026_, _07025_, _01262_);
  nand (_07027_, _07026_, _07016_);
  nand (_07028_, _07027_, _01274_);
  nand (_07029_, _07028_, _07005_);
  nand (_07030_, _07029_, _01241_);
  nand (_07031_, _07030_, _06983_);
  nand (_07032_, _07031_, _01245_);
  nor (_07033_, _01296_, _23277_);
  nor (_07034_, _01290_, _23279_);
  nor (_07035_, _07034_, _07033_);
  nand (_07036_, _07035_, _01204_);
  nor (_07037_, _01290_, _23283_);
  nor (_07038_, _01296_, _23281_);
  nor (_07039_, _07038_, _07037_);
  nand (_07040_, _07039_, _01206_);
  nand (_07041_, _07040_, _07036_);
  nand (_07042_, _07041_, _01262_);
  nor (_07043_, _01296_, _23269_);
  nor (_07044_, _01290_, _23271_);
  nor (_07045_, _07044_, _07043_);
  nand (_07046_, _07045_, _01204_);
  nor (_07047_, _01290_, _23275_);
  nor (_07048_, _01296_, _23273_);
  nor (_07051_, _07048_, _07047_);
  nand (_07052_, _07051_, _01206_);
  nand (_07053_, _07052_, _07046_);
  nand (_07054_, _07053_, _01260_);
  nand (_07055_, _07054_, _07042_);
  nand (_07056_, _07055_, _01274_);
  nand (_07057_, _01290_, _23260_);
  nand (_07058_, _01296_, _23262_);
  nand (_07059_, _07058_, _07057_);
  nand (_07060_, _07059_, _01204_);
  nand (_07061_, _01296_, _23267_);
  nand (_07062_, _01290_, _23265_);
  nand (_07063_, _07062_, _07061_);
  nand (_07064_, _07063_, _01206_);
  nand (_07065_, _07064_, _07060_);
  nand (_07066_, _07065_, _01262_);
  nand (_07067_, _01290_, _23141_);
  nand (_07068_, _01296_, _23183_);
  nand (_07069_, _07068_, _07067_);
  nand (_07070_, _07069_, _01204_);
  nand (_07071_, _01296_, _23258_);
  nand (_07072_, _01290_, _23225_);
  nand (_07073_, _07072_, _07071_);
  nand (_07074_, _07073_, _01206_);
  nand (_07075_, _07074_, _07070_);
  nand (_07076_, _07075_, _01260_);
  nand (_07077_, _07076_, _07066_);
  nand (_07078_, _07077_, _01275_);
  nand (_07079_, _07078_, _07056_);
  nand (_07080_, _07079_, _01241_);
  nor (_07081_, _01296_, _23047_);
  nor (_07082_, _01290_, _23089_);
  nor (_07083_, _07082_, _07081_);
  nand (_07084_, _07083_, _01206_);
  nand (_07085_, _01290_, _22963_);
  nand (_07086_, _01296_, _23005_);
  nand (_07087_, _07086_, _07085_);
  nand (_07088_, _07087_, _01204_);
  nand (_07089_, _07088_, _07084_);
  nand (_07090_, _07089_, _01262_);
  nor (_07092_, _01296_, _22878_);
  nor (_07093_, _01290_, _22920_);
  nor (_07094_, _07093_, _07092_);
  nand (_07095_, _07094_, _01206_);
  nand (_07096_, _01290_, _22794_);
  nand (_07097_, _01296_, _22836_);
  nand (_07098_, _07097_, _07096_);
  nand (_07099_, _07098_, _01204_);
  nand (_07100_, _07099_, _07095_);
  nand (_07101_, _07100_, _01260_);
  nand (_07102_, _07101_, _07090_);
  nand (_07103_, _07102_, _01274_);
  nand (_07104_, _01296_, _22668_);
  nand (_07105_, _01290_, _22626_);
  nand (_07106_, _07105_, _07104_);
  nand (_07107_, _07106_, _01204_);
  nand (_07108_, _01290_, _22710_);
  nand (_07109_, _01296_, _22752_);
  nand (_07110_, _07109_, _07108_);
  nand (_07111_, _07110_, _01206_);
  nand (_07112_, _07111_, _07107_);
  nand (_07113_, _07112_, _01262_);
  nand (_07114_, _01296_, _22499_);
  nand (_07115_, _01290_, _22457_);
  nand (_07116_, _07115_, _07114_);
  nand (_07117_, _07116_, _01204_);
  nand (_07118_, _01290_, _22542_);
  nand (_07119_, _01296_, _22584_);
  nand (_07120_, _07119_, _07118_);
  nand (_07121_, _07120_, _01206_);
  nand (_07122_, _07121_, _07117_);
  nand (_07123_, _07122_, _01260_);
  nand (_07124_, _07123_, _07113_);
  nand (_07125_, _07124_, _01275_);
  nand (_07126_, _07125_, _07103_);
  nand (_07127_, _07126_, _01308_);
  nand (_07128_, _07127_, _07080_);
  nand (_07129_, _07128_, _01244_);
  nand (_07130_, _07129_, _07032_);
  nor (_07131_, _07130_, _01235_);
  nor (_07133_, _07131_, _06933_);
  nor (_07134_, _07133_, _28718_);
  nor (_07135_, _07134_, _06738_);
  nor (_07136_, _07135_, _06280_);
  not (_07137_, _04666_);
  nand (_07138_, _06280_, _07137_);
  nand (_07139_, _07138_, _29344_);
  nor (_12837_, _07139_, _07136_);
  nor (_12878_, _28788_, _23698_);
  nor (_12919_, _28900_, _23698_);
  nor (_12960_, _28775_, _23698_);
  nor (_13001_, _28913_, _23698_);
  nand (_13042_, _28978_, _29344_);
  nand (_13083_, _28185_, _29344_);
  nand (_13125_, _28009_, _29344_);
  nor (_13166_, _28768_, _23698_);
  not (_07140_, _28664_);
  nor (_13207_, _07140_, _23698_);
  nor (_07141_, _00146_, _29040_);
  nor (_07142_, _31257_, _27981_);
  nand (_07143_, _07142_, _27977_);
  nor (_07144_, _07143_, _00164_);
  not (_07145_, _30773_);
  nand (_07146_, _07143_, _07145_);
  nand (_07147_, _07146_, _29040_);
  nor (_07148_, _07147_, _07144_);
  nor (_07149_, _07148_, _07141_);
  nor (_13248_, _07149_, _23698_);
  nor (_07150_, _02221_, _29040_);
  nor (_07151_, _07143_, _02217_);
  nand (_07152_, _07143_, _30274_);
  nand (_07153_, _07152_, _29040_);
  nor (_07154_, _07153_, _07151_);
  nor (_07155_, _07154_, _07150_);
  nor (_13289_, _07155_, _23698_);
  nor (_07156_, _31124_, _29040_);
  nor (_07157_, _07143_, _31067_);
  not (_07158_, _30780_);
  nand (_07159_, _07143_, _07158_);
  nand (_07160_, _07159_, _29040_);
  nor (_07162_, _07160_, _07157_);
  nor (_07163_, _07162_, _07156_);
  nor (_13330_, _07163_, _23698_);
  not (_07164_, _31174_);
  nor (_07165_, _07164_, _29040_);
  nor (_07166_, _07143_, _31328_);
  not (_07167_, _30783_);
  nand (_07168_, _07143_, _07167_);
  nand (_07169_, _07168_, _29040_);
  nor (_07170_, _07169_, _07166_);
  nor (_07171_, _07170_, _07165_);
  nor (_13371_, _07171_, _23698_);
  nand (_07172_, _00091_, _26791_);
  nor (_07173_, _07172_, _27955_);
  nor (_07174_, _07173_, _29039_);
  nor (_07175_, _07174_, _31419_);
  nand (_07176_, _07174_, _00255_);
  nand (_07177_, _07176_, _29344_);
  nor (_13412_, _07177_, _07175_);
  nor (_07178_, _07174_, _30828_);
  not (_07179_, _30797_);
  nand (_07180_, _07174_, _07179_);
  nand (_07181_, _07180_, _29344_);
  nor (_13453_, _07181_, _07178_);
  nor (_07182_, _00088_, _29040_);
  nor (_07183_, _07143_, _30692_);
  nand (_07184_, _07143_, _30560_);
  nand (_07185_, _07184_, _29040_);
  nor (_07186_, _07185_, _07183_);
  nor (_07187_, _07186_, _07182_);
  nor (_13494_, _07187_, _23698_);
  nor (_07188_, _31396_, _29040_);
  nor (_07189_, _07143_, _30828_);
  not (_07190_, _30765_);
  nand (_07191_, _07143_, _07190_);
  nand (_07192_, _07191_, _29040_);
  nor (_07193_, _07192_, _07189_);
  nor (_07194_, _07193_, _07188_);
  nor (_13536_, _07194_, _23698_);
  nor (_07195_, _07174_, _30692_);
  nand (_07197_, _07174_, _30572_);
  nand (_07198_, _07197_, _29344_);
  nor (_13577_, _07198_, _07195_);
  nor (_07199_, _07174_, _00164_);
  not (_07200_, _30803_);
  nand (_07201_, _07174_, _07200_);
  nand (_07202_, _07201_, _29344_);
  nor (_13618_, _07202_, _07199_);
  nor (_07203_, _07174_, _02217_);
  nand (_07204_, _07174_, _30266_);
  nand (_07205_, _07204_, _29344_);
  nor (_13655_, _07205_, _07203_);
  nor (_07206_, _07174_, _31067_);
  not (_07207_, _30809_);
  nand (_07208_, _07174_, _07207_);
  nand (_07209_, _07208_, _29344_);
  nor (_13692_, _07209_, _07206_);
  nor (_07210_, _07174_, _31328_);
  not (_07211_, _30812_);
  nand (_07212_, _07174_, _07211_);
  nand (_07213_, _07212_, _29344_);
  nor (_13728_, _07213_, _07210_);
  nor (_07214_, _00042_, _29040_);
  nor (_07215_, _07143_, _31419_);
  not (_07216_, _30761_);
  nand (_07217_, _07143_, _07216_);
  nand (_07218_, _07217_, _29040_);
  nor (_07219_, _07218_, _07215_);
  nor (_07220_, _07219_, _07214_);
  nor (_13763_, _07220_, _23698_);
  nor (_07221_, _31320_, _29040_);
  nor (_07222_, _07143_, _31253_);
  not (_07223_, _30736_);
  nand (_07224_, _07143_, _07223_);
  nand (_07225_, _07224_, _29040_);
  nor (_07226_, _07225_, _07222_);
  nor (_07227_, _07226_, _07221_);
  nor (_13796_, _07227_, _23698_);
  nor (_07228_, _07174_, _31253_);
  not (_07229_, _30743_);
  nand (_07231_, _07174_, _07229_);
  nand (_07232_, _07231_, _29344_);
  nor (_13830_, _07232_, _07228_);
  not (_07233_, _02099_);
  nand (_07234_, _07233_, _27961_);
  nor (_07235_, _07234_, _30944_);
  nand (_07236_, _07234_, _00400_);
  nand (_07237_, _07236_, _27586_);
  nor (_07238_, _07237_, _07235_);
  nor (_07239_, _27586_, _28157_);
  nor (_07240_, _07239_, _07238_);
  nor (_13863_, _07240_, _23698_);
  nor (_07241_, _30685_, _30677_);
  not (_07242_, _30653_);
  nand (_07243_, _30844_, _30788_);
  nor (_07244_, _07243_, _07242_);
  nand (_07245_, _07244_, _03556_);
  nor (_07246_, _07245_, _30362_);
  nand (_07247_, _07246_, _30199_);
  nor (_07248_, _07247_, _31342_);
  nor (_07249_, _07248_, _30195_);
  nor (_07250_, _30898_, _30896_);
  not (_07251_, _30891_);
  nand (_07252_, _30896_, _07251_);
  nand (_07253_, _07252_, _27564_);
  nor (_07254_, _07253_, _07250_);
  nand (_07255_, _30903_, _28337_);
  nor (_07256_, _30903_, _28331_);
  nor (_07257_, _07256_, _30011_);
  nand (_07258_, _07257_, _07255_);
  not (_07259_, _30685_);
  nor (_07260_, _27040_, _28096_);
  nand (_07261_, _07260_, _28578_);
  nor (_07262_, _27645_, _28500_);
  not (_07263_, _29347_);
  nand (_07264_, _29345_, _27849_);
  nor (_07265_, _07264_, _07263_);
  nand (_07266_, _07265_, _07262_);
  nor (_07267_, _07266_, _07261_);
  nor (_07268_, _07267_, _07259_);
  nand (_07270_, _07268_, _07258_);
  nor (_07271_, _07270_, _07254_);
  nand (_07272_, _07271_, _29977_);
  nor (_07273_, _07272_, _07249_);
  nor (_07274_, _07273_, _07241_);
  nor (_07275_, _07274_, _07233_);
  nand (_07276_, _00092_, _30677_);
  nand (_07277_, _07276_, _07233_);
  nor (_07278_, _07277_, _04354_);
  nor (_07279_, _07278_, _07275_);
  nor (_07280_, _07279_, _26901_);
  nand (_07281_, _26901_, _28540_);
  nand (_07282_, _07281_, _29344_);
  nor (_13898_, _07282_, _07280_);
  nor (_07284_, _02099_, _00105_);
  nand (_07285_, _07284_, _30943_);
  not (_07286_, _07284_);
  nand (_07287_, _07286_, _27627_);
  nand (_07288_, _07287_, _07285_);
  nor (_07289_, _07288_, _26901_);
  nor (_07290_, _07289_, _27720_);
  nor (_13931_, _07290_, _23698_);
  nand (_07291_, _07233_, _30953_);
  nor (_07292_, _07291_, _30944_);
  nand (_07293_, _07291_, _26644_);
  nand (_07294_, _07293_, _27586_);
  nor (_07295_, _07294_, _07292_);
  nor (_07296_, _07295_, _27588_);
  nor (_13964_, _07296_, _23698_);
  nor (_07297_, _02099_, _31071_);
  not (_07298_, _07297_);
  nor (_07299_, _07298_, _30943_);
  nand (_07300_, _07298_, _30705_);
  nand (_07301_, _07300_, _27586_);
  nor (_07302_, _07301_, _07299_);
  nand (_07303_, _26901_, _28598_);
  nand (_07304_, _07303_, _29344_);
  nor (_13998_, _07304_, _07302_);
  nand (_07305_, _31182_, _30666_);
  nand (_07306_, _07305_, _07233_);
  nor (_07308_, _07306_, _03807_);
  not (_07309_, _30689_);
  nor (_07310_, _07309_, _07259_);
  nand (_07311_, _30364_, _27564_);
  nand (_07312_, _30010_, _30370_);
  nand (_07313_, _07312_, _07311_);
  nand (_07314_, _07313_, _07310_);
  nand (_07315_, _07310_, _30103_);
  nand (_07316_, _07315_, _30666_);
  nand (_07317_, _07316_, _07314_);
  nor (_07318_, _07317_, _07233_);
  nor (_07319_, _07318_, _07308_);
  nor (_07320_, _07319_, _26901_);
  nand (_07321_, _26901_, _28639_);
  nand (_07322_, _07321_, _29344_);
  nor (_14031_, _07322_, _07320_);
  nor (_07323_, _30943_, _29242_);
  nand (_07324_, _29242_, _30702_);
  nand (_07325_, _07324_, _02099_);
  nor (_07326_, _07325_, _07323_);
  nand (_07327_, _31259_, _30702_);
  nand (_07328_, _07327_, _04174_);
  nor (_07329_, _07328_, _02099_);
  nor (_07330_, _07329_, _07326_);
  nor (_07331_, _07330_, _26901_);
  nand (_07332_, _26901_, _28481_);
  nand (_07333_, _07332_, _29344_);
  nor (_14064_, _07333_, _07331_);
  nor (_07334_, _00785_, _26895_);
  nand (_07335_, _07334_, _30943_);
  nor (_07336_, _00775_, _00889_);
  nor (_07337_, _07336_, _30459_);
  nor (_07338_, _07337_, _29297_);
  nand (_07339_, _07338_, _07335_);
  nand (_07340_, _07336_, _27888_);
  nand (_07341_, _07340_, _26787_);
  nor (_07342_, _07341_, _07337_);
  nand (_07343_, _29294_, _30459_);
  nand (_07344_, _07343_, _29344_);
  nor (_07345_, _07344_, _07342_);
  nand (_14097_, _07345_, _07339_);
  nor (_07347_, _00785_, _31399_);
  nand (_07348_, _07347_, _30943_);
  nor (_07349_, _07347_, _30497_);
  nor (_07350_, _07349_, _29297_);
  nand (_07351_, _07350_, _07348_);
  nand (_07352_, _07336_, _28157_);
  nor (_07353_, _07336_, _30497_);
  nor (_07354_, _07353_, _26789_);
  nand (_07355_, _07354_, _07352_);
  nand (_07356_, _29294_, _30497_);
  nand (_07357_, _07356_, _07355_);
  nor (_07358_, _07357_, _23698_);
  nand (_14131_, _07358_, _07351_);
  nor (_07359_, _00785_, _00092_);
  nand (_07360_, _07359_, _30943_);
  nor (_07361_, _07359_, _30331_);
  nor (_07362_, _07361_, _29297_);
  nand (_07363_, _07362_, _07360_);
  nand (_07364_, _07336_, _28540_);
  nor (_07365_, _07336_, _30331_);
  nor (_07366_, _07365_, _26789_);
  nand (_07367_, _07366_, _07364_);
  nand (_07368_, _29294_, _30331_);
  nand (_07369_, _07368_, _07367_);
  nor (_07370_, _07369_, _23698_);
  nand (_14164_, _07370_, _07363_);
  nor (_07371_, _00785_, _00105_);
  nand (_07372_, _07371_, _30943_);
  nor (_07373_, _07371_, _30396_);
  nor (_07374_, _07373_, _29297_);
  nand (_07375_, _07374_, _07372_);
  nand (_07376_, _07336_, _27718_);
  nor (_07377_, _07336_, _30396_);
  nor (_07378_, _07377_, _26789_);
  nand (_07379_, _07378_, _07376_);
  nand (_07380_, _29294_, _30396_);
  nand (_07381_, _07380_, _07379_);
  nor (_07382_, _07381_, _23698_);
  nand (_14197_, _07382_, _07375_);
  nor (_07384_, _00889_, _27955_);
  nand (_07385_, _07384_, _30943_);
  nor (_07386_, _07384_, _30301_);
  nor (_07387_, _07386_, _29297_);
  nand (_07388_, _07387_, _07385_);
  nand (_07389_, _07384_, _27888_);
  nor (_07390_, _07386_, _26789_);
  nand (_07391_, _07390_, _07389_);
  nand (_07392_, _29294_, _30301_);
  nand (_07393_, _07392_, _07391_);
  nor (_07394_, _07393_, _23698_);
  nand (_14231_, _07394_, _07388_);
  not (_07395_, _30947_);
  nor (_07396_, _07395_, _04293_);
  not (_07397_, _07396_);
  nor (_07398_, _00092_, _07397_);
  nand (_07399_, _07398_, _30943_);
  nor (_07400_, _07398_, _30339_);
  nor (_07401_, _07400_, _29297_);
  nand (_07402_, _07401_, _07399_);
  nand (_07403_, _07384_, _28540_);
  nor (_07404_, _07384_, _30339_);
  nor (_07405_, _07404_, _26789_);
  nand (_07406_, _07405_, _07403_);
  nand (_07407_, _29294_, _30339_);
  nand (_07408_, _07407_, _07406_);
  nor (_07409_, _07408_, _23698_);
  nand (_14265_, _07409_, _07402_);
  nor (_07410_, _00105_, _07397_);
  nand (_07411_, _07410_, _30943_);
  nor (_07412_, _07410_, _30358_);
  nor (_07413_, _07412_, _29297_);
  nand (_07414_, _07413_, _07411_);
  nand (_07415_, _07384_, _27718_);
  nor (_07416_, _07384_, _30358_);
  nor (_07417_, _07416_, _26789_);
  nand (_07418_, _07417_, _07415_);
  nand (_07419_, _29294_, _30358_);
  nand (_07420_, _07419_, _07418_);
  nor (_07421_, _07420_, _23698_);
  nand (_14298_, _07421_, _07414_);
  nand (_07424_, _30943_, _27965_);
  nor (_07425_, _27965_, _30325_);
  nor (_07426_, _07425_, _29297_);
  nand (_07427_, _07426_, _07424_);
  nand (_07428_, _07384_, _28157_);
  nor (_07429_, _07384_, _30325_);
  nor (_07430_, _07429_, _26789_);
  nand (_07431_, _07430_, _07428_);
  nand (_07432_, _29294_, _30325_);
  nand (_07433_, _07432_, _07431_);
  nor (_07434_, _07433_, _23698_);
  nand (_14331_, _07434_, _07427_);
  nor (_07435_, _30954_, _07397_);
  nand (_07436_, _07435_, _30943_);
  nor (_07437_, _07435_, _30374_);
  nor (_07438_, _07437_, _29297_);
  nand (_07439_, _07438_, _07436_);
  nand (_07440_, _07384_, _27584_);
  nor (_07441_, _07384_, _30374_);
  nor (_07442_, _07441_, _26789_);
  nand (_07443_, _07442_, _07440_);
  nand (_07444_, _29294_, _30374_);
  nand (_07445_, _07444_, _07443_);
  nor (_07446_, _07445_, _23698_);
  nand (_14364_, _07446_, _07439_);
  nand (_07447_, _00769_, _30947_);
  nor (_07448_, _07447_, _00092_);
  nand (_07449_, _07448_, _30943_);
  nor (_07450_, _07448_, _30428_);
  nor (_07451_, _07450_, _29297_);
  nand (_07452_, _07451_, _07449_);
  nand (_07453_, _04937_, _30881_);
  not (_07454_, _07453_);
  nand (_07455_, _07454_, _28540_);
  nor (_07456_, _07454_, _30428_);
  nor (_07457_, _07456_, _26789_);
  nand (_07458_, _07457_, _07455_);
  nand (_07459_, _29294_, _30428_);
  nand (_07460_, _07459_, _07458_);
  nor (_07462_, _07460_, _23698_);
  nand (_14398_, _07462_, _07452_);
  nor (_07463_, _07447_, _31399_);
  nand (_07464_, _07463_, _30943_);
  nor (_07465_, _07463_, _30402_);
  nor (_07466_, _07465_, _29297_);
  nand (_07467_, _07466_, _07464_);
  nand (_07468_, _07454_, _28157_);
  nor (_07469_, _07454_, _30402_);
  nor (_07470_, _07469_, _26789_);
  nand (_07471_, _07470_, _07468_);
  nand (_07472_, _29294_, _30402_);
  nand (_07473_, _07472_, _07471_);
  nor (_07474_, _07473_, _23698_);
  nand (_14431_, _07474_, _07467_);
  nor (_07475_, _07447_, _26895_);
  nand (_07476_, _07475_, _30943_);
  nor (_07477_, _07454_, _30379_);
  nor (_07478_, _07477_, _29297_);
  nand (_07479_, _07478_, _07476_);
  nand (_07480_, _07454_, _27888_);
  nand (_07481_, _07480_, _26787_);
  nor (_07482_, _07481_, _07477_);
  nand (_07483_, _29294_, _30379_);
  nand (_07484_, _07483_, _29344_);
  nor (_07485_, _07484_, _07482_);
  nand (_14464_, _07485_, _07479_);
  nor (_07486_, _00785_, _30954_);
  nand (_07487_, _07486_, _30943_);
  nor (_07488_, _07486_, _30471_);
  nor (_07489_, _07488_, _29297_);
  nand (_07490_, _07489_, _07487_);
  nand (_07491_, _07336_, _27584_);
  nor (_07492_, _07336_, _30471_);
  nor (_07493_, _07492_, _26789_);
  nand (_07494_, _07493_, _07491_);
  nand (_07495_, _29294_, _30471_);
  nand (_07496_, _07495_, _07494_);
  nor (_07497_, _07496_, _23698_);
  nand (_14497_, _07497_, _07490_);
  nor (_07499_, _00785_, _31071_);
  nand (_07500_, _07499_, _30943_);
  nor (_07501_, _07499_, _30297_);
  nor (_07502_, _07501_, _29297_);
  nand (_07503_, _07502_, _07500_);
  nand (_07504_, _07336_, _28598_);
  nor (_07505_, _07336_, _30297_);
  nor (_07506_, _07505_, _26789_);
  nand (_07507_, _07506_, _07504_);
  nand (_07508_, _29294_, _30297_);
  nand (_07509_, _07508_, _07507_);
  nor (_07510_, _07509_, _23698_);
  nand (_14531_, _07510_, _07503_);
  nor (_07511_, _00785_, _31182_);
  nand (_07512_, _07511_, _30943_);
  nor (_07513_, _07511_, _30346_);
  nor (_07514_, _07513_, _29297_);
  nand (_07515_, _07514_, _07512_);
  nand (_07516_, _07336_, _28639_);
  nor (_07517_, _07336_, _30346_);
  nor (_07518_, _07517_, _26789_);
  nand (_07519_, _07518_, _07516_);
  nand (_07520_, _29294_, _30346_);
  nand (_07521_, _07520_, _07519_);
  nor (_07522_, _07521_, _23698_);
  nand (_14566_, _07522_, _07515_);
  nand (_07523_, _00783_, _04292_);
  nor (_07524_, _07523_, _31071_);
  nand (_07525_, _07524_, _30943_);
  nor (_07526_, _07524_, _30512_);
  nor (_07527_, _07526_, _29297_);
  nand (_07528_, _07527_, _07525_);
  nor (_07529_, _04304_, _00889_);
  nand (_07530_, _07529_, _28598_);
  nor (_07531_, _07529_, _30512_);
  nor (_07532_, _07531_, _26789_);
  nand (_07533_, _07532_, _07530_);
  nand (_07534_, _29294_, _30512_);
  nand (_07535_, _07534_, _07533_);
  nor (_07536_, _07535_, _23698_);
  nand (_14599_, _07536_, _07528_);
  nor (_07538_, _07523_, _31182_);
  nand (_07540_, _07538_, _30943_);
  nor (_07541_, _07538_, _30313_);
  nor (_07542_, _07541_, _29297_);
  nand (_07544_, _07542_, _07540_);
  nand (_07545_, _07529_, _28639_);
  nor (_07547_, _07529_, _30313_);
  nor (_07548_, _07547_, _26789_);
  nand (_07550_, _07548_, _07545_);
  nand (_07551_, _29294_, _30313_);
  nand (_07553_, _07551_, _07550_);
  nor (_07554_, _07553_, _23698_);
  nand (_14632_, _07554_, _07544_);
  nor (_07555_, _07523_, _00105_);
  nand (_07556_, _07555_, _30943_);
  nor (_07557_, _07555_, _30478_);
  nor (_07559_, _07557_, _29297_);
  nand (_07560_, _07559_, _07556_);
  nand (_07562_, _07529_, _27718_);
  nor (_07563_, _07529_, _30478_);
  nor (_07564_, _07563_, _26789_);
  nand (_07565_, _07564_, _07562_);
  nand (_07566_, _29294_, _30478_);
  nand (_07567_, _07566_, _07565_);
  nor (_07568_, _07567_, _23698_);
  nand (_14666_, _07568_, _07560_);
  nor (_07570_, _07523_, _30954_);
  nand (_07571_, _07570_, _30943_);
  nor (_07573_, _07570_, _30490_);
  nor (_07574_, _07573_, _29297_);
  nand (_07575_, _07574_, _07571_);
  nand (_07576_, _07529_, _27584_);
  nor (_07577_, _07529_, _30490_);
  nor (_07578_, _07577_, _26789_);
  nand (_07579_, _07578_, _07576_);
  nand (_07580_, _29294_, _30490_);
  nand (_07581_, _07580_, _07579_);
  nor (_07582_, _07581_, _23698_);
  nand (_14699_, _07582_, _07575_);
  nor (_07584_, _07523_, _00092_);
  nand (_07585_, _07584_, _30943_);
  nor (_07586_, _07584_, _30466_);
  nor (_07587_, _07586_, _29297_);
  nand (_07588_, _07587_, _07585_);
  nand (_07589_, _07529_, _28540_);
  nor (_07590_, _07529_, _30466_);
  nor (_07591_, _07590_, _26789_);
  nand (_07592_, _07591_, _07589_);
  nand (_07593_, _29294_, _30466_);
  nand (_07594_, _07593_, _07592_);
  nor (_07595_, _07594_, _23698_);
  nand (_14732_, _07595_, _07588_);
  nor (_07596_, _07523_, _26895_);
  nand (_07597_, _07596_, _30943_);
  nor (_07598_, _07529_, _30440_);
  nor (_07599_, _07598_, _29297_);
  nand (_07600_, _07599_, _07597_);
  nand (_07601_, _07529_, _27888_);
  nand (_07602_, _07601_, _26787_);
  nor (_07603_, _07602_, _07598_);
  nand (_07604_, _29294_, _30440_);
  nand (_07606_, _07604_, _29344_);
  nor (_07608_, _07606_, _07603_);
  nand (_14765_, _07608_, _07600_);
  nor (_07609_, _07523_, _31399_);
  nand (_07610_, _07609_, _30943_);
  nor (_07611_, _07609_, _30451_);
  nor (_07612_, _07611_, _29297_);
  nand (_07613_, _07612_, _07610_);
  nand (_07614_, _07529_, _28157_);
  nor (_07615_, _07529_, _30451_);
  nor (_07616_, _07615_, _26789_);
  nand (_07617_, _07616_, _07614_);
  nand (_07618_, _29294_, _30451_);
  nand (_07619_, _07618_, _07617_);
  nor (_07620_, _07619_, _23698_);
  nand (_14798_, _07620_, _07613_);
  nor (_07621_, _31182_, _07397_);
  nand (_07622_, _07621_, _30943_);
  nor (_07624_, _07621_, _30409_);
  nor (_07625_, _07624_, _29297_);
  nand (_07626_, _07625_, _07622_);
  nand (_07627_, _07384_, _28639_);
  nor (_07628_, _07384_, _30409_);
  nor (_07629_, _07628_, _26789_);
  nand (_07630_, _07629_, _07627_);
  nand (_07631_, _29294_, _30409_);
  nand (_07632_, _07631_, _07630_);
  nor (_07633_, _07632_, _23698_);
  nand (_14827_, _07633_, _07626_);
  nor (_07634_, _31071_, _07397_);
  nand (_07635_, _07634_, _30943_);
  nor (_07636_, _07634_, _30392_);
  nor (_07637_, _07636_, _29297_);
  nand (_07639_, _07637_, _07635_);
  nand (_07640_, _07384_, _28598_);
  nor (_07641_, _07384_, _30392_);
  nor (_07642_, _07641_, _26789_);
  nand (_07643_, _07642_, _07640_);
  nand (_07644_, _29294_, _30392_);
  nand (_07645_, _07644_, _07643_);
  nor (_07646_, _07645_, _23698_);
  nand (_14854_, _07646_, _07639_);
  nor (_07647_, _07523_, _31259_);
  nand (_07648_, _07647_, _30943_);
  nor (_07649_, _07647_, _30279_);
  nor (_07651_, _07649_, _29297_);
  nand (_07652_, _07651_, _07648_);
  nand (_07653_, _07529_, _28481_);
  nor (_07654_, _07529_, _30279_);
  nor (_07655_, _07654_, _26789_);
  nand (_07656_, _07655_, _07653_);
  nand (_07657_, _29294_, _30279_);
  nand (_07659_, _07657_, _07656_);
  nor (_07660_, _07659_, _23698_);
  nand (_14883_, _07660_, _07652_);
  nor (_07661_, _31259_, _07397_);
  nand (_07662_, _07661_, _30943_);
  nor (_07663_, _07661_, _30424_);
  nor (_07665_, _07663_, _29297_);
  nand (_07666_, _07665_, _07662_);
  nand (_07667_, _07384_, _28481_);
  nor (_07668_, _07384_, _30424_);
  nor (_07669_, _07668_, _26789_);
  nand (_07670_, _07669_, _07667_);
  nand (_07671_, _29294_, _30424_);
  nand (_07672_, _07671_, _07670_);
  nor (_07673_, _07672_, _23698_);
  nand (_14911_, _07673_, _07666_);
  nor (_07674_, _07447_, _00105_);
  nand (_07675_, _07674_, _30943_);
  nor (_07677_, _07674_, _30456_);
  nor (_07678_, _07677_, _29297_);
  nand (_07680_, _07678_, _07675_);
  nand (_07681_, _07454_, _27718_);
  nor (_07682_, _07454_, _30456_);
  nor (_07684_, _07682_, _26789_);
  nand (_07685_, _07684_, _07681_);
  nand (_07686_, _29294_, _30456_);
  nand (_07687_, _07686_, _07685_);
  nor (_07688_, _07687_, _23698_);
  nand (_14938_, _07688_, _07680_);
  nor (_07689_, _07447_, _30954_);
  nand (_07691_, _07689_, _30943_);
  nor (_07692_, _07689_, _30483_);
  nor (_07693_, _07692_, _29297_);
  nand (_07694_, _07693_, _07691_);
  nand (_07695_, _07454_, _27584_);
  nor (_07696_, _07454_, _30483_);
  nor (_07697_, _07696_, _26789_);
  nand (_07698_, _07697_, _07695_);
  nand (_07699_, _29294_, _30483_);
  nand (_07700_, _07699_, _07698_);
  nor (_07701_, _07700_, _23698_);
  nand (_14966_, _07701_, _07694_);
  nor (_07702_, _07447_, _31071_);
  nand (_07703_, _07702_, _30943_);
  nor (_07705_, _07702_, _30517_);
  nor (_07706_, _07705_, _29297_);
  nand (_07709_, _07706_, _07703_);
  nand (_07710_, _07454_, _28598_);
  nor (_07711_, _07454_, _30517_);
  nor (_07712_, _07711_, _26789_);
  nand (_07713_, _07712_, _07710_);
  nand (_07714_, _29294_, _30517_);
  nand (_07715_, _07714_, _07713_);
  nor (_07716_, _07715_, _23698_);
  nand (_14994_, _07716_, _07709_);
  nor (_07717_, _07447_, _31182_);
  nand (_07719_, _07717_, _30943_);
  nor (_07720_, _07717_, _30321_);
  nor (_07721_, _07720_, _29297_);
  nand (_07722_, _07721_, _07719_);
  nand (_07723_, _07454_, _28639_);
  nor (_07725_, _07454_, _30321_);
  nor (_07727_, _07725_, _26789_);
  nand (_07728_, _07727_, _07723_);
  nand (_07729_, _29294_, _30321_);
  nand (_07730_, _07729_, _07728_);
  nor (_07732_, _07730_, _23698_);
  nand (_15021_, _07732_, _07722_);
  nand (_07733_, _00786_, _30943_);
  nor (_07734_, _00786_, _30290_);
  nor (_07735_, _07734_, _29297_);
  nand (_07736_, _07735_, _07733_);
  nand (_07737_, _07336_, _28481_);
  nor (_07738_, _07336_, _30290_);
  nor (_07739_, _07738_, _26789_);
  nand (_07741_, _07739_, _07737_);
  nand (_07742_, _29294_, _30290_);
  nand (_07744_, _07742_, _07741_);
  nor (_07745_, _07744_, _23698_);
  nand (_15049_, _07745_, _07736_);
  nor (_07746_, _07447_, _31259_);
  nand (_07747_, _07746_, _30943_);
  nor (_07748_, _07746_, _30285_);
  nor (_07749_, _07748_, _29297_);
  nand (_07750_, _07749_, _07747_);
  nand (_07751_, _07454_, _28481_);
  nor (_07753_, _07454_, _30285_);
  nor (_07754_, _07753_, _26789_);
  nand (_07755_, _07754_, _07751_);
  nand (_07756_, _29294_, _30285_);
  nand (_07757_, _07756_, _07755_);
  nor (_07758_, _07757_, _23698_);
  nand (_15077_, _07758_, _07750_);
  nand (_07759_, _01290_, _27897_);
  nand (_07760_, _01296_, _23569_);
  nand (_07761_, _07760_, _07759_);
  nand (_07762_, _07761_, _01206_);
  nand (_07763_, _01296_, _23555_);
  nand (_07764_, _01290_, _27925_);
  nand (_07765_, _07764_, _07763_);
  nand (_07766_, _07765_, _01204_);
  nand (_07767_, _07766_, _07762_);
  nand (_07768_, _07767_, _01260_);
  nand (_07769_, _01290_, _27812_);
  nand (_07770_, _01296_, _27784_);
  nand (_07771_, _07770_, _07769_);
  nand (_07772_, _07771_, _01206_);
  nand (_07773_, _01296_, _27840_);
  nand (_07774_, _01290_, _27869_);
  nand (_07775_, _07774_, _07773_);
  nand (_07776_, _07775_, _01204_);
  nand (_07778_, _07776_, _07772_);
  nand (_07779_, _07778_, _01262_);
  nand (_07781_, _07779_, _07768_);
  nand (_07782_, _07781_, _01275_);
  nand (_07783_, _01290_, _27755_);
  nand (_07784_, _01296_, _27727_);
  nand (_07785_, _07784_, _07783_);
  nand (_07786_, _07785_, _01204_);
  nor (_07788_, _01296_, _27698_);
  nor (_07789_, _01290_, _27670_);
  nor (_07790_, _07789_, _07788_);
  nand (_07791_, _07790_, _01206_);
  nand (_07792_, _07791_, _07786_);
  nand (_07793_, _07792_, _01260_);
  nand (_07794_, _01290_, _23584_);
  nand (_07796_, _01296_, _27642_);
  nand (_07797_, _07796_, _07794_);
  nand (_07798_, _07797_, _01204_);
  nor (_07799_, _01296_, _27613_);
  nor (_07800_, _01290_, _27585_);
  nor (_07801_, _07800_, _07799_);
  nand (_07802_, _07801_, _01206_);
  nand (_07803_, _07802_, _07798_);
  nand (_07804_, _07803_, _01262_);
  nand (_07805_, _07804_, _07793_);
  nand (_07806_, _07805_, _01274_);
  nand (_07807_, _07806_, _07782_);
  nand (_07808_, _07807_, _01308_);
  nand (_07809_, _01290_, _27557_);
  nand (_07810_, _01296_, _27527_);
  nand (_07811_, _07810_, _07809_);
  nand (_07812_, _07811_, _01204_);
  nand (_07813_, _01296_, _23598_);
  nand (_07815_, _01290_, _27499_);
  nand (_07816_, _07815_, _07813_);
  nand (_07818_, _07816_, _01206_);
  nand (_07819_, _07818_, _07812_);
  nand (_07820_, _07819_, _01260_);
  nand (_07821_, _01290_, _23692_);
  nand (_07822_, _01296_, _23612_);
  nand (_07823_, _07822_, _07821_);
  nand (_07824_, _07823_, _01204_);
  nand (_07825_, _01296_, _27442_);
  nand (_07826_, _01290_, _27471_);
  nand (_07827_, _07826_, _07825_);
  nand (_07828_, _07827_, _01206_);
  nand (_07829_, _07828_, _07824_);
  nand (_07830_, _07829_, _01262_);
  nand (_07831_, _07830_, _07820_);
  nand (_07833_, _07831_, _01275_);
  nor (_07834_, _01296_, _27414_);
  nor (_07836_, _01290_, _27386_);
  nor (_07837_, _07836_, _07834_);
  nand (_07838_, _07837_, _01204_);
  nor (_07839_, _01290_, _27329_);
  nor (_07842_, _01296_, _27357_);
  nor (_07843_, _07842_, _07839_);
  nand (_07844_, _07843_, _01206_);
  nand (_07845_, _07844_, _07838_);
  nand (_07846_, _07845_, _01260_);
  nor (_07847_, _01296_, _27301_);
  nor (_07848_, _01290_, _27272_);
  nor (_07849_, _07848_, _07847_);
  nor (_07850_, _07849_, _01206_);
  nor (_07851_, _01290_, _27216_);
  nor (_07852_, _01296_, _27244_);
  nor (_07853_, _07852_, _07851_);
  nor (_07854_, _07853_, _01204_);
  nor (_07855_, _07854_, _07850_);
  nand (_07856_, _07855_, _01262_);
  nand (_07857_, _07856_, _07846_);
  nand (_07858_, _07857_, _01274_);
  nand (_07859_, _07858_, _07833_);
  nand (_07861_, _07859_, _01241_);
  nand (_07862_, _07861_, _07808_);
  nand (_07864_, _07862_, _01245_);
  nand (_07865_, _01290_, _28408_);
  nand (_07866_, _01296_, _28380_);
  nand (_07867_, _07866_, _07865_);
  nand (_07868_, _07867_, _01204_);
  nand (_07869_, _01296_, _28294_);
  nand (_07870_, _01290_, _28352_);
  nand (_07871_, _07870_, _07869_);
  nand (_07872_, _07871_, _01206_);
  nand (_07874_, _07872_, _07868_);
  nand (_07875_, _07874_, _01260_);
  nand (_07876_, _01290_, _28265_);
  nand (_07877_, _01296_, _28237_);
  nand (_07879_, _07877_, _07876_);
  nand (_07881_, _07879_, _01204_);
  nand (_07882_, _01296_, _28152_);
  nand (_07883_, _01290_, _28180_);
  nand (_07884_, _07883_, _07882_);
  nand (_07885_, _07884_, _01206_);
  nand (_07886_, _07885_, _07881_);
  nand (_07888_, _07886_, _01262_);
  nand (_07889_, _07888_, _07875_);
  nand (_07890_, _07889_, _01275_);
  nor (_07891_, _01296_, _28124_);
  nor (_07892_, _01290_, _28095_);
  nor (_07893_, _07892_, _07891_);
  nand (_07894_, _07893_, _01204_);
  nor (_07895_, _01290_, _23497_);
  nor (_07896_, _01296_, _28067_);
  nor (_07898_, _07896_, _07895_);
  nand (_07899_, _07898_, _01206_);
  nand (_07900_, _07899_, _07894_);
  nand (_07901_, _07900_, _01260_);
  nor (_07903_, _01296_, _23483_);
  nor (_07904_, _01290_, _23469_);
  nor (_07905_, _07904_, _07903_);
  nand (_07906_, _07905_, _01204_);
  nor (_07907_, _01290_, _23440_);
  nor (_07908_, _01296_, _23454_);
  nor (_07909_, _07908_, _07907_);
  nand (_07910_, _07909_, _01206_);
  nand (_07912_, _07910_, _07906_);
  nand (_07913_, _07912_, _01262_);
  nand (_07914_, _07913_, _07901_);
  nand (_07916_, _07914_, _01274_);
  nand (_07917_, _07916_, _07890_);
  nand (_07918_, _07917_, _01308_);
  nand (_07919_, _01290_, _23426_);
  nand (_07920_, _01296_, _23411_);
  nand (_07921_, _07920_, _07919_);
  nand (_07922_, _07921_, _01204_);
  nand (_07923_, _01296_, _23383_);
  nand (_07924_, _01290_, _23397_);
  nand (_07925_, _07924_, _07923_);
  nand (_07926_, _07925_, _01206_);
  nand (_07927_, _07926_, _07922_);
  nand (_07928_, _07927_, _01260_);
  nand (_07930_, _01290_, _23368_);
  nand (_07931_, _01296_, _23354_);
  nand (_07932_, _07931_, _07930_);
  nand (_07934_, _07932_, _01204_);
  nand (_07935_, _01296_, _28209_);
  nand (_07936_, _01290_, _29296_);
  nand (_07937_, _07936_, _07935_);
  nand (_07938_, _07937_, _01206_);
  nand (_07939_, _07938_, _07934_);
  nand (_07940_, _07939_, _01262_);
  nand (_07941_, _07940_, _07928_);
  nand (_07942_, _07941_, _01275_);
  nor (_07943_, _01296_, _28322_);
  nor (_07944_, _01290_, _23526_);
  nor (_07945_, _07944_, _07943_);
  nand (_07946_, _07945_, _01204_);
  nor (_07947_, _01290_, _28039_);
  nor (_07948_, _01296_, _23512_);
  nor (_07949_, _07948_, _07947_);
  nand (_07950_, _07949_, _01206_);
  nand (_07951_, _07950_, _07946_);
  nand (_07952_, _07951_, _01260_);
  nor (_07953_, _01296_, _28010_);
  nor (_07954_, _01290_, _27982_);
  nor (_07955_, _07954_, _07953_);
  nand (_07956_, _07955_, _01204_);
  nor (_07957_, _01290_, _23541_);
  nor (_07958_, _01296_, _27954_);
  nor (_07959_, _07958_, _07957_);
  nand (_07960_, _07959_, _01206_);
  nand (_07961_, _07960_, _07956_);
  nand (_07962_, _07961_, _01262_);
  nand (_07963_, _07962_, _07952_);
  nand (_07964_, _07963_, _01274_);
  nand (_07965_, _07964_, _07942_);
  nand (_07966_, _07965_, _01241_);
  nand (_07967_, _07966_, _07918_);
  nand (_07968_, _07967_, _01244_);
  nand (_07969_, _07968_, _07864_);
  nor (_07970_, _07969_, _01231_);
  nand (_07971_, _01296_, _26251_);
  nand (_07972_, _01290_, _26279_);
  nand (_07973_, _07972_, _07971_);
  nand (_07975_, _07973_, _01204_);
  nand (_07976_, _01290_, _26222_);
  nand (_07977_, _01296_, _26194_);
  nand (_07978_, _07977_, _07976_);
  nand (_07979_, _07978_, _01206_);
  nand (_07980_, _07979_, _07975_);
  nand (_07981_, _07980_, _01260_);
  nand (_07982_, _01296_, _26137_);
  nand (_07983_, _01290_, _26166_);
  nand (_07984_, _07983_, _07982_);
  nand (_07985_, _07984_, _01204_);
  nand (_07986_, _01290_, _26109_);
  nand (_07987_, _01296_, _26081_);
  nand (_07988_, _07987_, _07986_);
  nand (_07989_, _07988_, _01206_);
  nand (_07990_, _07989_, _07985_);
  nand (_07991_, _07990_, _01262_);
  nand (_07992_, _07991_, _07981_);
  nand (_07993_, _07992_, _01275_);
  nor (_07994_, _01296_, _25995_);
  nor (_07995_, _01290_, _25967_);
  nor (_07996_, _07995_, _07994_);
  nand (_07997_, _07996_, _01206_);
  nand (_07998_, _01290_, _26052_);
  nand (_07999_, _01296_, _26024_);
  nand (_08000_, _07999_, _07998_);
  nand (_08001_, _08000_, _01204_);
  nand (_08002_, _08001_, _07997_);
  nand (_08003_, _08002_, _01260_);
  nor (_08004_, _01296_, _25881_);
  nor (_08005_, _01290_, _25853_);
  nor (_08007_, _08005_, _08004_);
  nand (_08009_, _08007_, _01206_);
  nand (_08011_, _01290_, _25939_);
  nand (_08013_, _01296_, _25909_);
  nand (_08015_, _08013_, _08011_);
  nand (_08017_, _08015_, _01204_);
  nand (_08019_, _08017_, _08009_);
  nand (_08021_, _08019_, _01262_);
  nand (_08023_, _08021_, _08003_);
  nand (_08026_, _08023_, _01274_);
  nand (_08028_, _08026_, _07993_);
  nand (_08030_, _08028_, _01308_);
  nand (_08032_, _01290_, _25824_);
  nand (_08034_, _01296_, _25796_);
  nand (_08036_, _08034_, _08032_);
  nand (_08038_, _08036_, _01204_);
  nand (_08039_, _01296_, _25739_);
  nand (_08040_, _01290_, _25768_);
  nand (_08041_, _08040_, _08039_);
  nand (_08042_, _08041_, _01206_);
  nand (_08043_, _08042_, _08038_);
  nand (_08044_, _08043_, _01260_);
  nand (_08045_, _01290_, _25711_);
  nand (_08046_, _01296_, _25683_);
  nand (_08047_, _08046_, _08045_);
  nand (_08048_, _08047_, _01204_);
  nand (_08049_, _01296_, _25626_);
  nand (_08050_, _01290_, _25654_);
  nand (_08051_, _08050_, _08049_);
  nand (_08052_, _08051_, _01206_);
  nand (_08053_, _08052_, _08048_);
  nand (_08054_, _08053_, _01262_);
  nand (_08055_, _08054_, _08044_);
  nand (_08056_, _08055_, _01275_);
  nor (_08057_, _01296_, _25598_);
  nor (_08058_, _01290_, _25578_);
  nor (_08059_, _08058_, _08057_);
  nand (_08060_, _08059_, _01204_);
  nor (_08061_, _01290_, _25550_);
  nor (_08062_, _01296_, _25564_);
  nor (_08063_, _08062_, _08061_);
  nand (_08064_, _08063_, _01206_);
  nand (_08065_, _08064_, _08060_);
  nand (_08066_, _08065_, _01260_);
  nor (_08067_, _01296_, _25535_);
  nor (_08068_, _01290_, _25521_);
  nor (_08069_, _08068_, _08067_);
  nand (_08070_, _08069_, _01204_);
  nor (_08071_, _01290_, _25492_);
  nor (_08073_, _01296_, _25506_);
  nor (_08074_, _08073_, _08071_);
  nand (_08075_, _08074_, _01206_);
  nand (_08076_, _08075_, _08070_);
  nand (_08077_, _08076_, _01262_);
  nand (_08078_, _08077_, _08066_);
  nand (_08079_, _08078_, _01274_);
  nand (_08080_, _08079_, _08056_);
  nand (_08081_, _08080_, _01241_);
  nand (_08082_, _08081_, _08030_);
  nand (_08083_, _08082_, _01245_);
  nor (_08084_, _01296_, _26392_);
  nor (_08085_, _01290_, _26364_);
  nor (_08086_, _08085_, _08084_);
  nand (_08087_, _08086_, _01204_);
  nor (_08088_, _01290_, _26307_);
  nor (_08089_, _01296_, _26336_);
  nor (_08090_, _08089_, _08088_);
  nand (_08091_, _08090_, _01206_);
  nand (_08092_, _08091_, _08087_);
  nand (_08093_, _08092_, _01262_);
  nor (_08094_, _01296_, _26506_);
  nor (_08095_, _01290_, _26477_);
  nor (_08096_, _08095_, _08094_);
  nand (_08097_, _08096_, _01204_);
  nor (_08098_, _01290_, _26421_);
  nor (_08099_, _01296_, _26449_);
  nor (_08100_, _08099_, _08098_);
  nand (_08101_, _08100_, _01206_);
  nand (_08102_, _08101_, _08097_);
  nand (_08103_, _08102_, _01260_);
  nand (_08104_, _08103_, _08093_);
  nand (_08105_, _08104_, _01274_);
  nand (_08106_, _01290_, _26619_);
  nand (_08107_, _01296_, _26591_);
  nand (_08108_, _08107_, _08106_);
  nand (_08110_, _08108_, _01204_);
  nand (_08111_, _01296_, _26534_);
  nand (_08112_, _01290_, _26562_);
  nand (_08113_, _08112_, _08111_);
  nand (_08115_, _08113_, _01206_);
  nand (_08116_, _08115_, _08110_);
  nand (_08117_, _08116_, _01262_);
  nand (_08118_, _01290_, _26734_);
  nand (_08119_, _01296_, _26704_);
  nand (_08120_, _08119_, _08118_);
  nand (_08121_, _08120_, _01204_);
  nand (_08122_, _01296_, _26648_);
  nand (_08123_, _01290_, _26676_);
  nand (_08124_, _08123_, _08122_);
  nand (_08125_, _08124_, _01206_);
  nand (_08126_, _08125_, _08121_);
  nand (_08127_, _08126_, _01260_);
  nand (_08128_, _08127_, _08117_);
  nand (_08129_, _08128_, _01275_);
  nand (_08130_, _08129_, _08105_);
  nand (_08131_, _08130_, _01241_);
  nor (_08132_, _01296_, _26790_);
  nor (_08133_, _01290_, _26762_);
  nor (_08134_, _08133_, _08132_);
  nand (_08136_, _08134_, _01206_);
  nand (_08137_, _01290_, _26847_);
  nand (_08138_, _01296_, _26819_);
  nand (_08139_, _08138_, _08137_);
  nand (_08140_, _08139_, _01204_);
  nand (_08141_, _08140_, _08136_);
  nand (_08142_, _08141_, _01262_);
  nor (_08143_, _01296_, _26904_);
  nor (_08144_, _01290_, _26875_);
  nor (_08145_, _08144_, _08143_);
  nand (_08146_, _08145_, _01206_);
  nand (_08147_, _01290_, _26960_);
  nand (_08148_, _01296_, _26932_);
  nand (_08149_, _08148_, _08147_);
  nand (_08150_, _08149_, _01204_);
  nand (_08151_, _08150_, _08146_);
  nand (_08152_, _08151_, _01260_);
  nand (_08153_, _08152_, _08142_);
  nand (_08154_, _08153_, _01274_);
  nand (_08155_, _01296_, _27045_);
  nand (_08157_, _01290_, _27074_);
  nand (_08158_, _08157_, _08155_);
  nand (_08159_, _08158_, _01204_);
  nand (_08160_, _01290_, _27017_);
  nand (_08162_, _01296_, _26989_);
  nand (_08163_, _08162_, _08160_);
  nand (_08164_, _08163_, _01206_);
  nand (_08165_, _08164_, _08159_);
  nand (_08166_, _08165_, _01262_);
  nand (_08167_, _01296_, _27159_);
  nand (_08168_, _01290_, _27187_);
  nand (_08169_, _08168_, _08167_);
  nand (_08170_, _08169_, _01204_);
  nand (_08171_, _01290_, _27130_);
  nand (_08172_, _01296_, _27102_);
  nand (_08173_, _08172_, _08171_);
  nand (_08174_, _08173_, _01206_);
  nand (_08175_, _08174_, _08170_);
  nand (_08176_, _08175_, _01260_);
  nand (_08177_, _08176_, _08166_);
  nand (_08179_, _08177_, _01275_);
  nand (_08180_, _08179_, _08154_);
  nand (_08181_, _08180_, _01308_);
  nand (_08182_, _08181_, _08131_);
  nand (_08183_, _08182_, _01244_);
  nand (_08184_, _08183_, _08083_);
  nor (_08185_, _08184_, _01235_);
  nor (_08186_, _08185_, _07970_);
  nor (_08187_, _08186_, _28717_);
  nand (_08188_, _01290_, _24844_);
  nand (_08189_, _01296_, _24830_);
  nand (_08190_, _08189_, _08188_);
  nand (_08191_, _08190_, _01204_);
  nand (_08192_, _01296_, _24801_);
  nand (_08193_, _01290_, _24816_);
  nand (_08194_, _08193_, _08192_);
  nand (_08195_, _08194_, _01206_);
  nand (_08196_, _08195_, _08191_);
  nand (_08197_, _08196_, _01260_);
  nand (_08198_, _01290_, _24787_);
  nand (_08200_, _01296_, _24773_);
  nand (_08201_, _08200_, _08198_);
  nand (_08202_, _08201_, _01204_);
  nand (_08203_, _01296_, _24744_);
  nand (_08205_, _01290_, _24758_);
  nand (_08206_, _08205_, _08203_);
  nand (_08207_, _08206_, _01206_);
  nand (_08208_, _08207_, _08202_);
  nand (_08209_, _08208_, _01262_);
  nand (_08210_, _08209_, _08197_);
  nand (_08211_, _08210_, _01275_);
  nor (_08212_, _01296_, _24730_);
  nor (_08213_, _01290_, _24715_);
  nor (_08214_, _08213_, _08212_);
  nand (_08215_, _08214_, _01204_);
  nor (_08216_, _01290_, _24687_);
  nor (_08218_, _01296_, _24701_);
  nor (_08219_, _08218_, _08216_);
  nand (_08220_, _08219_, _01206_);
  nand (_08221_, _08220_, _08215_);
  nand (_08222_, _08221_, _01260_);
  nor (_08223_, _01296_, _24672_);
  nor (_08224_, _01290_, _24658_);
  nor (_08225_, _08224_, _08223_);
  nand (_08226_, _08225_, _01204_);
  nor (_08227_, _01290_, _24629_);
  nor (_08228_, _01296_, _24643_);
  nor (_08229_, _08228_, _08227_);
  nand (_08231_, _08229_, _01206_);
  nand (_08232_, _08231_, _08226_);
  nand (_08233_, _08232_, _01262_);
  nand (_08234_, _08233_, _08222_);
  nand (_08235_, _08234_, _01274_);
  nand (_08236_, _08235_, _08211_);
  nand (_08237_, _08236_, _01241_);
  nand (_08238_, _01296_, _25061_);
  nand (_08239_, _01290_, _25075_);
  nand (_08240_, _08239_, _08238_);
  nand (_08241_, _08240_, _01204_);
  nand (_08242_, _01290_, _25046_);
  nand (_08245_, _01296_, _25032_);
  nand (_08246_, _08245_, _08242_);
  nand (_08247_, _08246_, _01206_);
  nand (_08248_, _08247_, _08241_);
  nand (_08249_, _08248_, _01260_);
  nand (_08250_, _01296_, _25003_);
  nand (_08251_, _01290_, _25018_);
  nand (_08252_, _08251_, _08250_);
  nand (_08253_, _08252_, _01204_);
  nand (_08254_, _01290_, _24989_);
  nand (_08255_, _01296_, _24975_);
  nand (_08256_, _08255_, _08254_);
  nand (_08257_, _08256_, _01206_);
  nand (_08258_, _08257_, _08253_);
  nand (_08259_, _08258_, _01262_);
  nand (_08260_, _08259_, _08249_);
  nand (_08261_, _08260_, _01275_);
  nor (_08262_, _01296_, _24930_);
  nor (_08263_, _01290_, _24916_);
  nor (_08264_, _08263_, _08262_);
  nand (_08265_, _08264_, _01206_);
  nand (_08266_, _01290_, _24960_);
  nand (_08267_, _01296_, _24946_);
  nand (_08268_, _08267_, _08266_);
  nand (_08270_, _08268_, _01204_);
  nand (_08271_, _08270_, _08265_);
  nand (_08272_, _08271_, _01260_);
  nor (_08273_, _01296_, _24873_);
  nor (_08274_, _01290_, _24859_);
  nor (_08275_, _08274_, _08273_);
  nand (_08276_, _08275_, _01206_);
  nand (_08277_, _01290_, _24902_);
  nand (_08278_, _01296_, _24887_);
  nand (_08279_, _08278_, _08277_);
  nand (_08280_, _08279_, _01204_);
  nand (_08281_, _08280_, _08276_);
  nand (_08283_, _08281_, _01262_);
  nand (_08284_, _08283_, _08272_);
  nand (_08285_, _08284_, _01274_);
  nand (_08286_, _08285_, _08261_);
  nand (_08289_, _08286_, _01308_);
  nand (_08290_, _08289_, _08237_);
  nand (_08291_, _08290_, _01245_);
  nand (_08292_, _01296_, _25463_);
  nand (_08293_, _01290_, _25478_);
  nand (_08294_, _08293_, _08292_);
  nand (_08295_, _08294_, _01204_);
  nand (_08296_, _01290_, _25449_);
  nand (_08298_, _01296_, _25435_);
  nand (_08299_, _08298_, _08296_);
  nand (_08300_, _08299_, _01206_);
  nand (_08301_, _08300_, _08295_);
  nand (_08302_, _08301_, _01260_);
  nand (_08303_, _01296_, _25406_);
  nand (_08304_, _01290_, _25420_);
  nand (_08305_, _08304_, _08303_);
  nand (_08306_, _08305_, _01204_);
  nand (_08307_, _01290_, _25392_);
  nand (_08308_, _01296_, _25377_);
  nand (_08309_, _08308_, _08307_);
  nand (_08311_, _08309_, _01206_);
  nand (_08312_, _08311_, _08306_);
  nand (_08313_, _08312_, _01262_);
  nand (_08314_, _08313_, _08302_);
  nand (_08315_, _08314_, _01275_);
  nor (_08316_, _01296_, _25333_);
  nor (_08317_, _01290_, _25319_);
  nor (_08318_, _08317_, _08316_);
  nand (_08319_, _08318_, _01206_);
  nand (_08320_, _01290_, _25363_);
  nand (_08321_, _01296_, _25349_);
  nand (_08322_, _08321_, _08320_);
  nand (_08323_, _08322_, _01204_);
  nand (_08324_, _08323_, _08319_);
  nand (_08325_, _08324_, _01260_);
  nor (_08326_, _01296_, _25276_);
  nor (_08328_, _01290_, _25262_);
  nor (_08329_, _08328_, _08326_);
  nand (_08330_, _08329_, _01206_);
  nand (_08331_, _01290_, _25305_);
  nand (_08333_, _01296_, _25290_);
  nand (_08334_, _08333_, _08331_);
  nand (_08335_, _08334_, _01204_);
  nand (_08336_, _08335_, _08330_);
  nand (_08337_, _08336_, _01262_);
  nand (_08338_, _08337_, _08325_);
  nand (_08339_, _08338_, _01274_);
  nand (_08340_, _08339_, _08315_);
  nand (_08342_, _08340_, _01308_);
  nand (_08343_, _01290_, _25247_);
  nand (_08344_, _01296_, _25233_);
  nand (_08345_, _08344_, _08343_);
  nand (_08346_, _08345_, _01204_);
  nand (_08347_, _01296_, _25204_);
  nand (_08348_, _01290_, _25218_);
  nand (_08349_, _08348_, _08347_);
  nand (_08350_, _08349_, _01206_);
  nand (_08351_, _08350_, _08346_);
  nand (_08352_, _08351_, _01260_);
  nand (_08353_, _01290_, _25190_);
  nand (_08355_, _01296_, _25175_);
  nand (_08356_, _08355_, _08353_);
  nand (_08357_, _08356_, _01204_);
  nand (_08358_, _01296_, _25147_);
  nand (_08359_, _01290_, _25161_);
  nand (_08360_, _08359_, _08358_);
  nand (_08361_, _08360_, _01206_);
  nand (_08362_, _08361_, _08357_);
  nand (_08363_, _08362_, _01262_);
  nand (_08364_, _08363_, _08352_);
  nand (_08365_, _08364_, _01275_);
  nor (_08366_, _01296_, _25132_);
  nor (_08368_, _01290_, _25118_);
  nor (_08369_, _08368_, _08366_);
  nand (_08370_, _08369_, _01204_);
  nor (_08372_, _01290_, _23670_);
  nor (_08373_, _01296_, _25104_);
  nor (_08374_, _08373_, _08372_);
  nand (_08376_, _08374_, _01206_);
  nand (_08377_, _08376_, _08370_);
  nand (_08379_, _08377_, _01260_);
  nor (_08381_, _01296_, _23641_);
  nor (_08382_, _01290_, _23627_);
  nor (_08383_, _08382_, _08381_);
  nand (_08385_, _08383_, _01204_);
  nor (_08386_, _01290_, _25089_);
  nor (_08387_, _01296_, _23655_);
  nor (_08389_, _08387_, _08386_);
  nand (_08390_, _08389_, _01206_);
  nand (_08391_, _08390_, _08385_);
  nand (_08393_, _08391_, _01262_);
  nand (_08394_, _08393_, _08379_);
  nand (_08396_, _08394_, _01274_);
  nand (_08397_, _08396_, _08365_);
  nand (_08399_, _08397_, _01241_);
  nand (_08401_, _08399_, _08342_);
  nand (_08402_, _08401_, _01244_);
  nand (_08404_, _08402_, _08291_);
  nor (_08406_, _08404_, _01231_);
  nand (_08407_, _01296_, _24140_);
  nand (_08409_, _01290_, _24155_);
  nand (_08411_, _08409_, _08407_);
  nand (_08413_, _08411_, _01204_);
  nand (_08415_, _01290_, _24126_);
  nand (_08417_, _01296_, _24112_);
  nand (_08419_, _08417_, _08415_);
  nand (_08421_, _08419_, _01206_);
  nand (_08423_, _08421_, _08413_);
  nand (_08425_, _08423_, _01260_);
  nand (_08427_, _01296_, _24082_);
  nand (_08428_, _01290_, _24096_);
  nand (_08430_, _08428_, _08427_);
  nand (_08432_, _08430_, _01204_);
  nand (_08433_, _01290_, _24067_);
  nand (_08435_, _01296_, _24053_);
  nand (_08437_, _08435_, _08433_);
  nand (_08438_, _08437_, _01206_);
  nand (_08440_, _08438_, _08432_);
  nand (_08442_, _08440_, _01262_);
  nand (_08443_, _08442_, _08425_);
  nand (_08446_, _08443_, _01275_);
  nor (_08448_, _01296_, _24010_);
  nor (_08449_, _01290_, _23996_);
  nor (_08451_, _08449_, _08448_);
  nand (_08453_, _08451_, _01206_);
  nand (_08454_, _01290_, _24039_);
  nand (_08456_, _01296_, _24024_);
  nand (_08458_, _08456_, _08454_);
  nand (_08459_, _08458_, _01204_);
  nand (_08461_, _08459_, _08453_);
  nand (_08462_, _08461_, _01260_);
  nor (_08463_, _01296_, _23953_);
  nor (_08464_, _01290_, _23938_);
  nor (_08465_, _08464_, _08463_);
  nand (_08466_, _08465_, _01206_);
  nand (_08467_, _01290_, _23981_);
  nand (_08468_, _01296_, _23967_);
  nand (_08470_, _08468_, _08467_);
  nand (_08471_, _08470_, _01204_);
  nand (_08473_, _08471_, _08466_);
  nand (_08475_, _08473_, _01262_);
  nand (_08476_, _08475_, _08462_);
  nand (_08478_, _08476_, _01274_);
  nand (_08480_, _08478_, _08446_);
  nand (_08481_, _08480_, _01308_);
  nand (_08483_, _01290_, _23924_);
  nand (_08485_, _01296_, _23910_);
  nand (_08486_, _08485_, _08483_);
  nand (_08488_, _08486_, _01204_);
  nand (_08490_, _01296_, _23881_);
  nand (_08491_, _01290_, _23895_);
  nand (_08493_, _08491_, _08490_);
  nand (_08495_, _08493_, _01206_);
  nand (_08496_, _08495_, _08488_);
  nand (_08498_, _08496_, _01260_);
  nand (_08500_, _01290_, _23867_);
  nand (_08501_, _01296_, _23852_);
  nand (_08503_, _08501_, _08500_);
  nand (_08505_, _08503_, _01204_);
  nand (_08507_, _01296_, _23824_);
  nand (_08509_, _01290_, _23838_);
  nand (_08511_, _08509_, _08507_);
  nand (_08513_, _08511_, _01206_);
  nand (_08514_, _08513_, _08505_);
  nand (_08516_, _08514_, _01262_);
  nand (_08518_, _08516_, _08498_);
  nand (_08519_, _08518_, _01275_);
  nor (_08521_, _01296_, _23809_);
  nor (_08522_, _01290_, _23795_);
  nor (_08524_, _08522_, _08521_);
  nand (_08526_, _08524_, _01204_);
  nor (_08527_, _01290_, _23766_);
  nor (_08529_, _01296_, _23780_);
  nor (_08531_, _08529_, _08527_);
  nand (_08532_, _08531_, _01206_);
  nand (_08534_, _08532_, _08526_);
  nand (_08536_, _08534_, _01260_);
  nor (_08537_, _01296_, _23752_);
  nor (_08539_, _01290_, _23737_);
  nor (_08541_, _08539_, _08537_);
  nand (_08542_, _08541_, _01204_);
  nor (_08544_, _01290_, _23709_);
  nor (_08546_, _01296_, _23723_);
  nor (_08547_, _08546_, _08544_);
  nand (_08549_, _08547_, _01206_);
  nand (_08551_, _08549_, _08542_);
  nand (_08552_, _08551_, _01262_);
  nand (_08554_, _08552_, _08536_);
  nand (_08555_, _08554_, _01274_);
  nand (_08557_, _08555_, _08519_);
  nand (_08559_, _08557_, _01241_);
  nand (_08560_, _08559_, _08481_);
  nand (_08561_, _08560_, _01245_);
  nor (_08562_, _01296_, _24212_);
  nor (_08563_, _01290_, _24198_);
  nor (_08564_, _08563_, _08562_);
  nand (_08566_, _08564_, _01204_);
  nor (_08568_, _01290_, _24169_);
  nor (_08569_, _01296_, _24183_);
  nor (_08571_, _08569_, _08568_);
  nand (_08574_, _08571_, _01206_);
  nand (_08575_, _08574_, _08566_);
  nand (_08577_, _08575_, _01262_);
  nor (_08579_, _01296_, _24269_);
  nor (_08580_, _01290_, _24255_);
  nor (_08581_, _08580_, _08579_);
  nand (_08582_, _08581_, _01204_);
  nor (_08583_, _01290_, _24226_);
  nor (_08584_, _01296_, _24241_);
  nor (_08585_, _08584_, _08583_);
  nand (_08586_, _08585_, _01206_);
  nand (_08587_, _08586_, _08582_);
  nand (_08588_, _08587_, _01260_);
  nand (_08589_, _08588_, _08577_);
  nand (_08590_, _08589_, _01274_);
  nand (_08591_, _01290_, _24327_);
  nand (_08592_, _01296_, _24312_);
  nand (_08593_, _08592_, _08591_);
  nand (_08594_, _08593_, _01204_);
  nand (_08595_, _01296_, _24284_);
  nand (_08596_, _01290_, _24298_);
  nand (_08597_, _08596_, _08595_);
  nand (_08598_, _08597_, _01206_);
  nand (_08599_, _08598_, _08594_);
  nand (_08600_, _08599_, _01262_);
  nand (_08601_, _01290_, _24384_);
  nand (_08602_, _01296_, _24370_);
  nand (_08603_, _08602_, _08601_);
  nand (_08604_, _08603_, _01204_);
  nand (_08605_, _01296_, _24341_);
  nand (_08606_, _01290_, _24355_);
  nand (_08607_, _08606_, _08605_);
  nand (_08608_, _08607_, _01206_);
  nand (_08609_, _08608_, _08604_);
  nand (_08610_, _08609_, _01260_);
  nand (_08611_, _08610_, _08600_);
  nand (_08612_, _08611_, _01275_);
  nand (_08613_, _08612_, _08590_);
  nand (_08614_, _08613_, _01241_);
  nor (_08615_, _01296_, _24413_);
  nor (_08617_, _01290_, _24399_);
  nor (_08618_, _08617_, _08615_);
  nand (_08619_, _08618_, _01206_);
  nand (_08620_, _01290_, _24442_);
  nand (_08621_, _01296_, _24427_);
  nand (_08622_, _08621_, _08620_);
  nand (_08623_, _08622_, _01204_);
  nand (_08624_, _08623_, _08619_);
  nand (_08625_, _08624_, _01262_);
  nor (_08626_, _01296_, _24470_);
  nor (_08627_, _01290_, _24456_);
  nor (_08628_, _08627_, _08626_);
  nand (_08629_, _08628_, _01206_);
  nand (_08630_, _01290_, _24499_);
  nand (_08631_, _01296_, _24485_);
  nand (_08632_, _08631_, _08630_);
  nand (_08633_, _08632_, _01204_);
  nand (_08634_, _08633_, _08629_);
  nand (_08635_, _08634_, _01260_);
  nand (_08636_, _08635_, _08625_);
  nand (_08637_, _08636_, _01274_);
  nand (_08638_, _01296_, _24543_);
  nand (_08639_, _01290_, _24557_);
  nand (_08640_, _08639_, _08638_);
  nand (_08641_, _08640_, _01204_);
  nand (_08642_, _01290_, _24529_);
  nand (_08643_, _01296_, _24513_);
  nand (_08644_, _08643_, _08642_);
  nand (_08645_, _08644_, _01206_);
  nand (_08646_, _08645_, _08641_);
  nand (_08647_, _08646_, _01262_);
  nand (_08648_, _01296_, _24600_);
  nand (_08649_, _01290_, _24615_);
  nand (_08650_, _08649_, _08648_);
  nand (_08651_, _08650_, _01204_);
  nand (_08652_, _01290_, _24586_);
  nand (_08653_, _01296_, _24572_);
  nand (_08654_, _08653_, _08652_);
  nand (_08655_, _08654_, _01206_);
  nand (_08656_, _08655_, _08651_);
  nand (_08658_, _08656_, _01260_);
  nand (_08659_, _08658_, _08647_);
  nand (_08660_, _08659_, _01275_);
  nand (_08661_, _08660_, _08637_);
  nand (_08662_, _08661_, _01308_);
  nand (_08663_, _08662_, _08614_);
  nand (_08664_, _08663_, _01244_);
  nand (_08665_, _08664_, _08561_);
  nor (_08666_, _08665_, _01235_);
  nor (_08667_, _08666_, _08406_);
  nor (_08668_, _08667_, _28718_);
  nor (_08669_, _08668_, _08187_);
  nor (_08670_, _08669_, _06280_);
  nand (_08671_, _06280_, _27105_);
  nand (_08672_, _08671_, _29344_);
  nor (_15104_, _08672_, _08670_);
  nand (_08673_, _01290_, _27561_);
  nand (_08674_, _01296_, _27531_);
  nand (_08675_, _08674_, _08673_);
  nand (_08676_, _08675_, _01204_);
  nand (_08677_, _01296_, _23600_);
  nand (_08678_, _01290_, _27503_);
  nand (_08679_, _08678_, _08677_);
  nand (_08680_, _08679_, _01206_);
  nand (_08681_, _08680_, _08676_);
  nand (_08682_, _08681_, _01260_);
  nand (_08683_, _01290_, _23694_);
  nand (_08684_, _01296_, _23614_);
  nand (_08685_, _08684_, _08683_);
  nand (_08686_, _08685_, _01204_);
  nand (_08687_, _01296_, _27446_);
  nand (_08688_, _01290_, _27475_);
  nand (_08689_, _08688_, _08687_);
  nand (_08690_, _08689_, _01206_);
  nand (_08691_, _08690_, _08686_);
  nand (_08692_, _08691_, _01262_);
  nand (_08693_, _08692_, _08682_);
  nand (_08694_, _08693_, _01275_);
  nor (_08695_, _01296_, _27418_);
  nor (_08697_, _01290_, _27390_);
  nor (_08700_, _08697_, _08695_);
  nand (_08701_, _08700_, _01204_);
  nor (_08703_, _01290_, _27333_);
  nor (_08705_, _01296_, _27361_);
  nor (_08706_, _08705_, _08703_);
  nand (_08708_, _08706_, _01206_);
  nand (_08710_, _08708_, _08701_);
  nand (_08712_, _08710_, _01260_);
  nor (_08714_, _01296_, _27305_);
  nor (_08715_, _01290_, _27276_);
  nor (_08716_, _08715_, _08714_);
  nand (_08717_, _08716_, _01204_);
  nor (_08718_, _01290_, _27220_);
  nor (_08719_, _01296_, _27248_);
  nor (_08720_, _08719_, _08718_);
  nand (_08721_, _08720_, _01206_);
  nand (_08722_, _08721_, _08717_);
  nand (_08723_, _08722_, _01262_);
  nand (_08724_, _08723_, _08712_);
  nand (_08725_, _08724_, _01274_);
  nand (_08726_, _08725_, _08694_);
  nand (_08727_, _08726_, _01241_);
  nand (_08728_, _01296_, _23557_);
  nand (_08730_, _01290_, _27929_);
  nand (_08732_, _08730_, _08728_);
  nand (_08733_, _08732_, _01204_);
  nand (_08735_, _01290_, _27901_);
  nand (_08737_, _01296_, _23571_);
  nand (_08738_, _08737_, _08735_);
  nand (_08739_, _08738_, _01206_);
  nand (_08740_, _08739_, _08733_);
  nand (_08741_, _08740_, _01260_);
  nand (_08742_, _01296_, _27844_);
  nand (_08743_, _01290_, _27873_);
  nand (_08744_, _08743_, _08742_);
  nand (_08745_, _08744_, _01204_);
  nand (_08746_, _01290_, _27816_);
  nand (_08747_, _01296_, _27788_);
  nand (_08748_, _08747_, _08746_);
  nand (_08749_, _08748_, _01206_);
  nand (_08751_, _08749_, _08745_);
  nand (_08752_, _08751_, _01262_);
  nand (_08753_, _08752_, _08741_);
  nand (_08754_, _08753_, _01275_);
  nor (_08755_, _01296_, _27703_);
  nor (_08756_, _01290_, _27674_);
  nor (_08757_, _08756_, _08755_);
  nand (_08758_, _08757_, _01206_);
  nand (_08759_, _01290_, _27759_);
  nand (_08760_, _01296_, _27731_);
  nand (_08761_, _08760_, _08759_);
  nand (_08762_, _08761_, _01204_);
  nand (_08763_, _08762_, _08758_);
  nand (_08764_, _08763_, _01260_);
  nor (_08765_, _01296_, _27617_);
  nor (_08766_, _01290_, _27589_);
  nor (_08767_, _08766_, _08765_);
  nand (_08768_, _08767_, _01206_);
  nand (_08769_, _01290_, _23586_);
  nand (_08770_, _01296_, _27646_);
  nand (_08771_, _08770_, _08769_);
  nand (_08772_, _08771_, _01204_);
  nand (_08773_, _08772_, _08768_);
  nand (_08774_, _08773_, _01262_);
  nand (_08775_, _08774_, _08764_);
  nand (_08776_, _08775_, _01274_);
  nand (_08777_, _08776_, _08754_);
  nand (_08778_, _08777_, _01308_);
  nand (_08779_, _08778_, _08727_);
  nand (_08780_, _08779_, _01245_);
  nand (_08781_, _01296_, _28384_);
  nand (_08782_, _01290_, _28412_);
  nand (_08783_, _08782_, _08781_);
  nand (_08784_, _08783_, _01204_);
  nand (_08785_, _01290_, _28356_);
  nand (_08786_, _01296_, _28298_);
  nand (_08787_, _08786_, _08785_);
  nand (_08788_, _08787_, _01206_);
  nand (_08789_, _08788_, _08784_);
  nand (_08790_, _08789_, _01260_);
  nand (_08793_, _01296_, _28241_);
  nand (_08794_, _01290_, _28270_);
  nand (_08795_, _08794_, _08793_);
  nand (_08796_, _08795_, _01204_);
  nand (_08797_, _01290_, _28184_);
  nand (_08798_, _01296_, _28156_);
  nand (_08799_, _08798_, _08797_);
  nand (_08800_, _08799_, _01206_);
  nand (_08801_, _08800_, _08796_);
  nand (_08802_, _08801_, _01262_);
  nand (_08803_, _08802_, _08790_);
  nand (_08804_, _08803_, _01275_);
  nor (_08805_, _01296_, _28071_);
  nor (_08806_, _01290_, _23500_);
  nor (_08807_, _08806_, _08805_);
  nand (_08808_, _08807_, _01206_);
  nand (_08810_, _01290_, _28128_);
  nand (_08812_, _01296_, _28099_);
  nand (_08813_, _08812_, _08810_);
  nand (_08815_, _08813_, _01204_);
  nand (_08817_, _08815_, _08808_);
  nand (_08819_, _08817_, _01260_);
  nor (_08821_, _01296_, _23456_);
  nor (_08822_, _01290_, _23442_);
  nor (_08823_, _08822_, _08821_);
  nand (_08824_, _08823_, _01206_);
  nand (_08826_, _01290_, _23485_);
  nand (_08828_, _01296_, _23471_);
  nand (_08829_, _08828_, _08826_);
  nand (_08831_, _08829_, _01204_);
  nand (_08833_, _08831_, _08824_);
  nand (_08834_, _08833_, _01262_);
  nand (_08836_, _08834_, _08819_);
  nand (_08838_, _08836_, _01274_);
  nand (_08839_, _08838_, _08804_);
  nand (_08840_, _08839_, _01308_);
  nand (_08841_, _01290_, _23428_);
  nand (_08842_, _01296_, _23413_);
  nand (_08843_, _08842_, _08841_);
  nand (_08844_, _08843_, _01204_);
  nand (_08846_, _01296_, _23385_);
  nand (_08848_, _01290_, _23399_);
  nand (_08850_, _08848_, _08846_);
  nand (_08851_, _08850_, _01206_);
  nand (_08853_, _08851_, _08844_);
  nand (_08855_, _08853_, _01260_);
  nand (_08856_, _01290_, _23370_);
  nand (_08857_, _01296_, _23356_);
  nand (_08858_, _08857_, _08856_);
  nand (_08860_, _08858_, _01204_);
  nand (_08862_, _01296_, _28213_);
  nand (_08863_, _01290_, _28457_);
  nand (_08865_, _08863_, _08862_);
  nand (_08867_, _08865_, _01206_);
  nand (_08868_, _08867_, _08860_);
  nand (_08869_, _08868_, _01262_);
  nand (_08870_, _08869_, _08855_);
  nand (_08871_, _08870_, _01275_);
  nor (_08872_, _01296_, _28326_);
  nor (_08873_, _01290_, _23528_);
  nor (_08874_, _08873_, _08872_);
  nand (_08875_, _08874_, _01204_);
  nor (_08877_, _01290_, _28043_);
  nor (_08879_, _01296_, _23514_);
  nor (_08880_, _08879_, _08877_);
  nand (_08881_, _08880_, _01206_);
  nand (_08882_, _08881_, _08875_);
  nand (_08883_, _08882_, _01260_);
  nor (_08884_, _01296_, _28014_);
  nor (_08885_, _01290_, _27986_);
  nor (_08886_, _08885_, _08884_);
  nand (_08887_, _08886_, _01204_);
  nor (_08888_, _01290_, _23543_);
  nor (_08889_, _01296_, _27958_);
  nor (_08890_, _08889_, _08888_);
  nand (_08891_, _08890_, _01206_);
  nand (_08892_, _08891_, _08887_);
  nand (_08893_, _08892_, _01262_);
  nand (_08894_, _08893_, _08883_);
  nand (_08896_, _08894_, _01274_);
  nand (_08899_, _08896_, _08871_);
  nand (_08901_, _08899_, _01241_);
  nand (_08903_, _08901_, _08840_);
  nand (_08904_, _08903_, _01244_);
  nand (_08906_, _08904_, _08780_);
  nor (_08908_, _08906_, _01231_);
  nand (_08909_, _01296_, _26255_);
  nand (_08910_, _01290_, _26283_);
  nand (_08912_, _08910_, _08909_);
  nand (_08914_, _08912_, _01204_);
  nand (_08915_, _01290_, _26226_);
  nand (_08917_, _01296_, _26198_);
  nand (_08919_, _08917_, _08915_);
  nand (_08920_, _08919_, _01206_);
  nand (_08922_, _08920_, _08914_);
  nand (_08924_, _08922_, _01260_);
  nand (_08925_, _01296_, _26141_);
  nand (_08927_, _01290_, _26170_);
  nand (_08929_, _08927_, _08925_);
  nand (_08930_, _08929_, _01204_);
  nand (_08931_, _01290_, _26113_);
  nand (_08933_, _01296_, _26085_);
  nand (_08935_, _08933_, _08931_);
  nand (_08937_, _08935_, _01206_);
  nand (_08939_, _08937_, _08930_);
  nand (_08940_, _08939_, _01262_);
  nand (_08941_, _08940_, _08924_);
  nand (_08943_, _08941_, _01275_);
  nor (_08945_, _01296_, _26000_);
  nor (_08946_, _01290_, _25971_);
  nor (_08947_, _08946_, _08945_);
  nand (_08948_, _08947_, _01206_);
  nand (_08949_, _01290_, _26056_);
  nand (_08951_, _01296_, _26028_);
  nand (_08953_, _08951_, _08949_);
  nand (_08954_, _08953_, _01204_);
  nand (_08955_, _08954_, _08948_);
  nand (_08956_, _08955_, _01260_);
  nor (_08957_, _01296_, _25885_);
  nor (_08958_, _01290_, _25857_);
  nor (_08960_, _08958_, _08957_);
  nand (_08961_, _08960_, _01206_);
  nand (_08962_, _01290_, _25943_);
  nand (_08963_, _01296_, _25913_);
  nand (_08964_, _08963_, _08962_);
  nand (_08965_, _08964_, _01204_);
  nand (_08966_, _08965_, _08961_);
  nand (_08967_, _08966_, _01262_);
  nand (_08968_, _08967_, _08956_);
  nand (_08970_, _08968_, _01274_);
  nand (_08972_, _08970_, _08943_);
  nand (_08973_, _08972_, _01308_);
  nand (_08974_, _01290_, _25828_);
  nand (_08975_, _01296_, _25800_);
  nand (_08976_, _08975_, _08974_);
  nand (_08977_, _08976_, _01204_);
  nand (_08978_, _01296_, _25743_);
  nand (_08979_, _01290_, _25772_);
  nand (_08981_, _08979_, _08978_);
  nand (_08983_, _08981_, _01206_);
  nand (_08984_, _08983_, _08977_);
  nand (_08985_, _08984_, _01260_);
  nand (_08987_, _01290_, _25715_);
  nand (_08989_, _01296_, _25687_);
  nand (_08990_, _08989_, _08987_);
  nand (_08991_, _08990_, _01204_);
  nand (_08992_, _01296_, _25630_);
  nand (_08994_, _01290_, _25658_);
  nand (_08996_, _08994_, _08992_);
  nand (_08997_, _08996_, _01206_);
  nand (_08999_, _08997_, _08991_);
  nand (_09001_, _08999_, _01262_);
  nand (_09002_, _09001_, _08985_);
  nand (_09004_, _09002_, _01275_);
  nor (_09006_, _01296_, _25602_);
  nor (_09007_, _01290_, _25580_);
  nor (_09008_, _09007_, _09006_);
  nand (_09009_, _09008_, _01204_);
  nor (_09011_, _01290_, _25552_);
  nor (_09013_, _01296_, _25566_);
  nor (_09015_, _09013_, _09011_);
  nand (_09017_, _09015_, _01206_);
  nand (_09019_, _09017_, _09009_);
  nand (_09020_, _09019_, _01260_);
  nor (_09022_, _01296_, _25537_);
  nor (_09024_, _01290_, _25523_);
  nor (_09025_, _09024_, _09022_);
  nand (_09026_, _09025_, _01204_);
  nor (_09027_, _01290_, _25494_);
  nor (_09028_, _01296_, _25509_);
  nor (_09029_, _09028_, _09027_);
  nand (_09030_, _09029_, _01206_);
  nand (_09031_, _09030_, _09026_);
  nand (_09033_, _09031_, _01262_);
  nand (_09035_, _09033_, _09020_);
  nand (_09036_, _09035_, _01274_);
  nand (_09038_, _09036_, _09004_);
  nand (_09040_, _09038_, _01241_);
  nand (_09041_, _09040_, _08973_);
  nand (_09042_, _09041_, _01245_);
  nor (_09044_, _01296_, _26396_);
  nor (_09046_, _01290_, _26368_);
  nor (_09047_, _09046_, _09044_);
  nand (_09049_, _09047_, _01204_);
  nor (_09051_, _01290_, _26311_);
  nor (_09052_, _01296_, _26340_);
  nor (_09053_, _09052_, _09051_);
  nand (_09055_, _09053_, _01206_);
  nand (_09057_, _09055_, _09049_);
  nand (_09059_, _09057_, _01262_);
  nor (_09061_, _01296_, _26510_);
  nor (_09062_, _01290_, _26481_);
  nor (_09063_, _09062_, _09061_);
  nand (_09064_, _09063_, _01204_);
  nor (_09065_, _01290_, _26425_);
  nor (_09066_, _01296_, _26453_);
  nor (_09067_, _09066_, _09065_);
  nand (_09068_, _09067_, _01206_);
  nand (_09069_, _09068_, _09064_);
  nand (_09070_, _09069_, _01260_);
  nand (_09072_, _09070_, _09059_);
  nand (_09073_, _09072_, _01274_);
  nand (_09074_, _01290_, _26623_);
  nand (_09075_, _01296_, _26595_);
  nand (_09076_, _09075_, _09074_);
  nand (_09077_, _09076_, _01204_);
  nand (_09078_, _01296_, _26538_);
  nand (_09079_, _01290_, _26567_);
  nand (_09080_, _09079_, _09078_);
  nand (_09081_, _09080_, _01206_);
  nand (_09082_, _09081_, _09077_);
  nand (_09083_, _09082_, _01262_);
  nand (_09084_, _01290_, _26738_);
  nand (_09085_, _01296_, _26708_);
  nand (_09086_, _09085_, _09084_);
  nand (_09087_, _09086_, _01204_);
  nand (_09088_, _01296_, _26652_);
  nand (_09089_, _01290_, _26680_);
  nand (_09090_, _09089_, _09088_);
  nand (_09091_, _09090_, _01206_);
  nand (_09092_, _09091_, _09087_);
  nand (_09093_, _09092_, _01260_);
  nand (_09094_, _09093_, _09083_);
  nand (_09095_, _09094_, _01275_);
  nand (_09096_, _09095_, _09073_);
  nand (_09097_, _09096_, _01241_);
  nor (_09098_, _01296_, _26794_);
  nor (_09099_, _01290_, _26766_);
  nor (_09100_, _09099_, _09098_);
  nand (_09101_, _09100_, _01206_);
  nand (_09102_, _01290_, _26851_);
  nand (_09103_, _01296_, _26823_);
  nand (_09104_, _09103_, _09102_);
  nand (_09105_, _09104_, _01204_);
  nand (_09106_, _09105_, _09101_);
  nand (_09107_, _09106_, _01262_);
  nor (_09108_, _01296_, _26908_);
  nor (_09109_, _01290_, _26879_);
  nor (_09110_, _09109_, _09108_);
  nand (_09111_, _09110_, _01206_);
  nand (_09113_, _01290_, _26964_);
  nand (_09114_, _01296_, _26936_);
  nand (_09115_, _09114_, _09113_);
  nand (_09116_, _09115_, _01204_);
  nand (_09117_, _09116_, _09111_);
  nand (_09118_, _09117_, _01260_);
  nand (_09119_, _09118_, _09107_);
  nand (_09120_, _09119_, _01274_);
  nand (_09121_, _01296_, _27049_);
  nand (_09122_, _01290_, _27078_);
  nand (_09123_, _09122_, _09121_);
  nand (_09124_, _09123_, _01204_);
  nand (_09125_, _01290_, _27021_);
  nand (_09126_, _01296_, _26993_);
  nand (_09127_, _09126_, _09125_);
  nand (_09128_, _09127_, _01206_);
  nand (_09129_, _09128_, _09124_);
  nand (_09130_, _09129_, _01262_);
  nand (_09131_, _01296_, _27163_);
  nand (_09132_, _01290_, _27191_);
  nand (_09133_, _09132_, _09131_);
  nand (_09134_, _09133_, _01204_);
  nand (_09135_, _01290_, _27135_);
  nand (_09136_, _01296_, _27106_);
  nand (_09137_, _09136_, _09135_);
  nand (_09138_, _09137_, _01206_);
  nand (_09139_, _09138_, _09134_);
  nand (_09140_, _09139_, _01260_);
  nand (_09141_, _09140_, _09130_);
  nand (_09142_, _09141_, _01275_);
  nand (_09143_, _09142_, _09120_);
  nand (_09145_, _09143_, _01308_);
  nand (_09146_, _09145_, _09097_);
  nand (_09148_, _09146_, _01244_);
  nand (_09149_, _09148_, _09042_);
  nor (_09151_, _09149_, _01235_);
  nor (_09152_, _09151_, _08908_);
  nor (_09154_, _09152_, _28717_);
  nand (_09155_, _01290_, _24846_);
  nand (_09157_, _01296_, _24832_);
  nand (_09159_, _09157_, _09155_);
  nand (_09161_, _09159_, _01204_);
  nand (_09162_, _01296_, _24803_);
  nand (_09164_, _01290_, _24818_);
  nand (_09165_, _09164_, _09162_);
  nand (_09166_, _09165_, _01206_);
  nand (_09167_, _09166_, _09161_);
  nand (_09168_, _09167_, _01260_);
  nand (_09169_, _01290_, _24789_);
  nand (_09170_, _01296_, _24775_);
  nand (_09171_, _09170_, _09169_);
  nand (_09172_, _09171_, _01204_);
  nand (_09173_, _01296_, _24746_);
  nand (_09174_, _01290_, _24760_);
  nand (_09175_, _09174_, _09173_);
  nand (_09176_, _09175_, _01206_);
  nand (_09177_, _09176_, _09172_);
  nand (_09178_, _09177_, _01262_);
  nand (_09179_, _09178_, _09168_);
  nand (_09181_, _09179_, _01275_);
  nor (_09182_, _01296_, _24732_);
  nor (_09184_, _01290_, _24717_);
  nor (_09185_, _09184_, _09182_);
  nand (_09187_, _09185_, _01204_);
  nor (_09188_, _01290_, _24689_);
  nor (_09190_, _01296_, _24703_);
  nor (_09191_, _09190_, _09188_);
  nand (_09193_, _09191_, _01206_);
  nand (_09194_, _09193_, _09187_);
  nand (_09196_, _09194_, _01260_);
  nor (_09197_, _01296_, _24674_);
  nor (_09199_, _01290_, _24660_);
  nor (_09200_, _09199_, _09197_);
  nand (_09201_, _09200_, _01204_);
  nor (_09202_, _01290_, _24631_);
  nor (_09203_, _01296_, _24646_);
  nor (_09204_, _09203_, _09202_);
  nand (_09205_, _09204_, _01206_);
  nand (_09206_, _09205_, _09201_);
  nand (_09207_, _09206_, _01262_);
  nand (_09209_, _09207_, _09196_);
  nand (_09210_, _09209_, _01274_);
  nand (_09211_, _09210_, _09181_);
  nand (_09212_, _09211_, _01241_);
  nand (_09213_, _01296_, _25063_);
  nand (_09214_, _01290_, _25077_);
  nand (_09215_, _09214_, _09213_);
  nand (_09217_, _09215_, _01204_);
  nand (_09218_, _01290_, _25048_);
  nand (_09220_, _01296_, _25034_);
  nand (_09221_, _09220_, _09218_);
  nand (_09223_, _09221_, _01206_);
  nand (_09224_, _09223_, _09217_);
  nand (_09226_, _09224_, _01260_);
  nand (_09227_, _01296_, _25005_);
  nand (_09229_, _01290_, _25020_);
  nand (_09230_, _09229_, _09227_);
  nand (_09232_, _09230_, _01204_);
  nand (_09233_, _01290_, _24991_);
  nand (_09235_, _01296_, _24977_);
  nand (_09236_, _09235_, _09233_);
  nand (_09237_, _09236_, _01206_);
  nand (_09238_, _09237_, _09232_);
  nand (_09239_, _09238_, _01262_);
  nand (_09240_, _09239_, _09226_);
  nand (_09241_, _09240_, _01275_);
  nor (_09242_, _01296_, _24934_);
  nor (_09243_, _01290_, _24918_);
  nor (_09244_, _09243_, _09242_);
  nand (_09245_, _09244_, _01206_);
  nand (_09246_, _01290_, _24962_);
  nand (_09247_, _01296_, _24948_);
  nand (_09248_, _09247_, _09246_);
  nand (_09249_, _09248_, _01204_);
  nand (_09250_, _09249_, _09245_);
  nand (_09252_, _09250_, _01260_);
  nor (_09253_, _01296_, _24875_);
  nor (_09255_, _01290_, _24861_);
  nor (_09256_, _09255_, _09253_);
  nand (_09258_, _09256_, _01206_);
  nand (_09260_, _01290_, _24904_);
  nand (_09262_, _01296_, _24889_);
  nand (_09263_, _09262_, _09260_);
  nand (_09265_, _09263_, _01204_);
  nand (_09266_, _09265_, _09258_);
  nand (_09268_, _09266_, _01262_);
  nand (_09269_, _09268_, _09252_);
  nand (_09271_, _09269_, _01274_);
  nand (_09272_, _09271_, _09241_);
  nand (_09273_, _09272_, _01308_);
  nand (_09274_, _09273_, _09212_);
  nand (_09275_, _09274_, _01245_);
  nand (_09276_, _01296_, _25465_);
  nand (_09277_, _01290_, _25480_);
  nand (_09278_, _09277_, _09276_);
  nand (_09279_, _09278_, _01204_);
  nand (_09280_, _01290_, _25451_);
  nand (_09281_, _01296_, _25437_);
  nand (_09282_, _09281_, _09280_);
  nand (_09283_, _09282_, _01206_);
  nand (_09284_, _09283_, _09279_);
  nand (_09285_, _09284_, _01260_);
  nand (_09286_, _01296_, _25408_);
  nand (_09288_, _01290_, _25422_);
  nand (_09289_, _09288_, _09286_);
  nand (_09291_, _09289_, _01204_);
  nand (_09292_, _01290_, _25394_);
  nand (_09294_, _01296_, _25379_);
  nand (_09295_, _09294_, _09292_);
  nand (_09297_, _09295_, _01206_);
  nand (_09298_, _09297_, _09291_);
  nand (_09300_, _09298_, _01262_);
  nand (_09301_, _09300_, _09285_);
  nand (_09303_, _09301_, _01275_);
  nor (_09304_, _01296_, _25335_);
  nor (_09306_, _01290_, _25321_);
  nor (_09307_, _09306_, _09304_);
  nand (_09308_, _09307_, _01206_);
  nand (_09309_, _01290_, _25365_);
  nand (_09310_, _01296_, _25351_);
  nand (_09313_, _09310_, _09309_);
  nand (_09314_, _09313_, _01204_);
  nand (_09315_, _09314_, _09308_);
  nand (_09316_, _09315_, _01260_);
  nor (_09317_, _01296_, _25278_);
  nor (_09318_, _01290_, _25264_);
  nor (_09319_, _09318_, _09317_);
  nand (_09320_, _09319_, _01206_);
  nand (_09321_, _01290_, _25307_);
  nand (_09322_, _01296_, _25292_);
  nand (_09323_, _09322_, _09321_);
  nand (_09325_, _09323_, _01204_);
  nand (_09326_, _09325_, _09320_);
  nand (_09328_, _09326_, _01262_);
  nand (_09329_, _09328_, _09316_);
  nand (_09331_, _09329_, _01274_);
  nand (_09332_, _09331_, _09303_);
  nand (_09334_, _09332_, _01308_);
  nand (_09335_, _01290_, _25249_);
  nand (_09337_, _01296_, _25235_);
  nand (_09338_, _09337_, _09335_);
  nand (_09340_, _09338_, _01204_);
  nand (_09341_, _01296_, _25206_);
  nand (_09343_, _01290_, _25221_);
  nand (_09344_, _09343_, _09341_);
  nand (_09345_, _09344_, _01206_);
  nand (_09346_, _09345_, _09340_);
  nand (_09347_, _09346_, _01260_);
  nand (_09348_, _01290_, _25192_);
  nand (_09349_, _01296_, _25177_);
  nand (_09350_, _09349_, _09348_);
  nand (_09351_, _09350_, _01204_);
  nand (_09352_, _01296_, _25149_);
  nand (_09353_, _01290_, _25163_);
  nand (_09354_, _09353_, _09352_);
  nand (_09355_, _09354_, _01206_);
  nand (_09356_, _09355_, _09351_);
  nand (_09357_, _09356_, _01262_);
  nand (_09358_, _09357_, _09347_);
  nand (_09360_, _09358_, _01275_);
  nor (_09362_, _01296_, _25134_);
  nor (_09364_, _01290_, _25120_);
  nor (_09365_, _09364_, _09362_);
  nand (_09367_, _09365_, _01204_);
  nor (_09368_, _01290_, _23672_);
  nor (_09370_, _01296_, _25106_);
  nor (_09371_, _09370_, _09368_);
  nand (_09373_, _09371_, _01206_);
  nand (_09374_, _09373_, _09367_);
  nand (_09376_, _09374_, _01260_);
  nor (_09377_, _01296_, _23643_);
  nor (_09379_, _01290_, _23629_);
  nor (_09380_, _09379_, _09377_);
  nand (_09381_, _09380_, _01204_);
  nor (_09382_, _01290_, _25091_);
  nor (_09383_, _01296_, _23657_);
  nor (_09384_, _09383_, _09382_);
  nand (_09385_, _09384_, _01206_);
  nand (_09386_, _09385_, _09381_);
  nand (_09387_, _09386_, _01262_);
  nand (_09388_, _09387_, _09376_);
  nand (_09389_, _09388_, _01274_);
  nand (_09390_, _09389_, _09360_);
  nand (_09391_, _09390_, _01241_);
  nand (_09392_, _09391_, _09334_);
  nand (_09393_, _09392_, _01244_);
  nand (_09394_, _09393_, _09275_);
  nor (_09396_, _09394_, _01231_);
  nand (_09397_, _01296_, _24142_);
  nand (_09399_, _01290_, _24157_);
  nand (_09400_, _09399_, _09397_);
  nand (_09402_, _09400_, _01204_);
  nand (_09403_, _01290_, _24128_);
  nand (_09405_, _01296_, _24114_);
  nand (_09406_, _09405_, _09403_);
  nand (_09408_, _09406_, _01206_);
  nand (_09409_, _09408_, _09402_);
  nand (_09411_, _09409_, _01260_);
  nand (_09412_, _01296_, _24084_);
  nand (_09414_, _01290_, _24098_);
  nand (_09416_, _09414_, _09412_);
  nand (_09417_, _09416_, _01204_);
  nand (_09418_, _01290_, _24070_);
  nand (_09419_, _01296_, _24055_);
  nand (_09420_, _09419_, _09418_);
  nand (_09421_, _09420_, _01206_);
  nand (_09422_, _09421_, _09417_);
  nand (_09423_, _09422_, _01262_);
  nand (_09424_, _09423_, _09411_);
  nand (_09425_, _09424_, _01275_);
  nor (_09426_, _01296_, _24012_);
  nor (_09427_, _01290_, _23998_);
  nor (_09428_, _09427_, _09426_);
  nand (_09429_, _09428_, _01206_);
  nand (_09430_, _01290_, _24041_);
  nand (_09432_, _01296_, _24026_);
  nand (_09433_, _09432_, _09430_);
  nand (_09435_, _09433_, _01204_);
  nand (_09436_, _09435_, _09429_);
  nand (_09438_, _09436_, _01260_);
  nor (_09439_, _01296_, _23955_);
  nor (_09441_, _01290_, _23940_);
  nor (_09442_, _09441_, _09439_);
  nand (_09444_, _09442_, _01206_);
  nand (_09445_, _01290_, _23983_);
  nand (_09447_, _01296_, _23969_);
  nand (_09448_, _09447_, _09445_);
  nand (_09450_, _09448_, _01204_);
  nand (_09451_, _09450_, _09444_);
  nand (_09452_, _09451_, _01262_);
  nand (_09453_, _09452_, _09438_);
  nand (_09454_, _09453_, _01274_);
  nand (_09455_, _09454_, _09425_);
  nand (_09456_, _09455_, _01308_);
  nand (_09457_, _01290_, _23926_);
  nand (_09458_, _01296_, _23912_);
  nand (_09459_, _09458_, _09457_);
  nand (_09460_, _09459_, _01204_);
  nand (_09461_, _01296_, _23883_);
  nand (_09462_, _01290_, _23897_);
  nand (_09464_, _09462_, _09461_);
  nand (_09465_, _09464_, _01206_);
  nand (_09466_, _09465_, _09460_);
  nand (_09468_, _09466_, _01260_);
  nand (_09469_, _01290_, _23869_);
  nand (_09471_, _01296_, _23854_);
  nand (_09472_, _09471_, _09469_);
  nand (_09474_, _09472_, _01204_);
  nand (_09475_, _01296_, _23826_);
  nand (_09477_, _01290_, _23840_);
  nand (_09478_, _09477_, _09475_);
  nand (_09480_, _09478_, _01206_);
  nand (_09481_, _09480_, _09474_);
  nand (_09483_, _09481_, _01262_);
  nand (_09484_, _09483_, _09468_);
  nand (_09486_, _09484_, _01275_);
  nor (_09487_, _01296_, _23811_);
  nor (_09488_, _01290_, _23797_);
  nor (_09489_, _09488_, _09487_);
  nand (_09490_, _09489_, _01204_);
  nor (_09491_, _01290_, _23768_);
  nor (_09492_, _01296_, _23783_);
  nor (_09493_, _09492_, _09491_);
  nand (_09494_, _09493_, _01206_);
  nand (_09495_, _09494_, _09490_);
  nand (_09496_, _09495_, _01260_);
  nor (_09497_, _01296_, _23754_);
  nor (_09498_, _01290_, _23739_);
  nor (_09499_, _09498_, _09497_);
  nand (_09500_, _09499_, _01204_);
  nor (_09501_, _01290_, _23711_);
  nor (_09503_, _01296_, _23725_);
  nor (_09504_, _09503_, _09501_);
  nand (_09506_, _09504_, _01206_);
  nand (_09507_, _09506_, _09500_);
  nand (_09509_, _09507_, _01262_);
  nand (_09510_, _09509_, _09496_);
  nand (_09512_, _09510_, _01274_);
  nand (_09513_, _09512_, _09486_);
  nand (_09515_, _09513_, _01241_);
  nand (_09517_, _09515_, _09456_);
  nand (_09519_, _09517_, _01245_);
  nor (_09520_, _01296_, _24214_);
  nor (_09522_, _01290_, _24200_);
  nor (_09523_, _09522_, _09520_);
  nand (_09524_, _09523_, _01204_);
  nor (_09525_, _01290_, _24171_);
  nor (_09526_, _01296_, _24185_);
  nor (_09527_, _09526_, _09525_);
  nand (_09528_, _09527_, _01206_);
  nand (_09529_, _09528_, _09524_);
  nand (_09530_, _09529_, _01262_);
  nor (_09531_, _01296_, _24271_);
  nor (_09532_, _01290_, _24257_);
  nor (_09533_, _09532_, _09531_);
  nand (_09534_, _09533_, _01204_);
  nor (_09535_, _01290_, _24228_);
  nor (_09536_, _01296_, _24243_);
  nor (_09537_, _09536_, _09535_);
  nand (_09539_, _09537_, _01206_);
  nand (_09540_, _09539_, _09534_);
  nand (_09542_, _09540_, _01260_);
  nand (_09543_, _09542_, _09530_);
  nand (_09545_, _09543_, _01274_);
  nand (_09546_, _01290_, _24329_);
  nand (_09548_, _01296_, _24314_);
  nand (_09549_, _09548_, _09546_);
  nand (_09551_, _09549_, _01204_);
  nand (_09552_, _01296_, _24286_);
  nand (_09554_, _01290_, _24300_);
  nand (_09555_, _09554_, _09552_);
  nand (_09557_, _09555_, _01206_);
  nand (_09558_, _09557_, _09551_);
  nand (_09559_, _09558_, _01262_);
  nand (_09560_, _01290_, _24386_);
  nand (_09561_, _01296_, _24372_);
  nand (_09562_, _09561_, _09560_);
  nand (_09563_, _09562_, _01204_);
  nand (_09564_, _01296_, _24343_);
  nand (_09565_, _01290_, _24358_);
  nand (_09567_, _09565_, _09564_);
  nand (_09568_, _09567_, _01206_);
  nand (_09569_, _09568_, _09563_);
  nand (_09570_, _09569_, _01260_);
  nand (_09571_, _09570_, _09559_);
  nand (_09572_, _09571_, _01275_);
  nand (_09573_, _09572_, _09545_);
  nand (_09575_, _09573_, _01241_);
  nor (_09576_, _01296_, _24415_);
  nor (_09578_, _01290_, _24401_);
  nor (_09579_, _09578_, _09576_);
  nand (_09581_, _09579_, _01206_);
  nand (_09582_, _01290_, _24444_);
  nand (_09584_, _01296_, _24429_);
  nand (_09585_, _09584_, _09582_);
  nand (_09587_, _09585_, _01204_);
  nand (_09588_, _09587_, _09581_);
  nand (_09590_, _09588_, _01262_);
  nor (_09591_, _01296_, _24472_);
  nor (_09593_, _01290_, _24458_);
  nor (_09594_, _09593_, _09591_);
  nand (_09595_, _09594_, _01206_);
  nand (_09596_, _01290_, _24501_);
  nand (_09597_, _01296_, _24487_);
  nand (_09598_, _09597_, _09596_);
  nand (_09599_, _09598_, _01204_);
  nand (_09600_, _09599_, _09595_);
  nand (_09601_, _09600_, _01260_);
  nand (_09602_, _09601_, _09590_);
  nand (_09603_, _09602_, _01274_);
  nand (_09604_, _01296_, _24545_);
  nand (_09605_, _01290_, _24559_);
  nand (_09606_, _09605_, _09604_);
  nand (_09607_, _09606_, _01204_);
  nand (_09608_, _01290_, _24531_);
  nand (_09610_, _01296_, _24515_);
  nand (_09611_, _09610_, _09608_);
  nand (_09613_, _09611_, _01206_);
  nand (_09614_, _09613_, _09607_);
  nand (_09616_, _09614_, _01262_);
  nand (_09618_, _01296_, _24602_);
  nand (_09620_, _01290_, _24617_);
  nand (_09621_, _09620_, _09618_);
  nand (_09623_, _09621_, _01204_);
  nand (_09624_, _01290_, _24588_);
  nand (_09626_, _01296_, _24574_);
  nand (_09627_, _09626_, _09624_);
  nand (_09629_, _09627_, _01206_);
  nand (_09630_, _09629_, _09623_);
  nand (_09631_, _09630_, _01260_);
  nand (_09632_, _09631_, _09616_);
  nand (_09633_, _09632_, _01275_);
  nand (_09634_, _09633_, _09603_);
  nand (_09635_, _09634_, _01308_);
  nand (_09636_, _09635_, _09575_);
  nand (_09637_, _09636_, _01244_);
  nand (_09638_, _09637_, _09519_);
  nor (_09639_, _09638_, _01235_);
  nor (_09640_, _09639_, _09396_);
  nor (_09641_, _09640_, _28718_);
  nor (_09642_, _09641_, _09154_);
  nor (_09643_, _09642_, _06280_);
  nand (_09645_, _06280_, _28102_);
  nand (_09647_, _09645_, _29344_);
  nor (_15132_, _09647_, _09643_);
  nand (_09650_, _01290_, _27565_);
  nand (_09652_, _01296_, _27535_);
  nand (_09653_, _09652_, _09650_);
  nand (_09655_, _09653_, _01204_);
  nand (_09656_, _01296_, _23602_);
  nand (_09658_, _01290_, _27507_);
  nand (_09659_, _09658_, _09656_);
  nand (_09661_, _09659_, _01206_);
  nand (_09662_, _09661_, _09655_);
  nand (_09664_, _09662_, _01260_);
  nand (_09665_, _01290_, _23696_);
  nand (_09667_, _01296_, _23616_);
  nand (_09668_, _09667_, _09665_);
  nand (_09670_, _09668_, _01204_);
  nand (_09671_, _01296_, _27450_);
  nand (_09674_, _01290_, _27479_);
  nand (_09675_, _09674_, _09671_);
  nand (_09676_, _09675_, _01206_);
  nand (_09677_, _09676_, _09670_);
  nand (_09678_, _09677_, _01262_);
  nand (_09679_, _09678_, _09664_);
  nand (_09680_, _09679_, _01275_);
  nor (_09681_, _01296_, _27422_);
  nor (_09682_, _01290_, _27394_);
  nor (_09683_, _09682_, _09681_);
  nand (_09684_, _09683_, _01204_);
  nor (_09685_, _01290_, _27337_);
  nor (_09686_, _01296_, _27365_);
  nor (_09687_, _09686_, _09685_);
  nand (_09688_, _09687_, _01206_);
  nand (_09689_, _09688_, _09684_);
  nand (_09690_, _09689_, _01260_);
  nor (_09691_, _01296_, _27309_);
  nor (_09692_, _01290_, _27280_);
  nor (_09693_, _09692_, _09691_);
  nand (_09694_, _09693_, _01204_);
  nor (_09695_, _01290_, _27224_);
  nor (_09697_, _01296_, _27252_);
  nor (_09699_, _09697_, _09695_);
  nand (_09701_, _09699_, _01206_);
  nand (_09703_, _09701_, _09694_);
  nand (_09705_, _09703_, _01262_);
  nand (_09706_, _09705_, _09690_);
  nand (_09707_, _09706_, _01274_);
  nand (_09708_, _09707_, _09680_);
  nand (_09709_, _09708_, _01241_);
  nand (_09710_, _01296_, _23559_);
  nand (_09711_, _01290_, _27933_);
  nand (_09712_, _09711_, _09710_);
  nand (_09713_, _09712_, _01204_);
  nand (_09714_, _01290_, _27905_);
  nand (_09715_, _01296_, _23573_);
  nand (_09716_, _09715_, _09714_);
  nand (_09717_, _09716_, _01206_);
  nand (_09718_, _09717_, _09713_);
  nand (_09720_, _09718_, _01260_);
  nand (_09721_, _01296_, _27848_);
  nand (_09722_, _01290_, _27877_);
  nand (_09723_, _09722_, _09721_);
  nand (_09724_, _09723_, _01204_);
  nand (_09725_, _01290_, _27820_);
  nand (_09726_, _01296_, _27792_);
  nand (_09727_, _09726_, _09725_);
  nand (_09728_, _09727_, _01206_);
  nand (_09729_, _09728_, _09724_);
  nand (_09730_, _09729_, _01262_);
  nand (_09731_, _09730_, _09720_);
  nand (_09732_, _09731_, _01275_);
  nor (_09733_, _01296_, _27707_);
  nor (_09734_, _01290_, _27678_);
  nor (_09735_, _09734_, _09733_);
  nand (_09736_, _09735_, _01206_);
  nand (_09737_, _01290_, _27763_);
  nand (_09738_, _01296_, _27735_);
  nand (_09739_, _09738_, _09737_);
  nand (_09740_, _09739_, _01204_);
  nand (_09741_, _09740_, _09736_);
  nand (_09742_, _09741_, _01260_);
  nor (_09743_, _01296_, _27622_);
  nor (_09744_, _01290_, _27593_);
  nor (_09745_, _09744_, _09743_);
  nand (_09746_, _09745_, _01206_);
  nand (_09747_, _01290_, _23588_);
  nand (_09748_, _01296_, _27650_);
  nand (_09749_, _09748_, _09747_);
  nand (_09750_, _09749_, _01204_);
  nand (_09751_, _09750_, _09746_);
  nand (_09752_, _09751_, _01262_);
  nand (_09753_, _09752_, _09742_);
  nand (_09754_, _09753_, _01274_);
  nand (_09755_, _09754_, _09732_);
  nand (_09756_, _09755_, _01308_);
  nand (_09757_, _09756_, _09709_);
  nand (_09758_, _09757_, _01245_);
  nand (_09759_, _01296_, _28388_);
  nand (_09761_, _01290_, _28416_);
  nand (_09762_, _09761_, _09759_);
  nand (_09763_, _09762_, _01204_);
  nand (_09764_, _01290_, _28360_);
  nand (_09765_, _01296_, _28302_);
  nand (_09766_, _09765_, _09764_);
  nand (_09767_, _09766_, _01206_);
  nand (_09768_, _09767_, _09763_);
  nand (_09769_, _09768_, _01260_);
  nand (_09770_, _01296_, _28245_);
  nand (_09771_, _01290_, _28274_);
  nand (_09772_, _09771_, _09770_);
  nand (_09773_, _09772_, _01204_);
  nand (_09774_, _01290_, _28189_);
  nand (_09775_, _01296_, _28160_);
  nand (_09776_, _09775_, _09774_);
  nand (_09777_, _09776_, _01206_);
  nand (_09778_, _09777_, _09773_);
  nand (_09779_, _09778_, _01262_);
  nand (_09780_, _09779_, _09769_);
  nand (_09781_, _09780_, _01275_);
  nor (_09782_, _01296_, _28075_);
  nor (_09783_, _01290_, _23502_);
  nor (_09784_, _09783_, _09782_);
  nand (_09785_, _09784_, _01206_);
  nand (_09786_, _01290_, _28132_);
  nand (_09787_, _01296_, _28103_);
  nand (_09788_, _09787_, _09786_);
  nand (_09789_, _09788_, _01204_);
  nand (_09790_, _09789_, _09785_);
  nand (_09791_, _09790_, _01260_);
  nor (_09792_, _01296_, _23459_);
  nor (_09793_, _01290_, _23444_);
  nor (_09794_, _09793_, _09792_);
  nand (_09795_, _09794_, _01206_);
  nand (_09796_, _01290_, _23487_);
  nand (_09797_, _01296_, _23473_);
  nand (_09798_, _09797_, _09796_);
  nand (_09799_, _09798_, _01204_);
  nand (_09800_, _09799_, _09795_);
  nand (_09803_, _09800_, _01262_);
  nand (_09804_, _09803_, _09791_);
  nand (_09805_, _09804_, _01274_);
  nand (_09806_, _09805_, _09781_);
  nand (_09807_, _09806_, _01308_);
  nand (_09808_, _01290_, _23430_);
  nand (_09809_, _01296_, _23415_);
  nand (_09810_, _09809_, _09808_);
  nand (_09811_, _09810_, _01204_);
  nand (_09812_, _01296_, _23387_);
  nand (_09813_, _01290_, _23401_);
  nand (_09814_, _09813_, _09812_);
  nand (_09815_, _09814_, _01206_);
  nand (_09816_, _09815_, _09811_);
  nand (_09817_, _09816_, _01260_);
  nand (_09818_, _01290_, _23372_);
  nand (_09819_, _01296_, _23358_);
  nand (_09820_, _09819_, _09818_);
  nand (_09821_, _09820_, _01204_);
  nand (_09822_, _01296_, _28217_);
  nand (_09823_, _01290_, _28453_);
  nand (_09824_, _09823_, _09822_);
  nand (_09825_, _09824_, _01206_);
  nand (_09826_, _09825_, _09821_);
  nand (_09827_, _09826_, _01262_);
  nand (_09828_, _09827_, _09817_);
  nand (_09829_, _09828_, _01275_);
  nor (_09830_, _01296_, _28330_);
  nor (_09831_, _01290_, _23530_);
  nor (_09832_, _09831_, _09830_);
  nand (_09833_, _09832_, _01204_);
  nor (_09834_, _01290_, _28047_);
  nor (_09835_, _01296_, _23516_);
  nor (_09836_, _09835_, _09834_);
  nand (_09837_, _09836_, _01206_);
  nand (_09838_, _09837_, _09833_);
  nand (_09839_, _09838_, _01260_);
  nor (_09840_, _01296_, _28018_);
  nor (_09841_, _01290_, _27990_);
  nor (_09842_, _09841_, _09840_);
  nand (_09844_, _09842_, _01204_);
  nor (_09845_, _01290_, _23545_);
  nor (_09846_, _01296_, _27962_);
  nor (_09847_, _09846_, _09845_);
  nand (_09848_, _09847_, _01206_);
  nand (_09849_, _09848_, _09844_);
  nand (_09850_, _09849_, _01262_);
  nand (_09851_, _09850_, _09839_);
  nand (_09852_, _09851_, _01274_);
  nand (_09853_, _09852_, _09829_);
  nand (_09854_, _09853_, _01241_);
  nand (_09855_, _09854_, _09807_);
  nand (_09856_, _09855_, _01244_);
  nand (_09857_, _09856_, _09758_);
  nor (_09858_, _09857_, _01231_);
  nand (_09859_, _01296_, _26259_);
  nand (_09860_, _01290_, _26287_);
  nand (_09861_, _09860_, _09859_);
  nand (_09862_, _09861_, _01204_);
  nand (_09863_, _01290_, _26230_);
  nand (_09864_, _01296_, _26202_);
  nand (_09865_, _09864_, _09863_);
  nand (_09866_, _09865_, _01206_);
  nand (_09867_, _09866_, _09862_);
  nand (_09868_, _09867_, _01260_);
  nand (_09869_, _01296_, _26145_);
  nand (_09870_, _01290_, _26174_);
  nand (_09871_, _09870_, _09869_);
  nand (_09872_, _09871_, _01204_);
  nand (_09873_, _01290_, _26117_);
  nand (_09874_, _01296_, _26089_);
  nand (_09875_, _09874_, _09873_);
  nand (_09876_, _09875_, _01206_);
  nand (_09877_, _09876_, _09872_);
  nand (_09878_, _09877_, _01262_);
  nand (_09879_, _09878_, _09868_);
  nand (_09880_, _09879_, _01275_);
  nor (_09881_, _01296_, _26004_);
  nor (_09882_, _01290_, _25975_);
  nor (_09883_, _09882_, _09881_);
  nand (_09885_, _09883_, _01206_);
  nand (_09886_, _01290_, _26060_);
  nand (_09887_, _01296_, _26032_);
  nand (_09888_, _09887_, _09886_);
  nand (_09889_, _09888_, _01204_);
  nand (_09890_, _09889_, _09885_);
  nand (_09891_, _09890_, _01260_);
  nor (_09892_, _01296_, _25889_);
  nor (_09893_, _01290_, _25861_);
  nor (_09894_, _09893_, _09892_);
  nand (_09895_, _09894_, _01206_);
  nand (_09896_, _01290_, _25947_);
  nand (_09897_, _01296_, _25919_);
  nand (_09898_, _09897_, _09896_);
  nand (_09899_, _09898_, _01204_);
  nand (_09900_, _09899_, _09895_);
  nand (_09901_, _09900_, _01262_);
  nand (_09902_, _09901_, _09891_);
  nand (_09903_, _09902_, _01274_);
  nand (_09904_, _09903_, _09880_);
  nand (_09905_, _09904_, _01308_);
  nand (_09906_, _01290_, _25832_);
  nand (_09907_, _01296_, _25804_);
  nand (_09908_, _09907_, _09906_);
  nand (_09909_, _09908_, _01204_);
  nand (_09910_, _01296_, _25747_);
  nand (_09911_, _01290_, _25776_);
  nand (_09912_, _09911_, _09910_);
  nand (_09913_, _09912_, _01206_);
  nand (_09914_, _09913_, _09909_);
  nand (_09915_, _09914_, _01260_);
  nand (_09916_, _01290_, _25719_);
  nand (_09917_, _01296_, _25691_);
  nand (_09918_, _09917_, _09916_);
  nand (_09919_, _09918_, _01204_);
  nand (_09920_, _01296_, _25634_);
  nand (_09921_, _01290_, _25662_);
  nand (_09922_, _09921_, _09920_);
  nand (_09923_, _09922_, _01206_);
  nand (_09924_, _09923_, _09919_);
  nand (_09926_, _09924_, _01262_);
  nand (_09927_, _09926_, _09915_);
  nand (_09928_, _09927_, _01275_);
  nor (_09929_, _01296_, _25606_);
  nor (_09930_, _01290_, _25582_);
  nor (_09931_, _09930_, _09929_);
  nand (_09932_, _09931_, _01204_);
  nor (_09933_, _01290_, _25554_);
  nor (_09934_, _01296_, _25568_);
  nor (_09935_, _09934_, _09933_);
  nand (_09936_, _09935_, _01206_);
  nand (_09937_, _09936_, _09932_);
  nand (_09938_, _09937_, _01260_);
  nor (_09939_, _01296_, _25539_);
  nor (_09940_, _01290_, _25525_);
  nor (_09941_, _09940_, _09939_);
  nand (_09942_, _09941_, _01204_);
  nor (_09943_, _01290_, _25496_);
  nor (_09944_, _01296_, _25511_);
  nor (_09945_, _09944_, _09943_);
  nand (_09946_, _09945_, _01206_);
  nand (_09947_, _09946_, _09942_);
  nand (_09948_, _09947_, _01262_);
  nand (_09949_, _09948_, _09938_);
  nand (_09950_, _09949_, _01274_);
  nand (_09951_, _09950_, _09928_);
  nand (_09952_, _09951_, _01241_);
  nand (_09953_, _09952_, _09905_);
  nand (_09954_, _09953_, _01245_);
  nor (_09955_, _01296_, _26400_);
  nor (_09956_, _01290_, _26372_);
  nor (_09957_, _09956_, _09955_);
  nand (_09958_, _09957_, _01204_);
  nor (_09959_, _01290_, _26315_);
  nor (_09960_, _01296_, _26344_);
  nor (_09961_, _09960_, _09959_);
  nand (_09962_, _09961_, _01206_);
  nand (_09963_, _09962_, _09958_);
  nand (_09964_, _09963_, _01262_);
  nor (_09965_, _01296_, _26514_);
  nor (_09967_, _01290_, _26486_);
  nor (_09968_, _09967_, _09965_);
  nand (_09969_, _09968_, _01204_);
  nor (_09970_, _01290_, _26429_);
  nor (_09971_, _01296_, _26457_);
  nor (_09972_, _09971_, _09970_);
  nand (_09973_, _09972_, _01206_);
  nand (_09974_, _09973_, _09969_);
  nand (_09975_, _09974_, _01260_);
  nand (_09976_, _09975_, _09964_);
  nand (_09977_, _09976_, _01274_);
  nand (_09978_, _01290_, _26627_);
  nand (_09979_, _01296_, _26599_);
  nand (_09980_, _09979_, _09978_);
  nand (_09981_, _09980_, _01204_);
  nand (_09982_, _01296_, _26542_);
  nand (_09983_, _01290_, _26571_);
  nand (_09984_, _09983_, _09982_);
  nand (_09985_, _09984_, _01206_);
  nand (_09986_, _09985_, _09981_);
  nand (_09987_, _09986_, _01262_);
  nand (_09988_, _01290_, _26742_);
  nand (_09989_, _01296_, _26712_);
  nand (_09990_, _09989_, _09988_);
  nand (_09991_, _09990_, _01204_);
  nand (_09992_, _01296_, _26656_);
  nand (_09993_, _01290_, _26684_);
  nand (_09994_, _09993_, _09992_);
  nand (_09995_, _09994_, _01206_);
  nand (_09996_, _09995_, _09991_);
  nand (_09997_, _09996_, _01260_);
  nand (_09998_, _09997_, _09987_);
  nand (_09999_, _09998_, _01275_);
  nand (_10000_, _09999_, _09977_);
  nand (_10001_, _10000_, _01241_);
  nor (_10002_, _01296_, _26798_);
  nor (_10003_, _01290_, _26770_);
  nor (_10004_, _10003_, _10002_);
  nand (_10005_, _10004_, _01206_);
  nand (_10006_, _01290_, _26855_);
  nand (_10008_, _01296_, _26827_);
  nand (_10009_, _10008_, _10006_);
  nand (_10010_, _10009_, _01204_);
  nand (_10011_, _10010_, _10005_);
  nand (_10012_, _10011_, _01262_);
  nor (_10013_, _01296_, _26912_);
  nor (_10014_, _01290_, _26883_);
  nor (_10015_, _10014_, _10013_);
  nand (_10016_, _10015_, _01206_);
  nand (_10017_, _01290_, _26968_);
  nand (_10018_, _01296_, _26940_);
  nand (_10019_, _10018_, _10017_);
  nand (_10020_, _10019_, _01204_);
  nand (_10021_, _10020_, _10016_);
  nand (_10022_, _10021_, _01260_);
  nand (_10023_, _10022_, _10012_);
  nand (_10024_, _10023_, _01274_);
  nand (_10025_, _01296_, _27054_);
  nand (_10026_, _01290_, _27082_);
  nand (_10027_, _10026_, _10025_);
  nand (_10028_, _10027_, _01204_);
  nand (_10029_, _01290_, _27025_);
  nand (_10030_, _01296_, _26997_);
  nand (_10031_, _10030_, _10029_);
  nand (_10032_, _10031_, _01206_);
  nand (_10033_, _10032_, _10028_);
  nand (_10034_, _10033_, _01262_);
  nand (_10035_, _01296_, _27167_);
  nand (_10036_, _01290_, _27195_);
  nand (_10037_, _10036_, _10035_);
  nand (_10038_, _10037_, _01204_);
  nand (_10039_, _01290_, _27139_);
  nand (_10040_, _01296_, _27110_);
  nand (_10041_, _10040_, _10039_);
  nand (_10042_, _10041_, _01206_);
  nand (_10043_, _10042_, _10038_);
  nand (_10044_, _10043_, _01260_);
  nand (_10045_, _10044_, _10034_);
  nand (_10046_, _10045_, _01275_);
  nand (_10047_, _10046_, _10024_);
  nand (_10049_, _10047_, _01308_);
  nand (_10050_, _10049_, _10001_);
  nand (_10051_, _10050_, _01244_);
  nand (_10052_, _10051_, _09954_);
  nor (_10053_, _10052_, _01235_);
  nor (_10054_, _10053_, _09858_);
  nor (_10055_, _10054_, _28717_);
  nand (_10056_, _01290_, _24848_);
  nand (_10057_, _01296_, _24834_);
  nand (_10058_, _10057_, _10056_);
  nand (_10059_, _10058_, _01204_);
  nand (_10060_, _01296_, _24805_);
  nand (_10061_, _01290_, _24820_);
  nand (_10062_, _10061_, _10060_);
  nand (_10063_, _10062_, _01206_);
  nand (_10064_, _10063_, _10059_);
  nand (_10065_, _10064_, _01260_);
  nand (_10066_, _01290_, _24791_);
  nand (_10067_, _01296_, _24777_);
  nand (_10068_, _10067_, _10066_);
  nand (_10069_, _10068_, _01204_);
  nand (_10070_, _01296_, _24748_);
  nand (_10071_, _01290_, _24762_);
  nand (_10072_, _10071_, _10070_);
  nand (_10073_, _10072_, _01206_);
  nand (_10074_, _10073_, _10069_);
  nand (_10075_, _10074_, _01262_);
  nand (_10076_, _10075_, _10065_);
  nand (_10077_, _10076_, _01275_);
  nor (_10078_, _01296_, _24734_);
  nor (_10079_, _01290_, _24719_);
  nor (_10080_, _10079_, _10078_);
  nand (_10081_, _10080_, _01204_);
  nor (_10082_, _01290_, _24691_);
  nor (_10083_, _01296_, _24705_);
  nor (_10084_, _10083_, _10082_);
  nand (_10085_, _10084_, _01206_);
  nand (_10086_, _10085_, _10081_);
  nand (_10087_, _10086_, _01260_);
  nor (_10088_, _01296_, _24676_);
  nor (_10090_, _01290_, _24662_);
  nor (_10091_, _10090_, _10088_);
  nand (_10092_, _10091_, _01204_);
  nor (_10093_, _01290_, _24633_);
  nor (_10094_, _01296_, _24648_);
  nor (_10095_, _10094_, _10093_);
  nand (_10096_, _10095_, _01206_);
  nand (_10097_, _10096_, _10092_);
  nand (_10098_, _10097_, _01262_);
  nand (_10099_, _10098_, _10087_);
  nand (_10100_, _10099_, _01274_);
  nand (_10101_, _10100_, _10077_);
  nand (_10102_, _10101_, _01241_);
  nand (_10103_, _01296_, _25065_);
  nand (_10104_, _01290_, _25079_);
  nand (_10105_, _10104_, _10103_);
  nand (_10106_, _10105_, _01204_);
  nand (_10107_, _01290_, _25050_);
  nand (_10108_, _01296_, _25036_);
  nand (_10109_, _10108_, _10107_);
  nand (_10110_, _10109_, _01206_);
  nand (_10111_, _10110_, _10106_);
  nand (_10112_, _10111_, _01260_);
  nand (_10113_, _01296_, _25007_);
  nand (_10114_, _01290_, _25022_);
  nand (_10115_, _10114_, _10113_);
  nand (_10116_, _10115_, _01204_);
  nand (_10117_, _01290_, _24993_);
  nand (_10118_, _01296_, _24979_);
  nand (_10119_, _10118_, _10117_);
  nand (_10120_, _10119_, _01206_);
  nand (_10121_, _10120_, _10116_);
  nand (_10122_, _10121_, _01262_);
  nand (_10123_, _10122_, _10112_);
  nand (_10124_, _10123_, _01275_);
  nor (_10125_, _01296_, _24936_);
  nor (_10126_, _01290_, _24920_);
  nor (_10127_, _10126_, _10125_);
  nand (_10128_, _10127_, _01206_);
  nand (_10129_, _01290_, _24964_);
  nand (_10131_, _01296_, _24950_);
  nand (_10132_, _10131_, _10129_);
  nand (_10133_, _10132_, _01204_);
  nand (_10134_, _10133_, _10128_);
  nand (_10135_, _10134_, _01260_);
  nor (_10136_, _01296_, _24877_);
  nor (_10137_, _01290_, _24863_);
  nor (_10138_, _10137_, _10136_);
  nand (_10139_, _10138_, _01206_);
  nand (_10140_, _01290_, _24906_);
  nand (_10141_, _01296_, _24892_);
  nand (_10142_, _10141_, _10140_);
  nand (_10143_, _10142_, _01204_);
  nand (_10144_, _10143_, _10139_);
  nand (_10145_, _10144_, _01262_);
  nand (_10146_, _10145_, _10135_);
  nand (_10147_, _10146_, _01274_);
  nand (_10148_, _10147_, _10124_);
  nand (_10149_, _10148_, _01308_);
  nand (_10150_, _10149_, _10102_);
  nand (_10151_, _10150_, _01245_);
  nand (_10152_, _01296_, _25468_);
  nand (_10153_, _01290_, _25482_);
  nand (_10154_, _10153_, _10152_);
  nand (_10155_, _10154_, _01204_);
  nand (_10156_, _01290_, _25453_);
  nand (_10157_, _01296_, _25439_);
  nand (_10158_, _10157_, _10156_);
  nand (_10159_, _10158_, _01206_);
  nand (_10160_, _10159_, _10155_);
  nand (_10161_, _10160_, _01260_);
  nand (_10162_, _01296_, _25410_);
  nand (_10163_, _01290_, _25424_);
  nand (_10164_, _10163_, _10162_);
  nand (_10165_, _10164_, _01204_);
  nand (_10166_, _01290_, _25396_);
  nand (_10167_, _01296_, _25381_);
  nand (_10168_, _10167_, _10166_);
  nand (_10169_, _10168_, _01206_);
  nand (_10170_, _10169_, _10165_);
  nand (_10172_, _10170_, _01262_);
  nand (_10173_, _10172_, _10161_);
  nand (_10174_, _10173_, _01275_);
  nor (_10175_, _01296_, _25337_);
  nor (_10176_, _01290_, _25323_);
  nor (_10177_, _10176_, _10175_);
  nand (_10178_, _10177_, _01206_);
  nand (_10179_, _01290_, _25367_);
  nand (_10180_, _01296_, _25353_);
  nand (_10181_, _10180_, _10179_);
  nand (_10182_, _10181_, _01204_);
  nand (_10183_, _10182_, _10178_);
  nand (_10184_, _10183_, _01260_);
  nor (_10185_, _01296_, _25280_);
  nor (_10186_, _01290_, _25266_);
  nor (_10187_, _10186_, _10185_);
  nand (_10188_, _10187_, _01206_);
  nand (_10189_, _01290_, _25309_);
  nand (_10190_, _01296_, _25294_);
  nand (_10191_, _10190_, _10189_);
  nand (_10192_, _10191_, _01204_);
  nand (_10193_, _10192_, _10188_);
  nand (_10194_, _10193_, _01262_);
  nand (_10195_, _10194_, _10184_);
  nand (_10196_, _10195_, _01274_);
  nand (_10197_, _10196_, _10174_);
  nand (_10198_, _10197_, _01308_);
  nand (_10199_, _01290_, _25251_);
  nand (_10200_, _01296_, _25237_);
  nand (_10201_, _10200_, _10199_);
  nand (_10202_, _10201_, _01204_);
  nand (_10203_, _01296_, _25208_);
  nand (_10204_, _01290_, _25223_);
  nand (_10205_, _10204_, _10203_);
  nand (_10206_, _10205_, _01206_);
  nand (_10207_, _10206_, _10202_);
  nand (_10208_, _10207_, _01260_);
  nand (_10209_, _01290_, _25194_);
  nand (_10210_, _01296_, _25180_);
  nand (_10211_, _10210_, _10209_);
  nand (_10214_, _10211_, _01204_);
  nand (_10215_, _01296_, _25151_);
  nand (_10216_, _01290_, _25165_);
  nand (_10217_, _10216_, _10215_);
  nand (_10218_, _10217_, _01206_);
  nand (_10220_, _10218_, _10214_);
  nand (_10221_, _10220_, _01262_);
  nand (_10222_, _10221_, _10208_);
  nand (_10223_, _10222_, _01275_);
  nor (_10224_, _01296_, _25136_);
  nor (_10225_, _01290_, _25122_);
  nor (_10226_, _10225_, _10224_);
  nand (_10227_, _10226_, _01204_);
  nor (_10228_, _01290_, _23674_);
  nor (_10229_, _01296_, _25108_);
  nor (_10230_, _10229_, _10228_);
  nand (_10231_, _10230_, _01206_);
  nand (_10232_, _10231_, _10227_);
  nand (_10233_, _10232_, _01260_);
  nor (_10234_, _01296_, _23645_);
  nor (_10235_, _01290_, _23631_);
  nor (_10236_, _10235_, _10234_);
  nand (_10237_, _10236_, _01204_);
  nor (_10238_, _01290_, _25093_);
  nor (_10239_, _01296_, _23659_);
  nor (_10240_, _10239_, _10238_);
  nand (_10241_, _10240_, _01206_);
  nand (_10242_, _10241_, _10237_);
  nand (_10243_, _10242_, _01262_);
  nand (_10244_, _10243_, _10233_);
  nand (_10245_, _10244_, _01274_);
  nand (_10246_, _10245_, _10223_);
  nand (_10247_, _10246_, _01241_);
  nand (_10248_, _10247_, _10198_);
  nand (_10249_, _10248_, _01244_);
  nand (_10250_, _10249_, _10151_);
  nor (_10251_, _10250_, _01231_);
  nand (_10252_, _01296_, _24144_);
  nand (_10253_, _01290_, _24159_);
  nand (_10254_, _10253_, _10252_);
  nand (_10256_, _10254_, _01204_);
  nand (_10257_, _01290_, _24130_);
  nand (_10259_, _01296_, _24116_);
  nand (_10260_, _10259_, _10257_);
  nand (_10261_, _10260_, _01206_);
  nand (_10262_, _10261_, _10256_);
  nand (_10263_, _10262_, _01260_);
  nand (_10264_, _01296_, _24086_);
  nand (_10265_, _01290_, _24100_);
  nand (_10266_, _10265_, _10264_);
  nand (_10267_, _10266_, _01204_);
  nand (_10268_, _01290_, _24072_);
  nand (_10269_, _01296_, _24057_);
  nand (_10270_, _10269_, _10268_);
  nand (_10271_, _10270_, _01206_);
  nand (_10273_, _10271_, _10267_);
  nand (_10274_, _10273_, _01262_);
  nand (_10275_, _10274_, _10263_);
  nand (_10276_, _10275_, _01275_);
  nor (_10277_, _01296_, _24014_);
  nor (_10278_, _01290_, _24000_);
  nor (_10279_, _10278_, _10277_);
  nand (_10280_, _10279_, _01206_);
  nand (_10281_, _01290_, _24043_);
  nand (_10282_, _01296_, _24029_);
  nand (_10283_, _10282_, _10281_);
  nand (_10284_, _10283_, _01204_);
  nand (_10285_, _10284_, _10280_);
  nand (_10286_, _10285_, _01260_);
  nor (_10287_, _01296_, _23957_);
  nor (_10288_, _01290_, _23942_);
  nor (_10289_, _10288_, _10287_);
  nand (_10290_, _10289_, _01206_);
  nand (_10291_, _01290_, _23985_);
  nand (_10292_, _01296_, _23971_);
  nand (_10293_, _10292_, _10291_);
  nand (_10294_, _10293_, _01204_);
  nand (_10295_, _10294_, _10290_);
  nand (_10296_, _10295_, _01262_);
  nand (_10297_, _10296_, _10286_);
  nand (_10299_, _10297_, _01274_);
  nand (_10300_, _10299_, _10276_);
  nand (_10301_, _10300_, _01308_);
  nand (_10302_, _01290_, _23928_);
  nand (_10303_, _01296_, _23914_);
  nand (_10304_, _10303_, _10302_);
  nand (_10305_, _10304_, _01204_);
  nand (_10306_, _01296_, _23885_);
  nand (_10307_, _01290_, _23899_);
  nand (_10308_, _10307_, _10306_);
  nand (_10309_, _10308_, _01206_);
  nand (_10310_, _10309_, _10305_);
  nand (_10311_, _10310_, _01260_);
  nand (_10312_, _01290_, _23871_);
  nand (_10313_, _01296_, _23856_);
  nand (_10314_, _10313_, _10312_);
  nand (_10315_, _10314_, _01204_);
  nand (_10316_, _01296_, _23828_);
  nand (_10317_, _01290_, _23842_);
  nand (_10318_, _10317_, _10316_);
  nand (_10319_, _10318_, _01206_);
  nand (_10320_, _10319_, _10315_);
  nand (_10321_, _10320_, _01262_);
  nand (_10322_, _10321_, _10311_);
  nand (_10323_, _10322_, _01275_);
  nor (_10324_, _01296_, _23813_);
  nor (_10325_, _01290_, _23799_);
  nor (_10326_, _10325_, _10324_);
  nand (_10327_, _10326_, _01204_);
  nor (_10328_, _01290_, _23770_);
  nor (_10329_, _01296_, _23785_);
  nor (_10330_, _10329_, _10328_);
  nand (_10331_, _10330_, _01206_);
  nand (_10332_, _10331_, _10327_);
  nand (_10333_, _10332_, _01260_);
  nor (_10334_, _01296_, _23756_);
  nor (_10335_, _01290_, _23742_);
  nor (_10336_, _10335_, _10334_);
  nand (_10337_, _10336_, _01204_);
  nor (_10338_, _01290_, _23713_);
  nor (_10340_, _01296_, _23727_);
  nor (_10341_, _10340_, _10338_);
  nand (_10342_, _10341_, _01206_);
  nand (_10343_, _10342_, _10337_);
  nand (_10344_, _10343_, _01262_);
  nand (_10345_, _10344_, _10333_);
  nand (_10346_, _10345_, _01274_);
  nand (_10347_, _10346_, _10323_);
  nand (_10348_, _10347_, _01241_);
  nand (_10349_, _10348_, _10301_);
  nand (_10350_, _10349_, _01245_);
  nor (_10351_, _01296_, _24216_);
  nor (_10352_, _01290_, _24202_);
  nor (_10353_, _10352_, _10351_);
  nand (_10354_, _10353_, _01204_);
  nor (_10355_, _01290_, _24173_);
  nor (_10356_, _01296_, _24187_);
  nor (_10357_, _10356_, _10355_);
  nand (_10358_, _10357_, _01206_);
  nand (_10359_, _10358_, _10354_);
  nand (_10360_, _10359_, _01262_);
  nor (_10361_, _01296_, _24273_);
  nor (_10362_, _01290_, _24259_);
  nor (_10363_, _10362_, _10361_);
  nand (_10364_, _10363_, _01204_);
  nor (_10365_, _01290_, _24230_);
  nor (_10366_, _01296_, _24245_);
  nor (_10367_, _10366_, _10365_);
  nand (_10368_, _10367_, _01206_);
  nand (_10369_, _10368_, _10364_);
  nand (_10370_, _10369_, _01260_);
  nand (_10371_, _10370_, _10360_);
  nand (_10372_, _10371_, _01274_);
  nand (_10373_, _01290_, _24331_);
  nand (_10374_, _01296_, _24317_);
  nand (_10375_, _10374_, _10373_);
  nand (_10376_, _10375_, _01204_);
  nand (_10377_, _01296_, _24288_);
  nand (_10378_, _01290_, _24302_);
  nand (_10379_, _10378_, _10377_);
  nand (_10381_, _10379_, _01206_);
  nand (_10382_, _10381_, _10376_);
  nand (_10383_, _10382_, _01262_);
  nand (_10384_, _01290_, _24388_);
  nand (_10385_, _01296_, _24374_);
  nand (_10386_, _10385_, _10384_);
  nand (_10387_, _10386_, _01204_);
  nand (_10388_, _01296_, _24345_);
  nand (_10389_, _01290_, _24360_);
  nand (_10390_, _10389_, _10388_);
  nand (_10391_, _10390_, _01206_);
  nand (_10392_, _10391_, _10387_);
  nand (_10393_, _10392_, _01260_);
  nand (_10394_, _10393_, _10383_);
  nand (_10395_, _10394_, _01275_);
  nand (_10396_, _10395_, _10372_);
  nand (_10397_, _10396_, _01241_);
  nor (_10398_, _01296_, _24417_);
  nor (_10399_, _01290_, _24403_);
  nor (_10400_, _10399_, _10398_);
  nand (_10401_, _10400_, _01206_);
  nand (_10402_, _01290_, _24446_);
  nand (_10403_, _01296_, _24431_);
  nand (_10404_, _10403_, _10402_);
  nand (_10405_, _10404_, _01204_);
  nand (_10406_, _10405_, _10401_);
  nand (_10407_, _10406_, _01262_);
  nor (_10408_, _01296_, _24474_);
  nor (_10409_, _01290_, _24460_);
  nor (_10410_, _10409_, _10408_);
  nand (_10411_, _10410_, _01206_);
  nand (_10412_, _01290_, _24503_);
  nand (_10413_, _01296_, _24489_);
  nand (_10414_, _10413_, _10412_);
  nand (_10415_, _10414_, _01204_);
  nand (_10416_, _10415_, _10411_);
  nand (_10417_, _10416_, _01260_);
  nand (_10418_, _10417_, _10407_);
  nand (_10419_, _10418_, _01274_);
  nand (_10420_, _01296_, _24547_);
  nand (_10422_, _01290_, _24561_);
  nand (_10423_, _10422_, _10420_);
  nand (_10424_, _10423_, _01204_);
  nand (_10425_, _01290_, _24533_);
  nand (_10426_, _01296_, _24517_);
  nand (_10427_, _10426_, _10425_);
  nand (_10428_, _10427_, _01206_);
  nand (_10429_, _10428_, _10424_);
  nand (_10430_, _10429_, _01262_);
  nand (_10431_, _01296_, _24605_);
  nand (_10432_, _01290_, _24619_);
  nand (_10433_, _10432_, _10431_);
  nand (_10434_, _10433_, _01204_);
  nand (_10435_, _01290_, _24590_);
  nand (_10436_, _01296_, _24576_);
  nand (_10437_, _10436_, _10435_);
  nand (_10438_, _10437_, _01206_);
  nand (_10439_, _10438_, _10434_);
  nand (_10440_, _10439_, _01260_);
  nand (_10441_, _10440_, _10430_);
  nand (_10442_, _10441_, _01275_);
  nand (_10443_, _10442_, _10419_);
  nand (_10444_, _10443_, _01308_);
  nand (_10445_, _10444_, _10397_);
  nand (_10446_, _10445_, _01244_);
  nand (_10447_, _10446_, _10350_);
  nor (_10448_, _10447_, _01235_);
  nor (_10449_, _10448_, _10251_);
  nor (_10450_, _10449_, _28718_);
  nor (_10451_, _10450_, _10055_);
  nor (_10452_, _10451_, _06280_);
  nand (_10453_, _06280_, _28511_);
  nand (_10454_, _10453_, _29344_);
  nor (_15161_, _10454_, _10452_);
  nand (_10455_, _01290_, _27569_);
  nand (_10456_, _01296_, _27541_);
  nand (_10457_, _10456_, _10455_);
  nand (_10458_, _10457_, _01204_);
  nand (_10459_, _01296_, _23604_);
  nand (_10460_, _01290_, _27511_);
  nand (_10462_, _10460_, _10459_);
  nand (_10463_, _10462_, _01206_);
  nand (_10464_, _10463_, _10458_);
  nand (_10465_, _10464_, _01260_);
  nand (_10466_, _01290_, _23701_);
  nand (_10467_, _01296_, _23618_);
  nand (_10468_, _10467_, _10466_);
  nand (_10469_, _10468_, _01204_);
  nand (_10470_, _01296_, _27454_);
  nand (_10471_, _01290_, _27483_);
  nand (_10472_, _10471_, _10470_);
  nand (_10473_, _10472_, _01206_);
  nand (_10474_, _10473_, _10469_);
  nand (_10475_, _10474_, _01262_);
  nand (_10476_, _10475_, _10465_);
  nand (_10477_, _10476_, _01275_);
  nor (_10478_, _01296_, _27426_);
  nor (_10479_, _01290_, _27398_);
  nor (_10480_, _10479_, _10478_);
  nand (_10481_, _10480_, _01204_);
  nor (_10482_, _01290_, _27341_);
  nor (_10483_, _01296_, _27369_);
  nor (_10484_, _10483_, _10482_);
  nand (_10485_, _10484_, _01206_);
  nand (_10486_, _10485_, _10481_);
  nand (_10487_, _10486_, _01260_);
  nor (_10488_, _01296_, _27313_);
  nor (_10489_, _01290_, _27284_);
  nor (_10490_, _10489_, _10488_);
  nand (_10491_, _10490_, _01204_);
  nor (_10492_, _01290_, _27228_);
  nor (_10493_, _01296_, _27256_);
  nor (_10494_, _10493_, _10492_);
  nand (_10495_, _10494_, _01206_);
  nand (_10496_, _10495_, _10491_);
  nand (_10497_, _10496_, _01262_);
  nand (_10498_, _10497_, _10487_);
  nand (_10499_, _10498_, _01274_);
  nand (_10500_, _10499_, _10477_);
  nand (_10501_, _10500_, _01241_);
  nand (_10503_, _01296_, _23561_);
  nand (_10504_, _01290_, _27937_);
  nand (_10505_, _10504_, _10503_);
  nand (_10506_, _10505_, _01204_);
  nand (_10507_, _01290_, _27909_);
  nand (_10508_, _01296_, _23575_);
  nand (_10509_, _10508_, _10507_);
  nand (_10510_, _10509_, _01206_);
  nand (_10511_, _10510_, _10506_);
  nand (_10512_, _10511_, _01260_);
  nand (_10513_, _01296_, _27852_);
  nand (_10514_, _01290_, _27881_);
  nand (_10515_, _10514_, _10513_);
  nand (_10516_, _10515_, _01204_);
  nand (_10517_, _01290_, _27824_);
  nand (_10518_, _01296_, _27796_);
  nand (_10519_, _10518_, _10517_);
  nand (_10520_, _10519_, _01206_);
  nand (_10521_, _10520_, _10516_);
  nand (_10522_, _10521_, _01262_);
  nand (_10523_, _10522_, _10512_);
  nand (_10524_, _10523_, _01275_);
  nor (_10525_, _01296_, _27711_);
  nor (_10526_, _01290_, _27682_);
  nor (_10527_, _10526_, _10525_);
  nand (_10528_, _10527_, _01206_);
  nand (_10529_, _01290_, _27767_);
  nand (_10530_, _01296_, _27739_);
  nand (_10531_, _10530_, _10529_);
  nand (_10532_, _10531_, _01204_);
  nand (_10533_, _10532_, _10528_);
  nand (_10534_, _10533_, _01260_);
  nor (_10535_, _01296_, _27626_);
  nor (_10536_, _01290_, _27597_);
  nor (_10537_, _10536_, _10535_);
  nand (_10538_, _10537_, _01206_);
  nand (_10539_, _01290_, _23590_);
  nand (_10540_, _01296_, _27654_);
  nand (_10541_, _10540_, _10539_);
  nand (_10542_, _10541_, _01204_);
  nand (_10544_, _10542_, _10538_);
  nand (_10545_, _10544_, _01262_);
  nand (_10546_, _10545_, _10534_);
  nand (_10547_, _10546_, _01274_);
  nand (_10548_, _10547_, _10524_);
  nand (_10549_, _10548_, _01308_);
  nand (_10550_, _10549_, _10501_);
  nand (_10551_, _10550_, _01245_);
  nand (_10552_, _01296_, _28392_);
  nand (_10553_, _01290_, _28420_);
  nand (_10554_, _10553_, _10552_);
  nand (_10555_, _10554_, _01204_);
  nand (_10556_, _01290_, _28364_);
  nand (_10557_, _01296_, _28306_);
  nand (_10558_, _10557_, _10556_);
  nand (_10559_, _10558_, _01206_);
  nand (_10560_, _10559_, _10555_);
  nand (_10561_, _10560_, _01260_);
  nand (_10562_, _01296_, _28249_);
  nand (_10563_, _01290_, _28278_);
  nand (_10564_, _10563_, _10562_);
  nand (_10565_, _10564_, _01204_);
  nand (_10566_, _01290_, _28193_);
  nand (_10567_, _01296_, _28164_);
  nand (_10568_, _10567_, _10566_);
  nand (_10569_, _10568_, _01206_);
  nand (_10570_, _10569_, _10565_);
  nand (_10571_, _10570_, _01262_);
  nand (_10572_, _10571_, _10561_);
  nand (_10573_, _10572_, _01275_);
  nor (_10574_, _01296_, _28079_);
  nor (_10575_, _01290_, _23504_);
  nor (_10576_, _10575_, _10574_);
  nand (_10577_, _10576_, _01206_);
  nand (_10578_, _01290_, _28136_);
  nand (_10579_, _01296_, _28108_);
  nand (_10580_, _10579_, _10578_);
  nand (_10581_, _10580_, _01204_);
  nand (_10582_, _10581_, _10577_);
  nand (_10583_, _10582_, _01260_);
  nor (_10585_, _01296_, _23461_);
  nor (_10586_, _01290_, _23446_);
  nor (_10587_, _10586_, _10585_);
  nand (_10588_, _10587_, _01206_);
  nand (_10589_, _01290_, _23489_);
  nand (_10590_, _01296_, _23475_);
  nand (_10591_, _10590_, _10589_);
  nand (_10592_, _10591_, _01204_);
  nand (_10593_, _10592_, _10588_);
  nand (_10594_, _10593_, _01262_);
  nand (_10595_, _10594_, _10583_);
  nand (_10596_, _10595_, _01274_);
  nand (_10597_, _10596_, _10573_);
  nand (_10598_, _10597_, _01308_);
  nand (_10599_, _01290_, _23432_);
  nand (_10600_, _01296_, _23418_);
  nand (_10601_, _10600_, _10599_);
  nand (_10602_, _10601_, _01204_);
  nand (_10603_, _01296_, _23389_);
  nand (_10604_, _01290_, _23403_);
  nand (_10605_, _10604_, _10603_);
  nand (_10606_, _10605_, _01206_);
  nand (_10607_, _10606_, _10602_);
  nand (_10608_, _10607_, _01260_);
  nand (_10609_, _01290_, _23374_);
  nand (_10610_, _01296_, _23360_);
  nand (_10611_, _10610_, _10609_);
  nand (_10612_, _10611_, _01204_);
  nand (_10613_, _01296_, _28221_);
  nand (_10614_, _01290_, _28445_);
  nand (_10615_, _10614_, _10613_);
  nand (_10616_, _10615_, _01206_);
  nand (_10617_, _10616_, _10612_);
  nand (_10618_, _10617_, _01262_);
  nand (_10619_, _10618_, _10608_);
  nand (_10620_, _10619_, _01275_);
  nor (_10621_, _01296_, _28334_);
  nor (_10622_, _01290_, _23532_);
  nor (_10623_, _10622_, _10621_);
  nand (_10624_, _10623_, _01204_);
  nor (_10629_, _01290_, _28051_);
  nor (_10630_, _01296_, _23518_);
  nor (_10631_, _10630_, _10629_);
  nand (_10632_, _10631_, _01206_);
  nand (_10633_, _10632_, _10624_);
  nand (_10634_, _10633_, _01260_);
  nor (_10635_, _01296_, _28022_);
  nor (_10636_, _01290_, _27994_);
  nor (_10637_, _10636_, _10635_);
  nand (_10638_, _10637_, _01204_);
  nor (_10639_, _01290_, _23547_);
  nor (_10640_, _01296_, _27966_);
  nor (_10641_, _10640_, _10639_);
  nand (_10642_, _10641_, _01206_);
  nand (_10643_, _10642_, _10638_);
  nand (_10644_, _10643_, _01262_);
  nand (_10645_, _10644_, _10634_);
  nand (_10646_, _10645_, _01274_);
  nand (_10647_, _10646_, _10620_);
  nand (_10648_, _10647_, _01241_);
  nand (_10649_, _10648_, _10598_);
  nand (_10650_, _10649_, _01244_);
  nand (_10651_, _10650_, _10551_);
  nor (_10652_, _10651_, _01231_);
  nand (_10653_, _01296_, _26263_);
  nand (_10654_, _01290_, _26291_);
  nand (_10655_, _10654_, _10653_);
  nand (_10656_, _10655_, _01204_);
  nand (_10657_, _01290_, _26234_);
  nand (_10658_, _01296_, _26206_);
  nand (_10659_, _10658_, _10657_);
  nand (_10660_, _10659_, _01206_);
  nand (_10661_, _10660_, _10656_);
  nand (_10662_, _10661_, _01260_);
  nand (_10663_, _01296_, _26149_);
  nand (_10664_, _01290_, _26178_);
  nand (_10665_, _10664_, _10663_);
  nand (_10666_, _10665_, _01204_);
  nand (_10667_, _01290_, _26121_);
  nand (_10668_, _01296_, _26093_);
  nand (_10670_, _10668_, _10667_);
  nand (_10671_, _10670_, _01206_);
  nand (_10672_, _10671_, _10666_);
  nand (_10673_, _10672_, _01262_);
  nand (_10674_, _10673_, _10662_);
  nand (_10675_, _10674_, _01275_);
  nor (_10676_, _01296_, _26008_);
  nor (_10677_, _01290_, _25979_);
  nor (_10678_, _10677_, _10676_);
  nand (_10679_, _10678_, _01206_);
  nand (_10680_, _01290_, _26064_);
  nand (_10681_, _01296_, _26036_);
  nand (_10682_, _10681_, _10680_);
  nand (_10683_, _10682_, _01204_);
  nand (_10684_, _10683_, _10679_);
  nand (_10685_, _10684_, _01260_);
  nor (_10686_, _01296_, _25893_);
  nor (_10687_, _01290_, _25865_);
  nor (_10688_, _10687_, _10686_);
  nand (_10689_, _10688_, _01206_);
  nand (_10690_, _01290_, _25951_);
  nand (_10691_, _01296_, _25923_);
  nand (_10692_, _10691_, _10690_);
  nand (_10693_, _10692_, _01204_);
  nand (_10694_, _10693_, _10689_);
  nand (_10695_, _10694_, _01262_);
  nand (_10696_, _10695_, _10685_);
  nand (_10697_, _10696_, _01274_);
  nand (_10698_, _10697_, _10675_);
  nand (_10699_, _10698_, _01308_);
  nand (_10700_, _01290_, _25837_);
  nand (_10701_, _01296_, _25808_);
  nand (_10702_, _10701_, _10700_);
  nand (_10703_, _10702_, _01204_);
  nand (_10704_, _01296_, _25751_);
  nand (_10705_, _01290_, _25780_);
  nand (_10706_, _10705_, _10704_);
  nand (_10707_, _10706_, _01206_);
  nand (_10708_, _10707_, _10703_);
  nand (_10709_, _10708_, _01260_);
  nand (_10711_, _01290_, _25723_);
  nand (_10712_, _01296_, _25695_);
  nand (_10713_, _10712_, _10711_);
  nand (_10714_, _10713_, _01204_);
  nand (_10715_, _01296_, _25638_);
  nand (_10716_, _01290_, _25666_);
  nand (_10717_, _10716_, _10715_);
  nand (_10718_, _10717_, _01206_);
  nand (_10719_, _10718_, _10714_);
  nand (_10720_, _10719_, _01262_);
  nand (_10721_, _10720_, _10709_);
  nand (_10722_, _10721_, _01275_);
  nor (_10723_, _01296_, _25610_);
  nor (_10724_, _01290_, _25584_);
  nor (_10725_, _10724_, _10723_);
  nand (_10726_, _10725_, _01204_);
  nor (_10727_, _01290_, _25556_);
  nor (_10728_, _01296_, _25570_);
  nor (_10729_, _10728_, _10727_);
  nand (_10730_, _10729_, _01206_);
  nand (_10731_, _10730_, _10726_);
  nand (_10732_, _10731_, _01260_);
  nor (_10733_, _01296_, _25541_);
  nor (_10734_, _01290_, _25527_);
  nor (_10735_, _10734_, _10733_);
  nand (_10736_, _10735_, _01204_);
  nor (_10737_, _01290_, _25498_);
  nor (_10738_, _01296_, _25513_);
  nor (_10739_, _10738_, _10737_);
  nand (_10740_, _10739_, _01206_);
  nand (_10741_, _10740_, _10736_);
  nand (_10742_, _10741_, _01262_);
  nand (_10743_, _10742_, _10732_);
  nand (_10744_, _10743_, _01274_);
  nand (_10745_, _10744_, _10722_);
  nand (_10746_, _10745_, _01241_);
  nand (_10747_, _10746_, _10699_);
  nand (_10748_, _10747_, _01245_);
  nor (_10749_, _01296_, _26405_);
  nor (_10750_, _01290_, _26376_);
  nor (_10752_, _10750_, _10749_);
  nand (_10753_, _10752_, _01204_);
  nor (_10754_, _01290_, _26319_);
  nor (_10755_, _01296_, _26348_);
  nor (_10756_, _10755_, _10754_);
  nand (_10757_, _10756_, _01206_);
  nand (_10758_, _10757_, _10753_);
  nand (_10759_, _10758_, _01262_);
  nor (_10760_, _01296_, _26518_);
  nor (_10761_, _01290_, _26490_);
  nor (_10763_, _10761_, _10760_);
  nand (_10764_, _10763_, _01204_);
  nor (_10765_, _01290_, _26433_);
  nor (_10766_, _01296_, _26461_);
  nor (_10767_, _10766_, _10765_);
  nand (_10768_, _10767_, _01206_);
  nand (_10769_, _10768_, _10764_);
  nand (_10770_, _10769_, _01260_);
  nand (_10771_, _10770_, _10759_);
  nand (_10772_, _10771_, _01274_);
  nand (_10773_, _01290_, _26631_);
  nand (_10774_, _01296_, _26603_);
  nand (_10775_, _10774_, _10773_);
  nand (_10776_, _10775_, _01204_);
  nand (_10777_, _01296_, _26546_);
  nand (_10778_, _01290_, _26575_);
  nand (_10779_, _10778_, _10777_);
  nand (_10780_, _10779_, _01206_);
  nand (_10781_, _10780_, _10776_);
  nand (_10782_, _10781_, _01262_);
  nand (_10783_, _01290_, _26746_);
  nand (_10784_, _01296_, _26716_);
  nand (_10785_, _10784_, _10783_);
  nand (_10786_, _10785_, _01204_);
  nand (_10787_, _01296_, _26660_);
  nand (_10788_, _01290_, _26688_);
  nand (_10789_, _10788_, _10787_);
  nand (_10790_, _10789_, _01206_);
  nand (_10791_, _10790_, _10786_);
  nand (_10792_, _10791_, _01260_);
  nand (_10794_, _10792_, _10782_);
  nand (_10795_, _10794_, _01275_);
  nand (_10796_, _10795_, _10772_);
  nand (_10797_, _10796_, _01241_);
  nor (_10798_, _01296_, _26802_);
  nor (_10799_, _01290_, _26774_);
  nor (_10800_, _10799_, _10798_);
  nand (_10801_, _10800_, _01206_);
  nand (_10802_, _01290_, _26859_);
  nand (_10803_, _01296_, _26831_);
  nand (_10804_, _10803_, _10802_);
  nand (_10805_, _10804_, _01204_);
  nand (_10806_, _10805_, _10801_);
  nand (_10807_, _10806_, _01262_);
  nor (_10808_, _01296_, _26916_);
  nor (_10809_, _01290_, _26887_);
  nor (_10810_, _10809_, _10808_);
  nand (_10811_, _10810_, _01206_);
  nand (_10812_, _01290_, _26973_);
  nand (_10813_, _01296_, _26944_);
  nand (_10814_, _10813_, _10812_);
  nand (_10815_, _10814_, _01204_);
  nand (_10816_, _10815_, _10811_);
  nand (_10817_, _10816_, _01260_);
  nand (_10818_, _10817_, _10807_);
  nand (_10819_, _10818_, _01274_);
  nand (_10820_, _01296_, _27058_);
  nand (_10821_, _01290_, _27086_);
  nand (_10822_, _10821_, _10820_);
  nand (_10823_, _10822_, _01204_);
  nand (_10824_, _01290_, _27029_);
  nand (_10825_, _01296_, _27001_);
  nand (_10826_, _10825_, _10824_);
  nand (_10827_, _10826_, _01206_);
  nand (_10828_, _10827_, _10823_);
  nand (_10829_, _10828_, _01262_);
  nand (_10830_, _01296_, _27171_);
  nand (_10831_, _01290_, _27199_);
  nand (_10832_, _10831_, _10830_);
  nand (_10833_, _10832_, _01204_);
  nand (_10835_, _01290_, _27143_);
  nand (_10836_, _01296_, _27114_);
  nand (_10837_, _10836_, _10835_);
  nand (_10838_, _10837_, _01206_);
  nand (_10839_, _10838_, _10833_);
  nand (_10840_, _10839_, _01260_);
  nand (_10841_, _10840_, _10829_);
  nand (_10842_, _10841_, _01275_);
  nand (_10843_, _10842_, _10819_);
  nand (_10844_, _10843_, _01308_);
  nand (_10845_, _10844_, _10797_);
  nand (_10846_, _10845_, _01244_);
  nand (_10847_, _10846_, _10748_);
  nor (_10848_, _10847_, _01235_);
  nor (_10849_, _10848_, _10652_);
  nor (_10850_, _10849_, _28717_);
  nand (_10851_, _01290_, _24851_);
  nand (_10852_, _01296_, _24836_);
  nand (_10853_, _10852_, _10851_);
  nand (_10854_, _10853_, _01204_);
  nand (_10855_, _01296_, _24807_);
  nand (_10856_, _01290_, _24822_);
  nand (_10857_, _10856_, _10855_);
  nand (_10858_, _10857_, _01206_);
  nand (_10859_, _10858_, _10854_);
  nand (_10860_, _10859_, _01260_);
  nand (_10861_, _01290_, _24793_);
  nand (_10862_, _01296_, _24779_);
  nand (_10863_, _10862_, _10861_);
  nand (_10864_, _10863_, _01204_);
  nand (_10865_, _01296_, _24750_);
  nand (_10866_, _01290_, _24764_);
  nand (_10867_, _10866_, _10865_);
  nand (_10868_, _10867_, _01206_);
  nand (_10869_, _10868_, _10864_);
  nand (_10870_, _10869_, _01262_);
  nand (_10871_, _10870_, _10860_);
  nand (_10872_, _10871_, _01275_);
  nor (_10873_, _01296_, _24736_);
  nor (_10874_, _01290_, _24721_);
  nor (_10876_, _10874_, _10873_);
  nand (_10877_, _10876_, _01204_);
  nor (_10878_, _01290_, _24693_);
  nor (_10879_, _01296_, _24707_);
  nor (_10880_, _10879_, _10878_);
  nand (_10881_, _10880_, _01206_);
  nand (_10882_, _10881_, _10877_);
  nand (_10883_, _10882_, _01260_);
  nor (_10884_, _01296_, _24678_);
  nor (_10885_, _01290_, _24664_);
  nor (_10886_, _10885_, _10884_);
  nand (_10887_, _10886_, _01204_);
  nor (_10888_, _01290_, _24635_);
  nor (_10889_, _01296_, _24650_);
  nor (_10890_, _10889_, _10888_);
  nand (_10891_, _10890_, _01206_);
  nand (_10892_, _10891_, _10887_);
  nand (_10893_, _10892_, _01262_);
  nand (_10894_, _10893_, _10883_);
  nand (_10895_, _10894_, _01274_);
  nand (_10896_, _10895_, _10872_);
  nand (_10897_, _10896_, _01241_);
  nand (_10898_, _01296_, _25067_);
  nand (_10899_, _01290_, _25081_);
  nand (_10900_, _10899_, _10898_);
  nand (_10901_, _10900_, _01204_);
  nand (_10902_, _01290_, _25052_);
  nand (_10903_, _01296_, _25038_);
  nand (_10904_, _10903_, _10902_);
  nand (_10905_, _10904_, _01206_);
  nand (_10906_, _10905_, _10901_);
  nand (_10907_, _10906_, _01260_);
  nand (_10908_, _01296_, _25009_);
  nand (_10909_, _01290_, _25024_);
  nand (_10910_, _10909_, _10908_);
  nand (_10911_, _10910_, _01204_);
  nand (_10912_, _01290_, _24995_);
  nand (_10913_, _01296_, _24981_);
  nand (_10914_, _10913_, _10912_);
  nand (_10915_, _10914_, _01206_);
  nand (_10917_, _10915_, _10911_);
  nand (_10918_, _10917_, _01262_);
  nand (_10919_, _10918_, _10907_);
  nand (_10920_, _10919_, _01275_);
  nor (_10921_, _01296_, _24938_);
  nor (_10922_, _01290_, _24922_);
  nor (_10923_, _10922_, _10921_);
  nand (_10924_, _10923_, _01206_);
  nand (_10925_, _01290_, _24966_);
  nand (_10926_, _01296_, _24952_);
  nand (_10927_, _10926_, _10925_);
  nand (_10928_, _10927_, _01204_);
  nand (_10929_, _10928_, _10924_);
  nand (_10930_, _10929_, _01260_);
  nor (_10931_, _01296_, _24879_);
  nor (_10932_, _01290_, _24865_);
  nor (_10933_, _10932_, _10931_);
  nand (_10934_, _10933_, _01206_);
  nand (_10935_, _01290_, _24908_);
  nand (_10936_, _01296_, _24894_);
  nand (_10937_, _10936_, _10935_);
  nand (_10938_, _10937_, _01204_);
  nand (_10939_, _10938_, _10934_);
  nand (_10940_, _10939_, _01262_);
  nand (_10941_, _10940_, _10930_);
  nand (_10942_, _10941_, _01274_);
  nand (_10943_, _10942_, _10920_);
  nand (_10944_, _10943_, _01308_);
  nand (_10945_, _10944_, _10897_);
  nand (_10946_, _10945_, _01245_);
  nand (_10947_, _01296_, _25470_);
  nand (_10948_, _01290_, _25484_);
  nand (_10949_, _10948_, _10947_);
  nand (_10950_, _10949_, _01204_);
  nand (_10951_, _01290_, _25455_);
  nand (_10952_, _01296_, _25441_);
  nand (_10953_, _10952_, _10951_);
  nand (_10954_, _10953_, _01206_);
  nand (_10955_, _10954_, _10950_);
  nand (_10956_, _10955_, _01260_);
  nand (_10958_, _01296_, _25412_);
  nand (_10959_, _01290_, _25427_);
  nand (_10960_, _10959_, _10958_);
  nand (_10961_, _10960_, _01204_);
  nand (_10962_, _01290_, _25398_);
  nand (_10963_, _01296_, _25383_);
  nand (_10964_, _10963_, _10962_);
  nand (_10965_, _10964_, _01206_);
  nand (_10966_, _10965_, _10961_);
  nand (_10967_, _10966_, _01262_);
  nand (_10968_, _10967_, _10956_);
  nand (_10969_, _10968_, _01275_);
  nor (_10970_, _01296_, _25339_);
  nor (_10971_, _01290_, _25325_);
  nor (_10972_, _10971_, _10970_);
  nand (_10973_, _10972_, _01206_);
  nand (_10974_, _01290_, _25369_);
  nand (_10975_, _01296_, _25355_);
  nand (_10976_, _10975_, _10974_);
  nand (_10977_, _10976_, _01204_);
  nand (_10978_, _10977_, _10973_);
  nand (_10979_, _10978_, _01260_);
  nor (_10980_, _01296_, _25282_);
  nor (_10981_, _01290_, _25268_);
  nor (_10982_, _10981_, _10980_);
  nand (_10983_, _10982_, _01206_);
  nand (_10984_, _01290_, _25311_);
  nand (_10985_, _01296_, _25296_);
  nand (_10986_, _10985_, _10984_);
  nand (_10987_, _10986_, _01204_);
  nand (_10989_, _10987_, _10983_);
  nand (_10990_, _10989_, _01262_);
  nand (_10991_, _10990_, _10979_);
  nand (_10992_, _10991_, _01274_);
  nand (_10993_, _10992_, _10969_);
  nand (_10994_, _10993_, _01308_);
  nand (_10995_, _01290_, _25253_);
  nand (_10996_, _01296_, _25239_);
  nand (_10997_, _10996_, _10995_);
  nand (_10998_, _10997_, _01204_);
  nand (_10999_, _01296_, _25210_);
  nand (_11000_, _01290_, _25225_);
  nand (_11001_, _11000_, _10999_);
  nand (_11002_, _11001_, _01206_);
  nand (_11003_, _11002_, _10998_);
  nand (_11004_, _11003_, _01260_);
  nand (_11005_, _01290_, _25196_);
  nand (_11006_, _01296_, _25182_);
  nand (_11007_, _11006_, _11005_);
  nand (_11008_, _11007_, _01204_);
  nand (_11009_, _01296_, _25153_);
  nand (_11010_, _01290_, _25167_);
  nand (_11011_, _11010_, _11009_);
  nand (_11012_, _11011_, _01206_);
  nand (_11013_, _11012_, _11008_);
  nand (_11014_, _11013_, _01262_);
  nand (_11015_, _11014_, _11004_);
  nand (_11016_, _11015_, _01275_);
  nor (_11017_, _01296_, _25139_);
  nor (_11018_, _01290_, _25124_);
  nor (_11019_, _11018_, _11017_);
  nand (_11020_, _11019_, _01204_);
  nor (_11021_, _01290_, _23676_);
  nor (_11022_, _01296_, _25110_);
  nor (_11023_, _11022_, _11021_);
  nand (_11024_, _11023_, _01206_);
  nand (_11025_, _11024_, _11020_);
  nand (_11026_, _11025_, _01260_);
  nor (_11027_, _01296_, _23647_);
  nor (_11028_, _01290_, _23633_);
  nor (_11030_, _11028_, _11027_);
  nand (_11031_, _11030_, _01204_);
  nor (_11032_, _01290_, _25095_);
  nor (_11033_, _01296_, _23661_);
  nor (_11034_, _11033_, _11032_);
  nand (_11035_, _11034_, _01206_);
  nand (_11036_, _11035_, _11031_);
  nand (_11037_, _11036_, _01262_);
  nand (_11038_, _11037_, _11026_);
  nand (_11039_, _11038_, _01274_);
  nand (_11041_, _11039_, _11016_);
  nand (_11042_, _11041_, _01241_);
  nand (_11043_, _11042_, _10994_);
  nand (_11044_, _11043_, _01244_);
  nand (_11045_, _11044_, _10946_);
  nor (_11046_, _11045_, _01231_);
  nand (_11047_, _01296_, _24146_);
  nand (_11048_, _01290_, _24161_);
  nand (_11049_, _11048_, _11047_);
  nand (_11050_, _11049_, _01204_);
  nand (_11051_, _01290_, _24132_);
  nand (_11052_, _01296_, _24118_);
  nand (_11053_, _11052_, _11051_);
  nand (_11054_, _11053_, _01206_);
  nand (_11055_, _11054_, _11050_);
  nand (_11056_, _11055_, _01260_);
  nand (_11057_, _01296_, _24088_);
  nand (_11058_, _01290_, _24102_);
  nand (_11059_, _11058_, _11057_);
  nand (_11060_, _11059_, _01204_);
  nand (_11061_, _01290_, _24074_);
  nand (_11062_, _01296_, _24059_);
  nand (_11063_, _11062_, _11061_);
  nand (_11064_, _11063_, _01206_);
  nand (_11065_, _11064_, _11060_);
  nand (_11066_, _11065_, _01262_);
  nand (_11067_, _11066_, _11056_);
  nand (_11068_, _11067_, _01275_);
  nor (_11069_, _01296_, _24016_);
  nor (_11070_, _01290_, _24002_);
  nor (_11072_, _11070_, _11069_);
  nand (_11073_, _11072_, _01206_);
  nand (_11074_, _01290_, _24045_);
  nand (_11075_, _01296_, _24031_);
  nand (_11076_, _11075_, _11074_);
  nand (_11077_, _11076_, _01204_);
  nand (_11078_, _11077_, _11073_);
  nand (_11079_, _11078_, _01260_);
  nor (_11080_, _01296_, _23959_);
  nor (_11081_, _01290_, _23944_);
  nor (_11082_, _11081_, _11080_);
  nand (_11083_, _11082_, _01206_);
  nand (_11084_, _01290_, _23988_);
  nand (_11085_, _01296_, _23973_);
  nand (_11086_, _11085_, _11084_);
  nand (_11087_, _11086_, _01204_);
  nand (_11088_, _11087_, _11083_);
  nand (_11089_, _11088_, _01262_);
  nand (_11090_, _11089_, _11079_);
  nand (_11091_, _11090_, _01274_);
  nand (_11092_, _11091_, _11068_);
  nand (_11093_, _11092_, _01308_);
  nand (_11094_, _01290_, _23930_);
  nand (_11095_, _01296_, _23916_);
  nand (_11096_, _11095_, _11094_);
  nand (_11097_, _11096_, _01204_);
  nand (_11098_, _01296_, _23887_);
  nand (_11099_, _01290_, _23901_);
  nand (_11100_, _11099_, _11098_);
  nand (_11101_, _11100_, _01206_);
  nand (_11102_, _11101_, _11097_);
  nand (_11103_, _11102_, _01260_);
  nand (_11104_, _01290_, _23873_);
  nand (_11105_, _01296_, _23858_);
  nand (_11106_, _11105_, _11104_);
  nand (_11107_, _11106_, _01204_);
  nand (_11108_, _01296_, _23830_);
  nand (_11109_, _01290_, _23844_);
  nand (_11110_, _11109_, _11108_);
  nand (_11111_, _11110_, _01206_);
  nand (_11113_, _11111_, _11107_);
  nand (_11114_, _11113_, _01262_);
  nand (_11115_, _11114_, _11103_);
  nand (_11116_, _11115_, _01275_);
  nor (_11117_, _01296_, _23815_);
  nor (_11118_, _01290_, _23801_);
  nor (_11119_, _11118_, _11117_);
  nand (_11120_, _11119_, _01204_);
  nor (_11121_, _01290_, _23772_);
  nor (_11122_, _01296_, _23787_);
  nor (_11123_, _11122_, _11121_);
  nand (_11124_, _11123_, _01206_);
  nand (_11125_, _11124_, _11120_);
  nand (_11126_, _11125_, _01260_);
  nor (_11127_, _01296_, _23758_);
  nor (_11128_, _01290_, _23744_);
  nor (_11129_, _11128_, _11127_);
  nand (_11130_, _11129_, _01204_);
  nor (_11131_, _01290_, _23715_);
  nor (_11132_, _01296_, _23729_);
  nor (_11133_, _11132_, _11131_);
  nand (_11134_, _11133_, _01206_);
  nand (_11135_, _11134_, _11130_);
  nand (_11136_, _11135_, _01262_);
  nand (_11137_, _11136_, _11126_);
  nand (_11138_, _11137_, _01274_);
  nand (_11139_, _11138_, _11116_);
  nand (_11140_, _11139_, _01241_);
  nand (_11141_, _11140_, _11093_);
  nand (_11142_, _11141_, _01245_);
  nor (_11143_, _01296_, _24218_);
  nor (_11144_, _01290_, _24204_);
  nor (_11145_, _11144_, _11143_);
  nand (_11146_, _11145_, _01204_);
  nor (_11147_, _01290_, _24175_);
  nor (_11148_, _01296_, _24189_);
  nor (_11149_, _11148_, _11147_);
  nand (_11150_, _11149_, _01206_);
  nand (_11151_, _11150_, _11146_);
  nand (_11152_, _11151_, _01262_);
  nor (_11154_, _01296_, _24276_);
  nor (_11155_, _01290_, _24261_);
  nor (_11156_, _11155_, _11154_);
  nand (_11157_, _11156_, _01204_);
  nor (_11158_, _01290_, _24232_);
  nor (_11159_, _01296_, _24247_);
  nor (_11160_, _11159_, _11158_);
  nand (_11161_, _11160_, _01206_);
  nand (_11162_, _11161_, _11157_);
  nand (_11163_, _11162_, _01260_);
  nand (_11164_, _11163_, _11152_);
  nand (_11165_, _11164_, _01274_);
  nand (_11166_, _01290_, _24333_);
  nand (_11167_, _01296_, _24319_);
  nand (_11168_, _11167_, _11166_);
  nand (_11169_, _11168_, _01204_);
  nand (_11170_, _01296_, _24290_);
  nand (_11171_, _01290_, _24304_);
  nand (_11172_, _11171_, _11170_);
  nand (_11173_, _11172_, _01206_);
  nand (_11174_, _11173_, _11169_);
  nand (_11175_, _11174_, _01262_);
  nand (_11176_, _01290_, _24390_);
  nand (_11177_, _01296_, _24376_);
  nand (_11178_, _11177_, _11176_);
  nand (_11179_, _11178_, _01204_);
  nand (_11180_, _01296_, _24347_);
  nand (_11181_, _01290_, _24362_);
  nand (_11182_, _11181_, _11180_);
  nand (_11183_, _11182_, _01206_);
  nand (_11184_, _11183_, _11179_);
  nand (_11185_, _11184_, _01260_);
  nand (_11186_, _11185_, _11175_);
  nand (_11187_, _11186_, _01275_);
  nand (_11188_, _11187_, _11165_);
  nand (_11189_, _11188_, _01241_);
  nor (_11190_, _01296_, _24419_);
  nor (_11191_, _01290_, _24405_);
  nor (_11192_, _11191_, _11190_);
  nand (_11193_, _11192_, _01206_);
  nand (_11195_, _01290_, _24448_);
  nand (_11196_, _01296_, _24433_);
  nand (_11197_, _11196_, _11195_);
  nand (_11198_, _11197_, _01204_);
  nand (_11199_, _11198_, _11193_);
  nand (_11200_, _11199_, _01262_);
  nor (_11201_, _01296_, _24476_);
  nor (_11202_, _01290_, _24462_);
  nor (_11203_, _11202_, _11201_);
  nand (_11204_, _11203_, _01206_);
  nand (_11205_, _01290_, _24505_);
  nand (_11206_, _01296_, _24491_);
  nand (_11207_, _11206_, _11205_);
  nand (_11208_, _11207_, _01204_);
  nand (_11209_, _11208_, _11204_);
  nand (_11210_, _11209_, _01260_);
  nand (_11211_, _11210_, _11200_);
  nand (_11212_, _11211_, _01274_);
  nand (_11213_, _01296_, _24549_);
  nand (_11214_, _01290_, _24564_);
  nand (_11215_, _11214_, _11213_);
  nand (_11216_, _11215_, _01204_);
  nand (_11217_, _01290_, _24535_);
  nand (_11218_, _01296_, _24519_);
  nand (_11219_, _11218_, _11217_);
  nand (_11220_, _11219_, _01206_);
  nand (_11221_, _11220_, _11216_);
  nand (_11222_, _11221_, _01262_);
  nand (_11223_, _01296_, _24607_);
  nand (_11224_, _01290_, _24621_);
  nand (_11225_, _11224_, _11223_);
  nand (_11226_, _11225_, _01204_);
  nand (_11227_, _01290_, _24592_);
  nand (_11228_, _01296_, _24578_);
  nand (_11229_, _11228_, _11227_);
  nand (_11230_, _11229_, _01206_);
  nand (_11231_, _11230_, _11226_);
  nand (_11232_, _11231_, _01260_);
  nand (_11233_, _11232_, _11222_);
  nand (_11234_, _11233_, _01275_);
  nand (_11236_, _11234_, _11212_);
  nand (_11237_, _11236_, _01308_);
  nand (_11238_, _11237_, _11189_);
  nand (_11239_, _11238_, _01244_);
  nand (_11240_, _11239_, _11142_);
  nor (_11241_, _11240_, _01235_);
  nor (_11242_, _11241_, _11046_);
  nor (_11243_, _11242_, _28718_);
  nor (_11244_, _11243_, _10850_);
  nor (_11245_, _11244_, _06280_);
  nand (_11246_, _06280_, _27651_);
  nand (_11247_, _11246_, _29344_);
  nor (_15188_, _11247_, _11245_);
  nand (_11248_, _01290_, _27573_);
  nand (_11249_, _01296_, _27545_);
  nand (_11250_, _11249_, _11248_);
  nand (_11251_, _11250_, _01204_);
  nand (_11252_, _01296_, _23606_);
  nand (_11253_, _01290_, _27515_);
  nand (_11254_, _11253_, _11252_);
  nand (_11255_, _11254_, _01206_);
  nand (_11256_, _11255_, _11251_);
  nand (_11257_, _11256_, _01260_);
  nand (_11258_, _01290_, _23703_);
  nand (_11259_, _01296_, _23620_);
  nand (_11260_, _11259_, _11258_);
  nand (_11261_, _11260_, _01204_);
  nand (_11262_, _01296_, _27459_);
  nand (_11263_, _01290_, _27487_);
  nand (_11264_, _11263_, _11262_);
  nand (_11265_, _11264_, _01206_);
  nand (_11266_, _11265_, _11261_);
  nand (_11267_, _11266_, _01262_);
  nand (_11268_, _11267_, _11257_);
  nand (_11269_, _11268_, _01275_);
  nor (_11270_, _01296_, _27430_);
  nor (_11271_, _01290_, _27402_);
  nor (_11272_, _11271_, _11270_);
  nand (_11273_, _11272_, _01204_);
  nor (_11274_, _01290_, _27345_);
  nor (_11276_, _01296_, _27373_);
  nor (_11277_, _11276_, _11274_);
  nand (_11278_, _11277_, _01206_);
  nand (_11279_, _11278_, _11273_);
  nand (_11280_, _11279_, _01260_);
  nor (_11281_, _01296_, _27317_);
  nor (_11282_, _01290_, _27288_);
  nor (_11283_, _11282_, _11281_);
  nand (_11284_, _11283_, _01204_);
  nor (_11285_, _01290_, _27232_);
  nor (_11286_, _01296_, _27260_);
  nor (_11287_, _11286_, _11285_);
  nand (_11288_, _11287_, _01206_);
  nand (_11289_, _11288_, _11284_);
  nand (_11290_, _11289_, _01262_);
  nand (_11291_, _11290_, _11280_);
  nand (_11292_, _11291_, _01274_);
  nand (_11293_, _11292_, _11269_);
  nand (_11294_, _11293_, _01241_);
  nand (_11295_, _01296_, _23563_);
  nand (_11296_, _01290_, _27941_);
  nand (_11297_, _11296_, _11295_);
  nand (_11298_, _11297_, _01204_);
  nand (_11299_, _01290_, _27913_);
  nand (_11300_, _01296_, _23577_);
  nand (_11301_, _11300_, _11299_);
  nand (_11302_, _11301_, _01206_);
  nand (_11303_, _11302_, _11298_);
  nand (_11304_, _11303_, _01260_);
  nand (_11305_, _01296_, _27856_);
  nand (_11306_, _01290_, _27885_);
  nand (_11307_, _11306_, _11305_);
  nand (_11308_, _11307_, _01204_);
  nand (_11309_, _01290_, _27828_);
  nand (_11310_, _01296_, _27800_);
  nand (_11311_, _11310_, _11309_);
  nand (_11312_, _11311_, _01206_);
  nand (_11313_, _11312_, _11308_);
  nand (_11314_, _11313_, _01262_);
  nand (_11315_, _11314_, _11304_);
  nand (_11317_, _11315_, _01275_);
  nor (_11318_, _01296_, _27715_);
  nor (_11319_, _01290_, _27686_);
  nor (_11320_, _11319_, _11318_);
  nand (_11321_, _11320_, _01206_);
  nand (_11322_, _01290_, _27771_);
  nand (_11323_, _01296_, _27743_);
  nand (_11324_, _11323_, _11322_);
  nand (_11325_, _11324_, _01204_);
  nand (_11326_, _11325_, _11321_);
  nand (_11327_, _11326_, _01260_);
  nor (_11328_, _01296_, _27630_);
  nor (_11329_, _01290_, _27601_);
  nor (_11330_, _11329_, _11328_);
  nand (_11331_, _11330_, _01206_);
  nand (_11332_, _01290_, _23592_);
  nand (_11333_, _01296_, _27658_);
  nand (_11334_, _11333_, _11332_);
  nand (_11335_, _11334_, _01204_);
  nand (_11336_, _11335_, _11331_);
  nand (_11337_, _11336_, _01262_);
  nand (_11338_, _11337_, _11327_);
  nand (_11339_, _11338_, _01274_);
  nand (_11340_, _11339_, _11317_);
  nand (_11341_, _11340_, _01308_);
  nand (_11342_, _11341_, _11294_);
  nand (_11343_, _11342_, _01245_);
  nand (_11344_, _01296_, _28396_);
  nand (_11345_, _01290_, _28424_);
  nand (_11346_, _11345_, _11344_);
  nand (_11347_, _11346_, _01204_);
  nand (_11348_, _01290_, _28368_);
  nand (_11349_, _01296_, _28310_);
  nand (_11350_, _11349_, _11348_);
  nand (_11351_, _11350_, _01206_);
  nand (_11352_, _11351_, _11347_);
  nand (_11353_, _11352_, _01260_);
  nand (_11354_, _01296_, _28253_);
  nand (_11355_, _01290_, _28282_);
  nand (_11356_, _11355_, _11354_);
  nand (_11358_, _11356_, _01204_);
  nand (_11359_, _01290_, _28197_);
  nand (_11360_, _01296_, _28168_);
  nand (_11361_, _11360_, _11359_);
  nand (_11362_, _11361_, _01206_);
  nand (_11363_, _11362_, _11358_);
  nand (_11364_, _11363_, _01262_);
  nand (_11365_, _11364_, _11353_);
  nand (_11366_, _11365_, _01275_);
  nor (_11367_, _01296_, _28083_);
  nor (_11368_, _01290_, _23506_);
  nor (_11369_, _11368_, _11367_);
  nand (_11370_, _11369_, _01206_);
  nand (_11371_, _01290_, _28140_);
  nand (_11372_, _01296_, _28112_);
  nand (_11373_, _11372_, _11371_);
  nand (_11374_, _11373_, _01204_);
  nand (_11375_, _11374_, _11370_);
  nand (_11376_, _11375_, _01260_);
  nor (_11377_, _01296_, _23463_);
  nor (_11378_, _01290_, _23448_);
  nor (_11379_, _11378_, _11377_);
  nand (_11380_, _11379_, _01206_);
  nand (_11381_, _01290_, _23491_);
  nand (_11382_, _01296_, _23477_);
  nand (_11383_, _11382_, _11381_);
  nand (_11384_, _11383_, _01204_);
  nand (_11385_, _11384_, _11380_);
  nand (_11386_, _11385_, _01262_);
  nand (_11387_, _11386_, _11376_);
  nand (_11388_, _11387_, _01274_);
  nand (_11389_, _11388_, _11366_);
  nand (_11390_, _11389_, _01308_);
  nand (_11391_, _01290_, _23434_);
  nand (_11392_, _01296_, _23420_);
  nand (_11393_, _11392_, _11391_);
  nand (_11394_, _11393_, _01204_);
  nand (_11395_, _01296_, _23391_);
  nand (_11396_, _01290_, _23405_);
  nand (_11397_, _11396_, _11395_);
  nand (_11399_, _11397_, _01206_);
  nand (_11400_, _11399_, _11394_);
  nand (_11401_, _11400_, _01260_);
  nand (_11402_, _01290_, _23377_);
  nand (_11403_, _01296_, _23362_);
  nand (_11404_, _11403_, _11402_);
  nand (_11405_, _11404_, _01204_);
  nand (_11406_, _01296_, _28225_);
  nand (_11407_, _01290_, _28441_);
  nand (_11408_, _11407_, _11406_);
  nand (_11409_, _11408_, _01206_);
  nand (_11410_, _11409_, _11405_);
  nand (_11411_, _11410_, _01262_);
  nand (_11412_, _11411_, _11401_);
  nand (_11413_, _11412_, _01275_);
  nor (_11414_, _01296_, _28338_);
  nor (_11415_, _01290_, _23534_);
  nor (_11416_, _11415_, _11414_);
  nand (_11417_, _11416_, _01204_);
  nor (_11418_, _01290_, _28055_);
  nor (_11419_, _01296_, _23520_);
  nor (_11420_, _11419_, _11418_);
  nand (_11421_, _11420_, _01206_);
  nand (_11422_, _11421_, _11417_);
  nand (_11423_, _11422_, _01260_);
  nor (_11424_, _01296_, _28027_);
  nor (_11425_, _01290_, _27998_);
  nor (_11426_, _11425_, _11424_);
  nand (_11427_, _11426_, _01204_);
  nor (_11428_, _01290_, _23549_);
  nor (_11429_, _01296_, _27970_);
  nor (_11430_, _11429_, _11428_);
  nand (_11431_, _11430_, _01206_);
  nand (_11432_, _11431_, _11427_);
  nand (_11433_, _11432_, _01262_);
  nand (_11434_, _11433_, _11423_);
  nand (_11435_, _11434_, _01274_);
  nand (_11436_, _11435_, _11413_);
  nand (_11437_, _11436_, _01241_);
  nand (_11438_, _11437_, _11390_);
  nand (_11440_, _11438_, _01244_);
  nand (_11441_, _11440_, _11343_);
  nor (_11442_, _11441_, _01231_);
  nand (_11443_, _01296_, _26267_);
  nand (_11444_, _01290_, _26295_);
  nand (_11445_, _11444_, _11443_);
  nand (_11446_, _11445_, _01204_);
  nand (_11447_, _01290_, _26238_);
  nand (_11448_, _01296_, _26210_);
  nand (_11449_, _11448_, _11447_);
  nand (_11451_, _11449_, _01206_);
  nand (_11452_, _11451_, _11446_);
  nand (_11453_, _11452_, _01260_);
  nand (_11454_, _01296_, _26153_);
  nand (_11455_, _01290_, _26182_);
  nand (_11456_, _11455_, _11454_);
  nand (_11457_, _11456_, _01204_);
  nand (_11458_, _01290_, _26125_);
  nand (_11459_, _01296_, _26097_);
  nand (_11460_, _11459_, _11458_);
  nand (_11461_, _11460_, _01206_);
  nand (_11462_, _11461_, _11457_);
  nand (_11463_, _11462_, _01262_);
  nand (_11464_, _11463_, _11453_);
  nand (_11465_, _11464_, _01275_);
  nor (_11466_, _01296_, _26012_);
  nor (_11467_, _01290_, _25983_);
  nor (_11468_, _11467_, _11466_);
  nand (_11469_, _11468_, _01206_);
  nand (_11470_, _01290_, _26068_);
  nand (_11471_, _01296_, _26040_);
  nand (_11472_, _11471_, _11470_);
  nand (_11473_, _11472_, _01204_);
  nand (_11474_, _11473_, _11469_);
  nand (_11475_, _11474_, _01260_);
  nor (_11476_, _01296_, _25897_);
  nor (_11477_, _01290_, _25869_);
  nor (_11478_, _11477_, _11476_);
  nand (_11479_, _11478_, _01206_);
  nand (_11480_, _01290_, _25955_);
  nand (_11482_, _01296_, _25927_);
  nand (_11483_, _11482_, _11480_);
  nand (_11484_, _11483_, _01204_);
  nand (_11485_, _11484_, _11479_);
  nand (_11486_, _11485_, _01262_);
  nand (_11487_, _11486_, _11475_);
  nand (_11488_, _11487_, _01274_);
  nand (_11489_, _11488_, _11465_);
  nand (_11490_, _11489_, _01308_);
  nand (_11491_, _01290_, _25841_);
  nand (_11492_, _01296_, _25812_);
  nand (_11493_, _11492_, _11491_);
  nand (_11494_, _11493_, _01204_);
  nand (_11495_, _01296_, _25756_);
  nand (_11496_, _01290_, _25784_);
  nand (_11497_, _11496_, _11495_);
  nand (_11498_, _11497_, _01206_);
  nand (_11499_, _11498_, _11494_);
  nand (_11500_, _11499_, _01260_);
  nand (_11501_, _01290_, _25727_);
  nand (_11502_, _01296_, _25699_);
  nand (_11503_, _11502_, _11501_);
  nand (_11504_, _11503_, _01204_);
  nand (_11505_, _01296_, _25642_);
  nand (_11506_, _01290_, _25670_);
  nand (_11507_, _11506_, _11505_);
  nand (_11508_, _11507_, _01206_);
  nand (_11509_, _11508_, _11504_);
  nand (_11510_, _11509_, _01262_);
  nand (_11511_, _11510_, _11500_);
  nand (_11512_, _11511_, _01275_);
  nor (_11513_, _01296_, _25614_);
  nor (_11514_, _01290_, _25586_);
  nor (_11515_, _11514_, _11513_);
  nand (_11516_, _11515_, _01204_);
  nor (_11517_, _01290_, _25558_);
  nor (_11518_, _01296_, _25572_);
  nor (_11519_, _11518_, _11517_);
  nand (_11520_, _11519_, _01206_);
  nand (_11521_, _11520_, _11516_);
  nand (_11523_, _11521_, _01260_);
  nor (_11524_, _01296_, _25543_);
  nor (_11525_, _01290_, _25529_);
  nor (_11526_, _11525_, _11524_);
  nand (_11527_, _11526_, _01204_);
  nor (_11528_, _01290_, _25500_);
  nor (_11529_, _01296_, _25515_);
  nor (_11530_, _11529_, _11528_);
  nand (_11531_, _11530_, _01206_);
  nand (_11532_, _11531_, _11527_);
  nand (_11533_, _11532_, _01262_);
  nand (_11534_, _11533_, _11523_);
  nand (_11535_, _11534_, _01274_);
  nand (_11536_, _11535_, _11512_);
  nand (_11537_, _11536_, _01241_);
  nand (_11538_, _11537_, _11490_);
  nand (_11539_, _11538_, _01245_);
  nor (_11540_, _01296_, _26409_);
  nor (_11541_, _01290_, _26380_);
  nor (_11542_, _11541_, _11540_);
  nand (_11543_, _11542_, _01204_);
  nor (_11544_, _01290_, _26324_);
  nor (_11545_, _01296_, _26352_);
  nor (_11546_, _11545_, _11544_);
  nand (_11547_, _11546_, _01206_);
  nand (_11548_, _11547_, _11543_);
  nand (_11549_, _11548_, _01262_);
  nor (_11550_, _01296_, _26522_);
  nor (_11551_, _01290_, _26494_);
  nor (_11552_, _11551_, _11550_);
  nand (_11553_, _11552_, _01204_);
  nor (_11554_, _01290_, _26437_);
  nor (_11555_, _01296_, _26465_);
  nor (_11556_, _11555_, _11554_);
  nand (_11557_, _11556_, _01206_);
  nand (_11558_, _11557_, _11553_);
  nand (_11559_, _11558_, _01260_);
  nand (_11560_, _11559_, _11549_);
  nand (_11561_, _11560_, _01274_);
  nand (_11562_, _01290_, _26635_);
  nand (_11564_, _01296_, _26607_);
  nand (_11565_, _11564_, _11562_);
  nand (_11566_, _11565_, _01204_);
  nand (_11567_, _01296_, _26550_);
  nand (_11568_, _01290_, _26579_);
  nand (_11569_, _11568_, _11567_);
  nand (_11570_, _11569_, _01206_);
  nand (_11571_, _11570_, _11566_);
  nand (_11572_, _11571_, _01262_);
  nand (_11573_, _01290_, _26750_);
  nand (_11574_, _01296_, _26720_);
  nand (_11575_, _11574_, _11573_);
  nand (_11576_, _11575_, _01204_);
  nand (_11577_, _01296_, _26664_);
  nand (_11578_, _01290_, _26692_);
  nand (_11579_, _11578_, _11577_);
  nand (_11580_, _11579_, _01206_);
  nand (_11581_, _11580_, _11576_);
  nand (_11582_, _11581_, _01260_);
  nand (_11583_, _11582_, _11572_);
  nand (_11584_, _11583_, _01275_);
  nand (_11585_, _11584_, _11561_);
  nand (_11586_, _11585_, _01241_);
  nor (_11587_, _01296_, _26806_);
  nor (_11588_, _01290_, _26778_);
  nor (_11589_, _11588_, _11587_);
  nand (_11590_, _11589_, _01206_);
  nand (_11591_, _01290_, _26863_);
  nand (_11592_, _01296_, _26835_);
  nand (_11593_, _11592_, _11591_);
  nand (_11594_, _11593_, _01204_);
  nand (_11595_, _11594_, _11590_);
  nand (_11596_, _11595_, _01262_);
  nor (_11597_, _01296_, _26920_);
  nor (_11598_, _01290_, _26892_);
  nor (_11599_, _11598_, _11597_);
  nand (_11600_, _11599_, _01206_);
  nand (_11601_, _01290_, _26977_);
  nand (_11602_, _01296_, _26948_);
  nand (_11603_, _11602_, _11601_);
  nand (_11605_, _11603_, _01204_);
  nand (_11606_, _11605_, _11600_);
  nand (_11607_, _11606_, _01260_);
  nand (_11608_, _11607_, _11596_);
  nand (_11609_, _11608_, _01274_);
  nand (_11610_, _01296_, _27062_);
  nand (_11611_, _01290_, _27090_);
  nand (_11612_, _11611_, _11610_);
  nand (_11613_, _11612_, _01204_);
  nand (_11614_, _01290_, _27033_);
  nand (_11615_, _01296_, _27005_);
  nand (_11616_, _11615_, _11614_);
  nand (_11617_, _11616_, _01206_);
  nand (_11618_, _11617_, _11613_);
  nand (_11619_, _11618_, _01262_);
  nand (_11620_, _01296_, _27175_);
  nand (_11621_, _01290_, _27203_);
  nand (_11622_, _11621_, _11620_);
  nand (_11623_, _11622_, _01204_);
  nand (_11624_, _01290_, _27147_);
  nand (_11625_, _01296_, _27118_);
  nand (_11626_, _11625_, _11624_);
  nand (_11627_, _11626_, _01206_);
  nand (_11628_, _11627_, _11623_);
  nand (_11629_, _11628_, _01260_);
  nand (_11630_, _11629_, _11619_);
  nand (_11631_, _11630_, _01275_);
  nand (_11632_, _11631_, _11609_);
  nand (_11633_, _11632_, _01308_);
  nand (_11634_, _11633_, _11586_);
  nand (_11635_, _11634_, _01244_);
  nand (_11636_, _11635_, _11539_);
  nor (_11637_, _11636_, _01235_);
  nor (_11638_, _11637_, _11442_);
  nor (_11639_, _11638_, _28717_);
  nand (_11640_, _01290_, _24853_);
  nand (_11641_, _01296_, _24838_);
  nand (_11642_, _11641_, _11640_);
  nand (_11643_, _11642_, _01204_);
  nand (_11644_, _01296_, _24810_);
  nand (_11646_, _01290_, _24824_);
  nand (_11647_, _11646_, _11644_);
  nand (_11648_, _11647_, _01206_);
  nand (_11649_, _11648_, _11643_);
  nand (_11650_, _11649_, _01260_);
  nand (_11651_, _01290_, _24795_);
  nand (_11652_, _01296_, _24781_);
  nand (_11653_, _11652_, _11651_);
  nand (_11654_, _11653_, _01204_);
  nand (_11655_, _01296_, _24752_);
  nand (_11656_, _01290_, _24766_);
  nand (_11657_, _11656_, _11655_);
  nand (_11658_, _11657_, _01206_);
  nand (_11659_, _11658_, _11654_);
  nand (_11660_, _11659_, _01262_);
  nand (_11661_, _11660_, _11650_);
  nand (_11662_, _11661_, _01275_);
  nor (_11663_, _01296_, _24738_);
  nor (_11664_, _01290_, _24723_);
  nor (_11665_, _11664_, _11663_);
  nand (_11666_, _11665_, _01204_);
  nor (_11667_, _01290_, _24695_);
  nor (_11668_, _01296_, _24709_);
  nor (_11669_, _11668_, _11667_);
  nand (_11670_, _11669_, _01206_);
  nand (_11671_, _11670_, _11666_);
  nand (_11672_, _11671_, _01260_);
  nor (_11673_, _01296_, _24680_);
  nor (_11674_, _01290_, _24666_);
  nor (_11675_, _11674_, _11673_);
  nand (_11676_, _11675_, _01204_);
  nor (_11677_, _01290_, _24637_);
  nor (_11678_, _01296_, _24652_);
  nor (_11679_, _11678_, _11677_);
  nand (_11680_, _11679_, _01206_);
  nand (_11681_, _11680_, _11676_);
  nand (_11682_, _11681_, _01262_);
  nand (_11683_, _11682_, _11672_);
  nand (_11684_, _11683_, _01274_);
  nand (_11685_, _11684_, _11662_);
  nand (_11687_, _11685_, _01241_);
  nand (_11688_, _01296_, _25069_);
  nand (_11689_, _01290_, _25083_);
  nand (_11690_, _11689_, _11688_);
  nand (_11691_, _11690_, _01204_);
  nand (_11692_, _01290_, _25054_);
  nand (_11693_, _01296_, _25040_);
  nand (_11694_, _11693_, _11692_);
  nand (_11695_, _11694_, _01206_);
  nand (_11696_, _11695_, _11691_);
  nand (_11697_, _11696_, _01260_);
  nand (_11698_, _01296_, _25011_);
  nand (_11699_, _01290_, _25026_);
  nand (_11700_, _11699_, _11698_);
  nand (_11701_, _11700_, _01204_);
  nand (_11702_, _01290_, _24997_);
  nand (_11703_, _01296_, _24983_);
  nand (_11704_, _11703_, _11702_);
  nand (_11705_, _11704_, _01206_);
  nand (_11706_, _11705_, _11701_);
  nand (_11707_, _11706_, _01262_);
  nand (_11708_, _11707_, _11697_);
  nand (_11709_, _11708_, _01275_);
  nor (_11710_, _01296_, _24940_);
  nor (_11711_, _01290_, _24924_);
  nor (_11712_, _11711_, _11710_);
  nand (_11713_, _11712_, _01206_);
  nand (_11714_, _01290_, _24968_);
  nand (_11715_, _01296_, _24954_);
  nand (_11716_, _11715_, _11714_);
  nand (_11717_, _11716_, _01204_);
  nand (_11718_, _11717_, _11713_);
  nand (_11719_, _11718_, _01260_);
  nor (_11720_, _01296_, _24881_);
  nor (_11721_, _01290_, _24867_);
  nor (_11722_, _11721_, _11720_);
  nand (_11723_, _11722_, _01206_);
  nand (_11724_, _01290_, _24910_);
  nand (_11725_, _01296_, _24896_);
  nand (_11726_, _11725_, _11724_);
  nand (_11728_, _11726_, _01204_);
  nand (_11729_, _11728_, _11723_);
  nand (_11730_, _11729_, _01262_);
  nand (_11731_, _11730_, _11719_);
  nand (_11732_, _11731_, _01274_);
  nand (_11733_, _11732_, _11709_);
  nand (_11734_, _11733_, _01308_);
  nand (_11735_, _11734_, _11687_);
  nand (_11736_, _11735_, _01245_);
  nand (_11737_, _01296_, _25472_);
  nand (_11738_, _01290_, _25486_);
  nand (_11739_, _11738_, _11737_);
  nand (_11740_, _11739_, _01204_);
  nand (_11741_, _01290_, _25457_);
  nand (_11742_, _01296_, _25443_);
  nand (_11743_, _11742_, _11741_);
  nand (_11744_, _11743_, _01206_);
  nand (_11745_, _11744_, _11740_);
  nand (_11746_, _11745_, _01260_);
  nand (_11747_, _01296_, _25414_);
  nand (_11748_, _01290_, _25429_);
  nand (_11749_, _11748_, _11747_);
  nand (_11750_, _11749_, _01204_);
  nand (_11751_, _01290_, _25400_);
  nand (_11752_, _01296_, _25386_);
  nand (_11753_, _11752_, _11751_);
  nand (_11754_, _11753_, _01206_);
  nand (_11755_, _11754_, _11750_);
  nand (_11756_, _11755_, _01262_);
  nand (_11757_, _11756_, _11746_);
  nand (_11758_, _11757_, _01275_);
  nor (_11759_, _01296_, _25341_);
  nor (_11760_, _01290_, _25327_);
  nor (_11761_, _11760_, _11759_);
  nand (_11762_, _11761_, _01206_);
  nand (_11763_, _01290_, _25371_);
  nand (_11764_, _01296_, _25357_);
  nand (_11765_, _11764_, _11763_);
  nand (_11766_, _11765_, _01204_);
  nand (_11767_, _11766_, _11762_);
  nand (_11769_, _11767_, _01260_);
  nor (_11770_, _01296_, _25284_);
  nor (_11771_, _01290_, _25270_);
  nor (_11772_, _11771_, _11770_);
  nand (_11773_, _11772_, _01206_);
  nand (_11774_, _01290_, _25313_);
  nand (_11775_, _01296_, _25298_);
  nand (_11776_, _11775_, _11774_);
  nand (_11777_, _11776_, _01204_);
  nand (_11778_, _11777_, _11773_);
  nand (_11779_, _11778_, _01262_);
  nand (_11780_, _11779_, _11769_);
  nand (_11781_, _11780_, _01274_);
  nand (_11782_, _11781_, _11758_);
  nand (_11783_, _11782_, _01308_);
  nand (_11784_, _01290_, _25255_);
  nand (_11785_, _01296_, _25241_);
  nand (_11786_, _11785_, _11784_);
  nand (_11787_, _11786_, _01204_);
  nand (_11788_, _01296_, _25212_);
  nand (_11789_, _01290_, _25227_);
  nand (_11790_, _11789_, _11788_);
  nand (_11791_, _11790_, _01206_);
  nand (_11792_, _11791_, _11787_);
  nand (_11793_, _11792_, _01260_);
  nand (_11794_, _01290_, _25198_);
  nand (_11795_, _01296_, _25184_);
  nand (_11796_, _11795_, _11794_);
  nand (_11797_, _11796_, _01204_);
  nand (_11798_, _01296_, _25155_);
  nand (_11799_, _01290_, _25169_);
  nand (_11800_, _11799_, _11798_);
  nand (_11801_, _11800_, _01206_);
  nand (_11802_, _11801_, _11797_);
  nand (_11803_, _11802_, _01262_);
  nand (_11804_, _11803_, _11793_);
  nand (_11805_, _11804_, _01275_);
  nor (_11806_, _01296_, _25141_);
  nor (_11807_, _01290_, _25126_);
  nor (_11808_, _11807_, _11806_);
  nand (_11810_, _11808_, _01204_);
  nor (_11811_, _01290_, _23678_);
  nor (_11812_, _01296_, _25112_);
  nor (_11813_, _11812_, _11811_);
  nand (_11814_, _11813_, _01206_);
  nand (_11815_, _11814_, _11810_);
  nand (_11816_, _11815_, _01260_);
  nor (_11817_, _01296_, _23649_);
  nor (_11818_, _01290_, _23635_);
  nor (_11819_, _11818_, _11817_);
  nand (_11820_, _11819_, _01204_);
  nor (_11821_, _01290_, _25098_);
  nor (_11822_, _01296_, _23664_);
  nor (_11823_, _11822_, _11821_);
  nand (_11824_, _11823_, _01206_);
  nand (_11825_, _11824_, _11820_);
  nand (_11826_, _11825_, _01262_);
  nand (_11827_, _11826_, _11816_);
  nand (_11828_, _11827_, _01274_);
  nand (_11829_, _11828_, _11805_);
  nand (_11830_, _11829_, _01241_);
  nand (_11831_, _11830_, _11783_);
  nand (_11832_, _11831_, _01244_);
  nand (_11833_, _11832_, _11736_);
  nor (_11834_, _11833_, _01231_);
  nand (_11835_, _01296_, _24148_);
  nand (_11836_, _01290_, _24163_);
  nand (_11837_, _11836_, _11835_);
  nand (_11838_, _11837_, _01204_);
  nand (_11839_, _01290_, _24134_);
  nand (_11840_, _01296_, _24120_);
  nand (_11841_, _11840_, _11839_);
  nand (_11842_, _11841_, _01206_);
  nand (_11843_, _11842_, _11838_);
  nand (_11844_, _11843_, _01260_);
  nand (_11845_, _01296_, _24090_);
  nand (_11846_, _01290_, _24104_);
  nand (_11847_, _11846_, _11845_);
  nand (_11848_, _11847_, _01204_);
  nand (_11849_, _01290_, _24076_);
  nand (_11851_, _01296_, _24061_);
  nand (_11852_, _11851_, _11849_);
  nand (_11853_, _11852_, _01206_);
  nand (_11854_, _11853_, _11848_);
  nand (_11855_, _11854_, _01262_);
  nand (_11856_, _11855_, _11844_);
  nand (_11857_, _11856_, _01275_);
  nor (_11858_, _01296_, _24018_);
  nor (_11859_, _01290_, _24004_);
  nor (_11860_, _11859_, _11858_);
  nand (_11862_, _11860_, _01206_);
  nand (_11863_, _01290_, _24047_);
  nand (_11864_, _01296_, _24033_);
  nand (_11865_, _11864_, _11863_);
  nand (_11866_, _11865_, _01204_);
  nand (_11867_, _11866_, _11862_);
  nand (_11868_, _11867_, _01260_);
  nor (_11869_, _01296_, _23961_);
  nor (_11870_, _01290_, _23947_);
  nor (_11871_, _11870_, _11869_);
  nand (_11872_, _11871_, _01206_);
  nand (_11873_, _01290_, _23990_);
  nand (_11874_, _01296_, _23975_);
  nand (_11875_, _11874_, _11873_);
  nand (_11876_, _11875_, _01204_);
  nand (_11877_, _11876_, _11872_);
  nand (_11878_, _11877_, _01262_);
  nand (_11879_, _11878_, _11868_);
  nand (_11880_, _11879_, _01274_);
  nand (_11881_, _11880_, _11857_);
  nand (_11882_, _11881_, _01308_);
  nand (_11883_, _01290_, _23932_);
  nand (_11884_, _01296_, _23918_);
  nand (_11885_, _11884_, _11883_);
  nand (_11886_, _11885_, _01204_);
  nand (_11887_, _01296_, _23889_);
  nand (_11888_, _01290_, _23903_);
  nand (_11889_, _11888_, _11887_);
  nand (_11890_, _11889_, _01206_);
  nand (_11891_, _11890_, _11886_);
  nand (_11893_, _11891_, _01260_);
  nand (_11894_, _01290_, _23875_);
  nand (_11895_, _01296_, _23860_);
  nand (_11896_, _11895_, _11894_);
  nand (_11897_, _11896_, _01204_);
  nand (_11898_, _01296_, _23832_);
  nand (_11899_, _01290_, _23846_);
  nand (_11900_, _11899_, _11898_);
  nand (_11901_, _11900_, _01206_);
  nand (_11902_, _11901_, _11897_);
  nand (_11903_, _11902_, _01262_);
  nand (_11904_, _11903_, _11893_);
  nand (_11905_, _11904_, _01275_);
  nor (_11906_, _01296_, _23817_);
  nor (_11907_, _01290_, _23803_);
  nor (_11908_, _11907_, _11906_);
  nand (_11909_, _11908_, _01204_);
  nor (_11910_, _01290_, _23774_);
  nor (_11911_, _01296_, _23789_);
  nor (_11912_, _11911_, _11910_);
  nand (_11913_, _11912_, _01206_);
  nand (_11914_, _11913_, _11909_);
  nand (_11915_, _11914_, _01260_);
  nor (_11916_, _01296_, _23760_);
  nor (_11917_, _01290_, _23746_);
  nor (_11918_, _11917_, _11916_);
  nand (_11919_, _11918_, _01204_);
  nor (_11920_, _01290_, _23717_);
  nor (_11921_, _01296_, _23731_);
  nor (_11922_, _11921_, _11920_);
  nand (_11923_, _11922_, _01206_);
  nand (_11924_, _11923_, _11919_);
  nand (_11925_, _11924_, _01262_);
  nand (_11926_, _11925_, _11915_);
  nand (_11927_, _11926_, _01274_);
  nand (_11928_, _11927_, _11905_);
  nand (_11929_, _11928_, _01241_);
  nand (_11930_, _11929_, _11882_);
  nand (_11931_, _11930_, _01245_);
  nor (_11932_, _01296_, _24220_);
  nor (_11934_, _01290_, _24206_);
  nor (_11935_, _11934_, _11932_);
  nand (_11936_, _11935_, _01204_);
  nor (_11937_, _01290_, _24177_);
  nor (_11938_, _01296_, _24191_);
  nor (_11939_, _11938_, _11937_);
  nand (_11940_, _11939_, _01206_);
  nand (_11941_, _11940_, _11936_);
  nand (_11942_, _11941_, _01262_);
  nor (_11943_, _01296_, _24278_);
  nor (_11944_, _01290_, _24263_);
  nor (_11945_, _11944_, _11943_);
  nand (_11946_, _11945_, _01204_);
  nor (_11947_, _01290_, _24235_);
  nor (_11948_, _01296_, _24249_);
  nor (_11949_, _11948_, _11947_);
  nand (_11950_, _11949_, _01206_);
  nand (_11951_, _11950_, _11946_);
  nand (_11952_, _11951_, _01260_);
  nand (_11953_, _11952_, _11942_);
  nand (_11954_, _11953_, _01274_);
  nand (_11955_, _01290_, _24335_);
  nand (_11956_, _01296_, _24321_);
  nand (_11957_, _11956_, _11955_);
  nand (_11958_, _11957_, _01204_);
  nand (_11959_, _01296_, _24292_);
  nand (_11960_, _01290_, _24306_);
  nand (_11961_, _11960_, _11959_);
  nand (_11962_, _11961_, _01206_);
  nand (_11963_, _11962_, _11958_);
  nand (_11964_, _11963_, _01262_);
  nand (_11965_, _01290_, _24392_);
  nand (_11966_, _01296_, _24378_);
  nand (_11967_, _11966_, _11965_);
  nand (_11968_, _11967_, _01204_);
  nand (_11969_, _01296_, _24349_);
  nand (_11970_, _01290_, _24364_);
  nand (_11971_, _11970_, _11969_);
  nand (_11972_, _11971_, _01206_);
  nand (_11973_, _11972_, _11968_);
  nand (_11975_, _11973_, _01260_);
  nand (_11976_, _11975_, _11964_);
  nand (_11977_, _11976_, _01275_);
  nand (_11978_, _11977_, _11954_);
  nand (_11979_, _11978_, _01241_);
  nor (_11980_, _01296_, _24421_);
  nor (_11981_, _01290_, _24407_);
  nor (_11982_, _11981_, _11980_);
  nand (_11983_, _11982_, _01206_);
  nand (_11984_, _01290_, _24450_);
  nand (_11985_, _01296_, _24435_);
  nand (_11986_, _11985_, _11984_);
  nand (_11987_, _11986_, _01204_);
  nand (_11988_, _11987_, _11983_);
  nand (_11989_, _11988_, _01262_);
  nor (_11990_, _01296_, _24478_);
  nor (_11991_, _01290_, _24464_);
  nor (_11992_, _11991_, _11990_);
  nand (_11993_, _11992_, _01206_);
  nand (_11994_, _01290_, _24507_);
  nand (_11995_, _01296_, _24493_);
  nand (_11996_, _11995_, _11994_);
  nand (_11997_, _11996_, _01204_);
  nand (_11998_, _11997_, _11993_);
  nand (_11999_, _11998_, _01260_);
  nand (_12000_, _11999_, _11989_);
  nand (_12001_, _12000_, _01274_);
  nand (_12002_, _01296_, _24551_);
  nand (_12003_, _01290_, _24566_);
  nand (_12004_, _12003_, _12002_);
  nand (_12005_, _12004_, _01204_);
  nand (_12006_, _01290_, _24537_);
  nand (_12007_, _01296_, _24523_);
  nand (_12008_, _12007_, _12006_);
  nand (_12009_, _12008_, _01206_);
  nand (_12010_, _12009_, _12005_);
  nand (_12011_, _12010_, _01262_);
  nand (_12012_, _01296_, _24609_);
  nand (_12013_, _01290_, _24623_);
  nand (_12014_, _12013_, _12012_);
  nand (_12016_, _12014_, _01204_);
  nand (_12017_, _01290_, _24594_);
  nand (_12018_, _01296_, _24580_);
  nand (_12019_, _12018_, _12017_);
  nand (_12020_, _12019_, _01206_);
  nand (_12021_, _12020_, _12016_);
  nand (_12022_, _12021_, _01260_);
  nand (_12023_, _12022_, _12011_);
  nand (_12024_, _12023_, _01275_);
  nand (_12025_, _12024_, _12001_);
  nand (_12026_, _12025_, _01308_);
  nand (_12027_, _12026_, _11979_);
  nand (_12028_, _12027_, _01244_);
  nand (_12029_, _12028_, _11931_);
  nor (_12030_, _12029_, _01235_);
  nor (_12031_, _12030_, _11834_);
  nor (_12032_, _12031_, _28718_);
  nor (_12033_, _12032_, _11639_);
  nor (_12034_, _12033_, _06280_);
  nand (_12035_, _06280_, _27059_);
  nand (_12036_, _12035_, _29344_);
  nor (_15216_, _12036_, _12034_);
  nand (_12037_, _01290_, _27581_);
  nand (_12038_, _01296_, _27553_);
  nand (_12039_, _12038_, _12037_);
  nand (_12040_, _12039_, _01204_);
  nand (_12041_, _01296_, _23610_);
  nand (_12042_, _01290_, _27523_);
  nand (_12043_, _12042_, _12041_);
  nand (_12044_, _12043_, _01206_);
  nand (_12045_, _12044_, _12040_);
  nand (_12046_, _12045_, _01260_);
  nand (_12047_, _01290_, _23707_);
  nand (_12048_, _01296_, _23625_);
  nand (_12049_, _12048_, _12047_);
  nand (_12050_, _12049_, _01204_);
  nand (_12051_, _01296_, _27467_);
  nand (_12052_, _01290_, _27495_);
  nand (_12053_, _12052_, _12051_);
  nand (_12054_, _12053_, _01206_);
  nand (_12056_, _12054_, _12050_);
  nand (_12057_, _12056_, _01262_);
  nand (_12058_, _12057_, _12046_);
  nand (_12059_, _12058_, _01275_);
  nor (_12060_, _01296_, _27438_);
  nor (_12061_, _01290_, _27410_);
  nor (_12062_, _12061_, _12060_);
  nand (_12063_, _12062_, _01204_);
  nor (_12064_, _01290_, _27353_);
  nor (_12065_, _01296_, _27382_);
  nor (_12066_, _12065_, _12064_);
  nand (_12067_, _12066_, _01206_);
  nand (_12068_, _12067_, _12063_);
  nand (_12069_, _12068_, _01260_);
  nor (_12070_, _01296_, _27325_);
  nor (_12071_, _01290_, _27297_);
  nor (_12072_, _12071_, _12070_);
  nand (_12073_, _12072_, _01204_);
  nor (_12074_, _01290_, _27240_);
  nor (_12075_, _01296_, _27268_);
  nor (_12076_, _12075_, _12074_);
  nand (_12077_, _12076_, _01206_);
  nand (_12078_, _12077_, _12073_);
  nand (_12079_, _12078_, _01262_);
  nand (_12080_, _12079_, _12069_);
  nand (_12081_, _12080_, _01274_);
  nand (_12082_, _12081_, _12059_);
  nand (_12083_, _12082_, _01241_);
  nand (_12084_, _01296_, _23567_);
  nand (_12085_, _01290_, _27950_);
  nand (_12086_, _12085_, _12084_);
  nand (_12087_, _12086_, _01204_);
  nand (_12088_, _01290_, _27921_);
  nand (_12089_, _01296_, _23582_);
  nand (_12090_, _12089_, _12088_);
  nand (_12091_, _12090_, _01206_);
  nand (_12092_, _12091_, _12087_);
  nand (_12093_, _12092_, _01260_);
  nand (_12094_, _01296_, _27865_);
  nand (_12095_, _01290_, _27893_);
  nand (_12097_, _12095_, _12094_);
  nand (_12098_, _12097_, _01204_);
  nand (_12099_, _01290_, _27836_);
  nand (_12100_, _01296_, _27808_);
  nand (_12101_, _12100_, _12099_);
  nand (_12102_, _12101_, _01206_);
  nand (_12103_, _12102_, _12098_);
  nand (_12104_, _12103_, _01262_);
  nand (_12105_, _12104_, _12093_);
  nand (_12106_, _12105_, _01275_);
  nor (_12107_, _01296_, _27723_);
  nor (_12108_, _01290_, _27694_);
  nor (_12109_, _12108_, _12107_);
  nand (_12110_, _12109_, _01206_);
  nand (_12111_, _01290_, _27779_);
  nand (_12112_, _01296_, _27751_);
  nand (_12113_, _12112_, _12111_);
  nand (_12114_, _12113_, _01204_);
  nand (_12115_, _12114_, _12110_);
  nand (_12116_, _12115_, _01260_);
  nor (_12117_, _01296_, _27638_);
  nor (_12118_, _01290_, _27609_);
  nor (_12119_, _12118_, _12117_);
  nand (_12120_, _12119_, _01206_);
  nand (_12121_, _01290_, _23596_);
  nand (_12122_, _01296_, _27666_);
  nand (_12123_, _12122_, _12121_);
  nand (_12124_, _12123_, _01204_);
  nand (_12125_, _12124_, _12120_);
  nand (_12126_, _12125_, _01262_);
  nand (_12127_, _12126_, _12116_);
  nand (_12128_, _12127_, _01274_);
  nand (_12129_, _12128_, _12106_);
  nand (_12130_, _12129_, _01308_);
  nand (_12131_, _12130_, _12083_);
  nand (_12132_, _12131_, _01245_);
  nand (_12133_, _01296_, _28404_);
  nand (_12134_, _01290_, _28433_);
  nand (_12135_, _12134_, _12133_);
  nand (_12136_, _12135_, _01204_);
  nand (_12138_, _01290_, _28376_);
  nand (_12139_, _01296_, _28318_);
  nand (_12140_, _12139_, _12138_);
  nand (_12141_, _12140_, _01206_);
  nand (_12142_, _12141_, _12136_);
  nand (_12143_, _12142_, _01260_);
  nand (_12144_, _01296_, _28261_);
  nand (_12145_, _01290_, _28290_);
  nand (_12146_, _12145_, _12144_);
  nand (_12147_, _12146_, _01204_);
  nand (_12148_, _01290_, _28205_);
  nand (_12149_, _01296_, _28176_);
  nand (_12150_, _12149_, _12148_);
  nand (_12151_, _12150_, _01206_);
  nand (_12152_, _12151_, _12147_);
  nand (_12153_, _12152_, _01262_);
  nand (_12154_, _12153_, _12143_);
  nand (_12155_, _12154_, _01275_);
  nor (_12156_, _01296_, _28091_);
  nor (_12157_, _01290_, _23510_);
  nor (_12158_, _12157_, _12156_);
  nand (_12159_, _12158_, _01206_);
  nand (_12160_, _01290_, _28148_);
  nand (_12161_, _01296_, _28120_);
  nand (_12162_, _12161_, _12160_);
  nand (_12163_, _12162_, _01204_);
  nand (_12164_, _12163_, _12159_);
  nand (_12165_, _12164_, _01260_);
  nor (_12166_, _01296_, _23467_);
  nor (_12167_, _01290_, _23452_);
  nor (_12168_, _12167_, _12166_);
  nand (_12169_, _12168_, _01206_);
  nand (_12170_, _01290_, _23495_);
  nand (_12171_, _01296_, _23481_);
  nand (_12172_, _12171_, _12170_);
  nand (_12173_, _12172_, _01204_);
  nand (_12174_, _12173_, _12169_);
  nand (_12175_, _12174_, _01262_);
  nand (_12176_, _12175_, _12165_);
  nand (_12177_, _12176_, _01274_);
  nand (_12179_, _12177_, _12155_);
  nand (_12180_, _12179_, _01308_);
  nand (_12181_, _01290_, _23438_);
  nand (_12182_, _01296_, _23424_);
  nand (_12183_, _12182_, _12181_);
  nand (_12184_, _12183_, _01204_);
  nand (_12185_, _01296_, _23395_);
  nand (_12186_, _01290_, _23409_);
  nand (_12187_, _12186_, _12185_);
  nand (_12188_, _12187_, _01206_);
  nand (_12189_, _12188_, _12184_);
  nand (_12190_, _12189_, _01260_);
  nand (_12191_, _01290_, _23381_);
  nand (_12192_, _01296_, _23366_);
  nand (_12193_, _12192_, _12191_);
  nand (_12194_, _12193_, _01204_);
  nand (_12195_, _01296_, _28233_);
  nand (_12196_, _01290_, _28449_);
  nand (_12197_, _12196_, _12195_);
  nand (_12198_, _12197_, _01206_);
  nand (_12199_, _12198_, _12194_);
  nand (_12200_, _12199_, _01262_);
  nand (_12201_, _12200_, _12190_);
  nand (_12202_, _12201_, _01275_);
  nor (_12203_, _01296_, _28346_);
  nor (_12204_, _01290_, _23538_);
  nor (_12205_, _12204_, _12203_);
  nand (_12206_, _12205_, _01204_);
  nor (_12207_, _01290_, _28063_);
  nor (_12208_, _01296_, _23524_);
  nor (_12209_, _12208_, _12207_);
  nand (_12210_, _12209_, _01206_);
  nand (_12211_, _12210_, _12206_);
  nand (_12212_, _12211_, _01260_);
  nor (_12213_, _01296_, _28035_);
  nor (_12214_, _01290_, _28006_);
  nor (_12215_, _12214_, _12213_);
  nand (_12216_, _12215_, _01204_);
  nor (_12217_, _01290_, _23553_);
  nor (_12218_, _01296_, _27978_);
  nor (_12220_, _12218_, _12217_);
  nand (_12221_, _12220_, _01206_);
  nand (_12222_, _12221_, _12216_);
  nand (_12223_, _12222_, _01262_);
  nand (_12224_, _12223_, _12212_);
  nand (_12225_, _12224_, _01274_);
  nand (_12226_, _12225_, _12202_);
  nand (_12227_, _12226_, _01241_);
  nand (_12228_, _12227_, _12180_);
  nand (_12229_, _12228_, _01244_);
  nand (_12230_, _12229_, _12132_);
  nor (_12231_, _12230_, _01231_);
  nand (_12232_, _01296_, _26275_);
  nand (_12233_, _01290_, _26303_);
  nand (_12234_, _12233_, _12232_);
  nand (_12235_, _12234_, _01204_);
  nand (_12236_, _01290_, _26247_);
  nand (_12237_, _01296_, _26218_);
  nand (_12238_, _12237_, _12236_);
  nand (_12239_, _12238_, _01206_);
  nand (_12240_, _12239_, _12235_);
  nand (_12241_, _12240_, _01260_);
  nand (_12242_, _01296_, _26162_);
  nand (_12243_, _01290_, _26190_);
  nand (_12244_, _12243_, _12242_);
  nand (_12245_, _12244_, _01204_);
  nand (_12246_, _01290_, _26133_);
  nand (_12247_, _01296_, _26105_);
  nand (_12248_, _12247_, _12246_);
  nand (_12249_, _12248_, _01206_);
  nand (_12250_, _12249_, _12245_);
  nand (_12251_, _12250_, _01262_);
  nand (_12252_, _12251_, _12241_);
  nand (_12253_, _12252_, _01275_);
  nor (_12254_, _01296_, _26020_);
  nor (_12255_, _01290_, _25991_);
  nor (_12256_, _12255_, _12254_);
  nand (_12257_, _12256_, _01206_);
  nand (_12258_, _01290_, _26076_);
  nand (_12259_, _01296_, _26048_);
  nand (_12261_, _12259_, _12258_);
  nand (_12262_, _12261_, _01204_);
  nand (_12263_, _12262_, _12257_);
  nand (_12264_, _12263_, _01260_);
  nor (_12265_, _01296_, _25905_);
  nor (_12266_, _01290_, _25877_);
  nor (_12267_, _12266_, _12265_);
  nand (_12268_, _12267_, _01206_);
  nand (_12269_, _01290_, _25963_);
  nand (_12270_, _01296_, _25935_);
  nand (_12272_, _12270_, _12269_);
  nand (_12273_, _12272_, _01204_);
  nand (_12274_, _12273_, _12268_);
  nand (_12275_, _12274_, _01262_);
  nand (_12276_, _12275_, _12264_);
  nand (_12277_, _12276_, _01274_);
  nand (_12278_, _12277_, _12253_);
  nand (_12279_, _12278_, _01308_);
  nand (_12280_, _01290_, _25849_);
  nand (_12281_, _01296_, _25820_);
  nand (_12282_, _12281_, _12280_);
  nand (_12283_, _12282_, _01204_);
  nand (_12284_, _01296_, _25764_);
  nand (_12285_, _01290_, _25792_);
  nand (_12286_, _12285_, _12284_);
  nand (_12287_, _12286_, _01206_);
  nand (_12288_, _12287_, _12283_);
  nand (_12289_, _12288_, _01260_);
  nand (_12290_, _01290_, _25735_);
  nand (_12291_, _01296_, _25707_);
  nand (_12292_, _12291_, _12290_);
  nand (_12293_, _12292_, _01204_);
  nand (_12294_, _01296_, _25650_);
  nand (_12295_, _01290_, _25679_);
  nand (_12296_, _12295_, _12294_);
  nand (_12297_, _12296_, _01206_);
  nand (_12298_, _12297_, _12293_);
  nand (_12299_, _12298_, _01262_);
  nand (_12300_, _12299_, _12289_);
  nand (_12301_, _12300_, _01275_);
  nor (_12303_, _01296_, _25622_);
  nor (_12304_, _01290_, _25594_);
  nor (_12305_, _12304_, _12303_);
  nand (_12306_, _12305_, _01204_);
  nor (_12307_, _01290_, _25562_);
  nor (_12308_, _01296_, _25576_);
  nor (_12309_, _12308_, _12307_);
  nand (_12310_, _12309_, _01206_);
  nand (_12311_, _12310_, _12306_);
  nand (_12312_, _12311_, _01260_);
  nor (_12313_, _01296_, _25547_);
  nor (_12314_, _01290_, _25533_);
  nor (_12315_, _12314_, _12313_);
  nand (_12316_, _12315_, _01204_);
  nor (_12317_, _01290_, _25504_);
  nor (_12318_, _01296_, _25519_);
  nor (_12319_, _12318_, _12317_);
  nand (_12320_, _12319_, _01206_);
  nand (_12321_, _12320_, _12316_);
  nand (_12322_, _12321_, _01262_);
  nand (_12323_, _12322_, _12312_);
  nand (_12324_, _12323_, _01274_);
  nand (_12325_, _12324_, _12301_);
  nand (_12326_, _12325_, _01241_);
  nand (_12327_, _12326_, _12279_);
  nand (_12328_, _12327_, _01245_);
  nor (_12329_, _01296_, _26417_);
  nor (_12330_, _01290_, _26388_);
  nor (_12331_, _12330_, _12329_);
  nand (_12332_, _12331_, _01204_);
  nor (_12333_, _01290_, _26332_);
  nor (_12334_, _01296_, _26360_);
  nor (_12335_, _12334_, _12333_);
  nand (_12336_, _12335_, _01206_);
  nand (_12337_, _12336_, _12332_);
  nand (_12338_, _12337_, _01262_);
  nor (_12339_, _01296_, _26530_);
  nor (_12340_, _01290_, _26502_);
  nor (_12341_, _12340_, _12339_);
  nand (_12342_, _12341_, _01204_);
  nor (_12344_, _01290_, _26445_);
  nor (_12345_, _01296_, _26473_);
  nor (_12346_, _12345_, _12344_);
  nand (_12347_, _12346_, _01206_);
  nand (_12348_, _12347_, _12342_);
  nand (_12349_, _12348_, _01260_);
  nand (_12350_, _12349_, _12338_);
  nand (_12351_, _12350_, _01274_);
  nand (_12352_, _01290_, _26643_);
  nand (_12353_, _01296_, _26615_);
  nand (_12354_, _12353_, _12352_);
  nand (_12355_, _12354_, _01204_);
  nand (_12356_, _01296_, _26558_);
  nand (_12357_, _01290_, _26587_);
  nand (_12358_, _12357_, _12356_);
  nand (_12359_, _12358_, _01206_);
  nand (_12360_, _12359_, _12355_);
  nand (_12361_, _12360_, _01262_);
  nand (_12362_, _01290_, _26758_);
  nand (_12363_, _01296_, _26730_);
  nand (_12364_, _12363_, _12362_);
  nand (_12365_, _12364_, _01204_);
  nand (_12366_, _01296_, _26672_);
  nand (_12367_, _01290_, _26700_);
  nand (_12368_, _12367_, _12366_);
  nand (_12369_, _12368_, _01206_);
  nand (_12370_, _12369_, _12365_);
  nand (_12371_, _12370_, _01260_);
  nand (_12372_, _12371_, _12361_);
  nand (_12373_, _12372_, _01275_);
  nand (_12374_, _12373_, _12351_);
  nand (_12375_, _12374_, _01241_);
  nor (_12376_, _01296_, _26815_);
  nor (_12377_, _01290_, _26786_);
  nor (_12378_, _12377_, _12376_);
  nand (_12379_, _12378_, _01206_);
  nand (_12380_, _01290_, _26871_);
  nand (_12381_, _01296_, _26843_);
  nand (_12382_, _12381_, _12380_);
  nand (_12383_, _12382_, _01204_);
  nand (_12385_, _12383_, _12379_);
  nand (_12386_, _12385_, _01262_);
  nor (_12387_, _01296_, _26928_);
  nor (_12388_, _01290_, _26900_);
  nor (_12389_, _12388_, _12387_);
  nand (_12390_, _12389_, _01206_);
  nand (_12391_, _01290_, _26985_);
  nand (_12392_, _01296_, _26956_);
  nand (_12393_, _12392_, _12391_);
  nand (_12394_, _12393_, _01204_);
  nand (_12395_, _12394_, _12390_);
  nand (_12396_, _12395_, _01260_);
  nand (_12397_, _12396_, _12386_);
  nand (_12398_, _12397_, _01274_);
  nand (_12399_, _01296_, _27070_);
  nand (_12400_, _01290_, _27098_);
  nand (_12401_, _12400_, _12399_);
  nand (_12402_, _12401_, _01204_);
  nand (_12403_, _01290_, _27041_);
  nand (_12404_, _01296_, _27013_);
  nand (_12405_, _12404_, _12403_);
  nand (_12406_, _12405_, _01206_);
  nand (_12407_, _12406_, _12402_);
  nand (_12408_, _12407_, _01262_);
  nand (_12409_, _01296_, _27183_);
  nand (_12410_, _01290_, _27211_);
  nand (_12411_, _12410_, _12409_);
  nand (_12412_, _12411_, _01204_);
  nand (_12413_, _01290_, _27155_);
  nand (_12414_, _01296_, _27126_);
  nand (_12415_, _12414_, _12413_);
  nand (_12416_, _12415_, _01206_);
  nand (_12417_, _12416_, _12412_);
  nand (_12418_, _12417_, _01260_);
  nand (_12419_, _12418_, _12408_);
  nand (_12420_, _12419_, _01275_);
  nand (_12421_, _12420_, _12398_);
  nand (_12422_, _12421_, _01308_);
  nand (_12423_, _12422_, _12375_);
  nand (_12424_, _12423_, _01244_);
  nand (_12426_, _12424_, _12328_);
  nor (_12427_, _12426_, _01235_);
  nor (_12428_, _12427_, _12231_);
  nor (_12429_, _12428_, _28717_);
  nand (_12430_, _01290_, _24857_);
  nand (_12431_, _01296_, _24842_);
  nand (_12432_, _12431_, _12430_);
  nand (_12433_, _12432_, _01204_);
  nand (_12434_, _01296_, _24814_);
  nand (_12435_, _01290_, _24828_);
  nand (_12436_, _12435_, _12434_);
  nand (_12437_, _12436_, _01206_);
  nand (_12438_, _12437_, _12433_);
  nand (_12439_, _12438_, _01260_);
  nand (_12440_, _01290_, _24799_);
  nand (_12441_, _01296_, _24785_);
  nand (_12442_, _12441_, _12440_);
  nand (_12443_, _12442_, _01204_);
  nand (_12444_, _01296_, _24756_);
  nand (_12445_, _01290_, _24771_);
  nand (_12446_, _12445_, _12444_);
  nand (_12447_, _12446_, _01206_);
  nand (_12448_, _12447_, _12443_);
  nand (_12449_, _12448_, _01262_);
  nand (_12450_, _12449_, _12439_);
  nand (_12451_, _12450_, _01275_);
  nor (_12452_, _01296_, _24742_);
  nor (_12453_, _01290_, _24728_);
  nor (_12454_, _12453_, _12452_);
  nand (_12455_, _12454_, _01204_);
  nor (_12456_, _01290_, _24699_);
  nor (_12457_, _01296_, _24713_);
  nor (_12458_, _12457_, _12456_);
  nand (_12459_, _12458_, _01206_);
  nand (_12460_, _12459_, _12455_);
  nand (_12461_, _12460_, _01260_);
  nor (_12462_, _01296_, _24684_);
  nor (_12463_, _01290_, _24670_);
  nor (_12464_, _12463_, _12462_);
  nand (_12465_, _12464_, _01204_);
  nor (_12467_, _01290_, _24641_);
  nor (_12468_, _01296_, _24656_);
  nor (_12469_, _12468_, _12467_);
  nand (_12470_, _12469_, _01206_);
  nand (_12471_, _12470_, _12465_);
  nand (_12472_, _12471_, _01262_);
  nand (_12473_, _12472_, _12461_);
  nand (_12474_, _12473_, _01274_);
  nand (_12475_, _12474_, _12451_);
  nand (_12476_, _12475_, _01241_);
  nand (_12477_, _01296_, _25073_);
  nand (_12478_, _01290_, _25087_);
  nand (_12479_, _12478_, _12477_);
  nand (_12480_, _12479_, _01204_);
  nand (_12481_, _01290_, _25059_);
  nand (_12482_, _01296_, _25044_);
  nand (_12483_, _12482_, _12481_);
  nand (_12484_, _12483_, _01206_);
  nand (_12485_, _12484_, _12480_);
  nand (_12486_, _12485_, _01260_);
  nand (_12487_, _01296_, _25016_);
  nand (_12488_, _01290_, _25030_);
  nand (_12489_, _12488_, _12487_);
  nand (_12490_, _12489_, _01204_);
  nand (_12491_, _01290_, _25001_);
  nand (_12492_, _01296_, _24987_);
  nand (_12493_, _12492_, _12491_);
  nand (_12494_, _12493_, _01206_);
  nand (_12495_, _12494_, _12490_);
  nand (_12496_, _12495_, _01262_);
  nand (_12497_, _12496_, _12486_);
  nand (_12498_, _12497_, _01275_);
  nor (_12499_, _01296_, _24944_);
  nor (_12500_, _01290_, _24928_);
  nor (_12501_, _12500_, _12499_);
  nand (_12502_, _12501_, _01206_);
  nand (_12503_, _01290_, _24972_);
  nand (_12504_, _01296_, _24958_);
  nand (_12505_, _12504_, _12503_);
  nand (_12506_, _12505_, _01204_);
  nand (_12508_, _12506_, _12502_);
  nand (_12509_, _12508_, _01260_);
  nor (_12510_, _01296_, _24885_);
  nor (_12511_, _01290_, _24871_);
  nor (_12512_, _12511_, _12510_);
  nand (_12513_, _12512_, _01206_);
  nand (_12514_, _01290_, _24914_);
  nand (_12515_, _01296_, _24900_);
  nand (_12516_, _12515_, _12514_);
  nand (_12517_, _12516_, _01204_);
  nand (_12518_, _12517_, _12513_);
  nand (_12519_, _12518_, _01262_);
  nand (_12520_, _12519_, _12509_);
  nand (_12521_, _12520_, _01274_);
  nand (_12522_, _12521_, _12498_);
  nand (_12523_, _12522_, _01308_);
  nand (_12524_, _12523_, _12476_);
  nand (_12525_, _12524_, _01245_);
  nand (_12526_, _01296_, _25476_);
  nand (_12527_, _01290_, _25490_);
  nand (_12528_, _12527_, _12526_);
  nand (_12529_, _12528_, _01204_);
  nand (_12530_, _01290_, _25461_);
  nand (_12531_, _01296_, _25447_);
  nand (_12532_, _12531_, _12530_);
  nand (_12533_, _12532_, _01206_);
  nand (_12534_, _12533_, _12529_);
  nand (_12535_, _12534_, _01260_);
  nand (_12536_, _01296_, _25418_);
  nand (_12537_, _01290_, _25433_);
  nand (_12538_, _12537_, _12536_);
  nand (_12539_, _12538_, _01204_);
  nand (_12540_, _01290_, _25404_);
  nand (_12541_, _01296_, _25390_);
  nand (_12542_, _12541_, _12540_);
  nand (_12543_, _12542_, _01206_);
  nand (_12544_, _12543_, _12539_);
  nand (_12545_, _12544_, _01262_);
  nand (_12546_, _12545_, _12535_);
  nand (_12547_, _12546_, _01275_);
  nor (_12549_, _01296_, _25347_);
  nor (_12550_, _01290_, _25331_);
  nor (_12551_, _12550_, _12549_);
  nand (_12552_, _12551_, _01206_);
  nand (_12553_, _01290_, _25375_);
  nand (_12554_, _01296_, _25361_);
  nand (_12555_, _12554_, _12553_);
  nand (_12556_, _12555_, _01204_);
  nand (_12557_, _12556_, _12552_);
  nand (_12558_, _12557_, _01260_);
  nor (_12559_, _01296_, _25288_);
  nor (_12560_, _01290_, _25274_);
  nor (_12561_, _12560_, _12559_);
  nand (_12562_, _12561_, _01206_);
  nand (_12563_, _01290_, _25317_);
  nand (_12564_, _01296_, _25303_);
  nand (_12565_, _12564_, _12563_);
  nand (_12566_, _12565_, _01204_);
  nand (_12567_, _12566_, _12562_);
  nand (_12568_, _12567_, _01262_);
  nand (_12569_, _12568_, _12558_);
  nand (_12570_, _12569_, _01274_);
  nand (_12571_, _12570_, _12547_);
  nand (_12572_, _12571_, _01308_);
  nand (_12573_, _01290_, _25259_);
  nand (_12574_, _01296_, _25245_);
  nand (_12575_, _12574_, _12573_);
  nand (_12576_, _12575_, _01204_);
  nand (_12577_, _01296_, _25216_);
  nand (_12578_, _01290_, _25231_);
  nand (_12579_, _12578_, _12577_);
  nand (_12580_, _12579_, _01206_);
  nand (_12581_, _12580_, _12576_);
  nand (_12582_, _12581_, _01260_);
  nand (_12583_, _01290_, _25202_);
  nand (_12584_, _01296_, _25188_);
  nand (_12585_, _12584_, _12583_);
  nand (_12586_, _12585_, _01204_);
  nand (_12587_, _01296_, _25159_);
  nand (_12588_, _01290_, _25173_);
  nand (_12590_, _12588_, _12587_);
  nand (_12591_, _12590_, _01206_);
  nand (_12592_, _12591_, _12586_);
  nand (_12593_, _12592_, _01262_);
  nand (_12594_, _12593_, _12582_);
  nand (_12595_, _12594_, _01275_);
  nor (_12596_, _01296_, _25145_);
  nor (_12597_, _01290_, _25130_);
  nor (_12598_, _12597_, _12596_);
  nand (_12599_, _12598_, _01204_);
  nor (_12600_, _01290_, _23682_);
  nor (_12601_, _01296_, _25116_);
  nor (_12602_, _12601_, _12600_);
  nand (_12603_, _12602_, _01206_);
  nand (_12604_, _12603_, _12599_);
  nand (_12605_, _12604_, _01260_);
  nor (_12606_, _01296_, _23653_);
  nor (_12607_, _01290_, _23639_);
  nor (_12608_, _12607_, _12606_);
  nand (_12609_, _12608_, _01204_);
  nor (_12610_, _01290_, _25102_);
  nor (_12611_, _01296_, _23668_);
  nor (_12612_, _12611_, _12610_);
  nand (_12613_, _12612_, _01206_);
  nand (_12614_, _12613_, _12609_);
  nand (_12615_, _12614_, _01262_);
  nand (_12616_, _12615_, _12605_);
  nand (_12617_, _12616_, _01274_);
  nand (_12618_, _12617_, _12595_);
  nand (_12619_, _12618_, _01241_);
  nand (_12620_, _12619_, _12572_);
  nand (_12621_, _12620_, _01244_);
  nand (_12622_, _12621_, _12525_);
  nor (_12623_, _12622_, _01231_);
  nand (_12624_, _01296_, _24153_);
  nand (_12625_, _01290_, _24167_);
  nand (_12626_, _12625_, _12624_);
  nand (_12627_, _12626_, _01204_);
  nand (_12628_, _01290_, _24138_);
  nand (_12629_, _01296_, _24124_);
  nand (_12631_, _12629_, _12628_);
  nand (_12632_, _12631_, _01206_);
  nand (_12633_, _12632_, _12627_);
  nand (_12634_, _12633_, _01260_);
  nand (_12635_, _01296_, _24094_);
  nand (_12636_, _01290_, _24108_);
  nand (_12637_, _12636_, _12635_);
  nand (_12638_, _12637_, _01204_);
  nand (_12639_, _01290_, _24080_);
  nand (_12640_, _01296_, _24065_);
  nand (_12642_, _12640_, _12639_);
  nand (_12643_, _12642_, _01206_);
  nand (_12644_, _12643_, _12638_);
  nand (_12645_, _12644_, _01262_);
  nand (_12646_, _12645_, _12634_);
  nand (_12647_, _12646_, _01275_);
  nor (_12648_, _01296_, _24022_);
  nor (_12649_, _01290_, _24008_);
  nor (_12650_, _12649_, _12648_);
  nand (_12651_, _12650_, _01206_);
  nand (_12652_, _01290_, _24051_);
  nand (_12653_, _01296_, _24037_);
  nand (_12654_, _12653_, _12652_);
  nand (_12655_, _12654_, _01204_);
  nand (_12656_, _12655_, _12651_);
  nand (_12657_, _12656_, _01260_);
  nor (_12658_, _01296_, _23965_);
  nor (_12659_, _01290_, _23951_);
  nor (_12660_, _12659_, _12658_);
  nand (_12661_, _12660_, _01206_);
  nand (_12662_, _01290_, _23994_);
  nand (_12663_, _01296_, _23979_);
  nand (_12664_, _12663_, _12662_);
  nand (_12665_, _12664_, _01204_);
  nand (_12666_, _12665_, _12661_);
  nand (_12667_, _12666_, _01262_);
  nand (_12668_, _12667_, _12657_);
  nand (_12669_, _12668_, _01274_);
  nand (_12670_, _12669_, _12647_);
  nand (_12671_, _12670_, _01308_);
  nand (_12673_, _01290_, _23936_);
  nand (_12674_, _01296_, _23922_);
  nand (_12675_, _12674_, _12673_);
  nand (_12676_, _12675_, _01204_);
  nand (_12677_, _01296_, _23893_);
  nand (_12678_, _01290_, _23908_);
  nand (_12679_, _12678_, _12677_);
  nand (_12680_, _12679_, _01206_);
  nand (_12681_, _12680_, _12676_);
  nand (_12682_, _12681_, _01260_);
  nand (_12685_, _01290_, _23879_);
  nand (_12686_, _01296_, _23865_);
  nand (_12687_, _12686_, _12685_);
  nand (_12688_, _12687_, _01204_);
  nand (_12689_, _01296_, _23836_);
  nand (_12690_, _01290_, _23850_);
  nand (_12691_, _12690_, _12689_);
  nand (_12692_, _12691_, _01206_);
  nand (_12693_, _12692_, _12688_);
  nand (_12694_, _12693_, _01262_);
  nand (_12695_, _12694_, _12682_);
  nand (_12696_, _12695_, _01275_);
  nor (_12697_, _01296_, _23821_);
  nor (_12698_, _01290_, _23807_);
  nor (_12699_, _12698_, _12697_);
  nand (_12700_, _12699_, _01204_);
  nor (_12701_, _01290_, _23778_);
  nor (_12702_, _01296_, _23793_);
  nor (_12703_, _12702_, _12701_);
  nand (_12704_, _12703_, _01206_);
  nand (_12705_, _12704_, _12700_);
  nand (_12706_, _12705_, _01260_);
  nor (_12707_, _01296_, _23764_);
  nor (_12708_, _01290_, _23750_);
  nor (_12709_, _12708_, _12707_);
  nand (_12710_, _12709_, _01204_);
  nor (_12711_, _01290_, _23721_);
  nor (_12712_, _01296_, _23735_);
  nor (_12713_, _12712_, _12711_);
  nand (_12714_, _12713_, _01206_);
  nand (_12716_, _12714_, _12710_);
  nand (_12717_, _12716_, _01262_);
  nand (_12718_, _12717_, _12706_);
  nand (_12719_, _12718_, _01274_);
  nand (_12720_, _12719_, _12696_);
  nand (_12721_, _12720_, _01241_);
  nand (_12722_, _12721_, _12671_);
  nand (_12723_, _12722_, _01245_);
  nor (_12724_, _01296_, _24224_);
  nor (_12725_, _01290_, _24210_);
  nor (_12726_, _12725_, _12724_);
  nand (_12727_, _12726_, _01204_);
  nor (_12728_, _01290_, _24181_);
  nor (_12729_, _01296_, _24196_);
  nor (_12730_, _12729_, _12728_);
  nand (_12731_, _12730_, _01206_);
  nand (_12732_, _12731_, _12727_);
  nand (_12733_, _12732_, _01262_);
  nor (_12734_, _01296_, _24282_);
  nor (_12735_, _01290_, _24267_);
  nor (_12736_, _12735_, _12734_);
  nand (_12737_, _12736_, _01204_);
  nor (_12738_, _01290_, _24239_);
  nor (_12739_, _01296_, _24253_);
  nor (_12740_, _12739_, _12738_);
  nand (_12741_, _12740_, _01206_);
  nand (_12742_, _12741_, _12737_);
  nand (_12743_, _12742_, _01260_);
  nand (_12744_, _12743_, _12733_);
  nand (_12745_, _12744_, _01274_);
  nand (_12746_, _01290_, _24339_);
  nand (_12747_, _01296_, _24325_);
  nand (_12748_, _12747_, _12746_);
  nand (_12749_, _12748_, _01204_);
  nand (_12750_, _01296_, _24296_);
  nand (_12751_, _01290_, _24310_);
  nand (_12752_, _12751_, _12750_);
  nand (_12753_, _12752_, _01206_);
  nand (_12754_, _12753_, _12749_);
  nand (_12755_, _12754_, _01262_);
  nand (_12757_, _01290_, _24396_);
  nand (_12758_, _01296_, _24382_);
  nand (_12759_, _12758_, _12757_);
  nand (_12760_, _12759_, _01204_);
  nand (_12761_, _01296_, _24353_);
  nand (_12762_, _01290_, _24368_);
  nand (_12763_, _12762_, _12761_);
  nand (_12764_, _12763_, _01206_);
  nand (_12765_, _12764_, _12760_);
  nand (_12766_, _12765_, _01260_);
  nand (_12767_, _12766_, _12755_);
  nand (_12768_, _12767_, _01275_);
  nand (_12769_, _12768_, _12745_);
  nand (_12770_, _12769_, _01241_);
  nor (_12771_, _01296_, _24425_);
  nor (_12772_, _01290_, _24411_);
  nor (_12773_, _12772_, _12771_);
  nand (_12774_, _12773_, _01206_);
  nand (_12775_, _01290_, _24454_);
  nand (_12776_, _01296_, _24440_);
  nand (_12777_, _12776_, _12775_);
  nand (_12778_, _12777_, _01204_);
  nand (_12779_, _12778_, _12774_);
  nand (_12780_, _12779_, _01262_);
  nor (_12781_, _01296_, _24483_);
  nor (_12782_, _01290_, _24468_);
  nor (_12783_, _12782_, _12781_);
  nand (_12784_, _12783_, _01206_);
  nand (_12785_, _01290_, _24511_);
  nand (_12786_, _01296_, _24497_);
  nand (_12787_, _12786_, _12785_);
  nand (_12788_, _12787_, _01204_);
  nand (_12789_, _12788_, _12784_);
  nand (_12790_, _12789_, _01260_);
  nand (_12791_, _12790_, _12780_);
  nand (_12792_, _12791_, _01274_);
  nand (_12793_, _01296_, _24555_);
  nand (_12794_, _01290_, _24570_);
  nand (_12795_, _12794_, _12793_);
  nand (_12796_, _12795_, _01204_);
  nand (_12798_, _01290_, _24541_);
  nand (_12799_, _01296_, _24527_);
  nand (_12800_, _12799_, _12798_);
  nand (_12801_, _12800_, _01206_);
  nand (_12802_, _12801_, _12796_);
  nand (_12803_, _12802_, _01262_);
  nand (_12804_, _01296_, _24613_);
  nand (_12805_, _01290_, _24627_);
  nand (_12806_, _12805_, _12804_);
  nand (_12807_, _12806_, _01204_);
  nand (_12808_, _01290_, _24598_);
  nand (_12809_, _01296_, _24584_);
  nand (_12810_, _12809_, _12808_);
  nand (_12811_, _12810_, _01206_);
  nand (_12812_, _12811_, _12807_);
  nand (_12813_, _12812_, _01260_);
  nand (_12814_, _12813_, _12803_);
  nand (_12815_, _12814_, _01275_);
  nand (_12816_, _12815_, _12792_);
  nand (_12817_, _12816_, _01308_);
  nand (_12818_, _12817_, _12770_);
  nand (_12819_, _12818_, _01244_);
  nand (_12820_, _12819_, _12723_);
  nor (_12821_, _12820_, _01235_);
  nor (_12822_, _12821_, _12623_);
  nor (_12823_, _12822_, _28718_);
  nor (_12824_, _12823_, _12429_);
  nor (_12825_, _12824_, _06280_);
  not (_12826_, _23691_);
  nand (_12827_, _06280_, _12826_);
  nand (_12828_, _12827_, _29344_);
  nor (_15244_, _12828_, _12825_);
  nand (_12829_, _01290_, _27577_);
  nand (_12830_, _01296_, _27549_);
  nand (_12831_, _12830_, _12829_);
  nand (_12832_, _12831_, _01204_);
  nand (_12833_, _01296_, _23608_);
  nand (_12834_, _01290_, _27519_);
  nand (_12835_, _12834_, _12833_);
  nand (_12836_, _12835_, _01206_);
  nand (_12838_, _12836_, _12832_);
  nand (_12839_, _12838_, _01260_);
  nand (_12840_, _01290_, _23705_);
  nand (_12841_, _01296_, _23623_);
  nand (_12842_, _12841_, _12840_);
  nand (_12843_, _12842_, _01204_);
  nand (_12844_, _01296_, _27463_);
  nand (_12845_, _01290_, _27491_);
  nand (_12846_, _12845_, _12844_);
  nand (_12847_, _12846_, _01206_);
  nand (_12848_, _12847_, _12843_);
  nand (_12849_, _12848_, _01262_);
  nand (_12850_, _12849_, _12839_);
  nand (_12851_, _12850_, _01275_);
  nor (_12852_, _01296_, _27434_);
  nor (_12853_, _01290_, _27406_);
  nor (_12854_, _12853_, _12852_);
  nand (_12855_, _12854_, _01204_);
  nor (_12856_, _01290_, _27349_);
  nor (_12857_, _01296_, _27378_);
  nor (_12858_, _12857_, _12856_);
  nand (_12859_, _12858_, _01206_);
  nand (_12860_, _12859_, _12855_);
  nand (_12861_, _12860_, _01260_);
  nor (_12862_, _01296_, _27321_);
  nor (_12863_, _01290_, _27292_);
  nor (_12864_, _12863_, _12862_);
  nand (_12865_, _12864_, _01204_);
  nor (_12866_, _01290_, _27236_);
  nor (_12867_, _01296_, _27264_);
  nor (_12868_, _12867_, _12866_);
  nand (_12869_, _12868_, _01206_);
  nand (_12870_, _12869_, _12865_);
  nand (_12871_, _12870_, _01262_);
  nand (_12872_, _12871_, _12861_);
  nand (_12873_, _12872_, _01274_);
  nand (_12874_, _12873_, _12851_);
  nand (_12875_, _12874_, _01241_);
  nand (_12876_, _01296_, _23565_);
  nand (_12877_, _01290_, _27946_);
  nand (_12879_, _12877_, _12876_);
  nand (_12880_, _12879_, _01204_);
  nand (_12881_, _01290_, _27917_);
  nand (_12882_, _01296_, _23579_);
  nand (_12883_, _12882_, _12881_);
  nand (_12884_, _12883_, _01206_);
  nand (_12885_, _12884_, _12880_);
  nand (_12886_, _12885_, _01260_);
  nand (_12887_, _01296_, _27860_);
  nand (_12888_, _01290_, _27889_);
  nand (_12889_, _12888_, _12887_);
  nand (_12890_, _12889_, _01204_);
  nand (_12891_, _01290_, _27832_);
  nand (_12892_, _01296_, _27804_);
  nand (_12893_, _12892_, _12891_);
  nand (_12894_, _12893_, _01206_);
  nand (_12895_, _12894_, _12890_);
  nand (_12896_, _12895_, _01262_);
  nand (_12897_, _12896_, _12886_);
  nand (_12898_, _12897_, _01275_);
  nor (_12899_, _01296_, _27719_);
  nor (_12900_, _01290_, _27690_);
  nor (_12901_, _12900_, _12899_);
  nand (_12902_, _12901_, _01206_);
  nand (_12903_, _01290_, _27775_);
  nand (_12904_, _01296_, _27747_);
  nand (_12905_, _12904_, _12903_);
  nand (_12906_, _12905_, _01204_);
  nand (_12907_, _12906_, _12902_);
  nand (_12908_, _12907_, _01260_);
  nor (_12909_, _01296_, _27634_);
  nor (_12910_, _01290_, _27605_);
  nor (_12911_, _12910_, _12909_);
  nand (_12912_, _12911_, _01206_);
  nand (_12913_, _01290_, _23594_);
  nand (_12914_, _01296_, _27662_);
  nand (_12915_, _12914_, _12913_);
  nand (_12916_, _12915_, _01204_);
  nand (_12917_, _12916_, _12912_);
  nand (_12918_, _12917_, _01262_);
  nand (_12920_, _12918_, _12908_);
  nand (_12921_, _12920_, _01274_);
  nand (_12922_, _12921_, _12898_);
  nand (_12923_, _12922_, _01308_);
  nand (_12924_, _12923_, _12875_);
  nand (_12925_, _12924_, _01245_);
  nand (_12926_, _01296_, _28400_);
  nand (_12927_, _01290_, _28428_);
  nand (_12928_, _12927_, _12926_);
  nand (_12929_, _12928_, _01204_);
  nand (_12930_, _01290_, _28372_);
  nand (_12931_, _01296_, _28314_);
  nand (_12932_, _12931_, _12930_);
  nand (_12933_, _12932_, _01206_);
  nand (_12934_, _12933_, _12929_);
  nand (_12935_, _12934_, _01260_);
  nand (_12936_, _01296_, _28257_);
  nand (_12937_, _01290_, _28286_);
  nand (_12938_, _12937_, _12936_);
  nand (_12939_, _12938_, _01204_);
  nand (_12940_, _01290_, _28201_);
  nand (_12941_, _01296_, _28172_);
  nand (_12942_, _12941_, _12940_);
  nand (_12943_, _12942_, _01206_);
  nand (_12944_, _12943_, _12939_);
  nand (_12945_, _12944_, _01262_);
  nand (_12946_, _12945_, _12935_);
  nand (_12947_, _12946_, _01275_);
  nor (_12948_, _01296_, _28087_);
  nor (_12949_, _01290_, _23508_);
  nor (_12950_, _12949_, _12948_);
  nand (_12951_, _12950_, _01206_);
  nand (_12952_, _01290_, _28144_);
  nand (_12953_, _01296_, _28116_);
  nand (_12954_, _12953_, _12952_);
  nand (_12955_, _12954_, _01204_);
  nand (_12956_, _12955_, _12951_);
  nand (_12957_, _12956_, _01260_);
  nor (_12958_, _01296_, _23465_);
  nor (_12959_, _01290_, _23450_);
  nor (_12961_, _12959_, _12958_);
  nand (_12962_, _12961_, _01206_);
  nand (_12963_, _01290_, _23493_);
  nand (_12964_, _01296_, _23479_);
  nand (_12965_, _12964_, _12963_);
  nand (_12966_, _12965_, _01204_);
  nand (_12967_, _12966_, _12962_);
  nand (_12968_, _12967_, _01262_);
  nand (_12969_, _12968_, _12957_);
  nand (_12970_, _12969_, _01274_);
  nand (_12971_, _12970_, _12947_);
  nand (_12972_, _12971_, _01308_);
  nand (_12973_, _01290_, _23436_);
  nand (_12974_, _01296_, _23422_);
  nand (_12975_, _12974_, _12973_);
  nand (_12976_, _12975_, _01204_);
  nand (_12977_, _01296_, _23393_);
  nand (_12978_, _01290_, _23407_);
  nand (_12979_, _12978_, _12977_);
  nand (_12980_, _12979_, _01206_);
  nand (_12981_, _12980_, _12976_);
  nand (_12982_, _12981_, _01260_);
  nand (_12983_, _01290_, _23379_);
  nand (_12984_, _01296_, _23364_);
  nand (_12985_, _12984_, _12983_);
  nand (_12986_, _12985_, _01204_);
  nand (_12987_, _01296_, _28229_);
  nand (_12988_, _01290_, _28437_);
  nand (_12989_, _12988_, _12987_);
  nand (_12990_, _12989_, _01206_);
  nand (_12991_, _12990_, _12986_);
  nand (_12992_, _12991_, _01262_);
  nand (_12993_, _12992_, _12982_);
  nand (_12994_, _12993_, _01275_);
  nor (_12995_, _01296_, _28342_);
  nor (_12996_, _01290_, _23536_);
  nor (_12997_, _12996_, _12995_);
  nand (_12998_, _12997_, _01204_);
  nor (_12999_, _01290_, _28059_);
  nor (_13000_, _01296_, _23522_);
  nor (_13002_, _13000_, _12999_);
  nand (_13003_, _13002_, _01206_);
  nand (_13004_, _13003_, _12998_);
  nand (_13005_, _13004_, _01260_);
  nor (_13006_, _01296_, _28031_);
  nor (_13007_, _01290_, _28002_);
  nor (_13008_, _13007_, _13006_);
  nand (_13009_, _13008_, _01204_);
  nor (_13010_, _01290_, _23551_);
  nor (_13011_, _01296_, _27974_);
  nor (_13012_, _13011_, _13010_);
  nand (_13013_, _13012_, _01206_);
  nand (_13014_, _13013_, _13009_);
  nand (_13015_, _13014_, _01262_);
  nand (_13016_, _13015_, _13005_);
  nand (_13017_, _13016_, _01274_);
  nand (_13018_, _13017_, _12994_);
  nand (_13019_, _13018_, _01241_);
  nand (_13020_, _13019_, _12972_);
  nand (_13021_, _13020_, _01244_);
  nand (_13022_, _13021_, _12925_);
  nor (_13023_, _13022_, _01231_);
  nand (_13024_, _01296_, _26271_);
  nand (_13025_, _01290_, _26299_);
  nand (_13026_, _13025_, _13024_);
  nand (_13027_, _13026_, _01204_);
  nand (_13028_, _01290_, _26243_);
  nand (_13029_, _01296_, _26214_);
  nand (_13030_, _13029_, _13028_);
  nand (_13031_, _13030_, _01206_);
  nand (_13032_, _13031_, _13027_);
  nand (_13033_, _13032_, _01260_);
  nand (_13034_, _01296_, _26157_);
  nand (_13035_, _01290_, _26186_);
  nand (_13036_, _13035_, _13034_);
  nand (_13037_, _13036_, _01204_);
  nand (_13038_, _01290_, _26129_);
  nand (_13039_, _01296_, _26101_);
  nand (_13040_, _13039_, _13038_);
  nand (_13041_, _13040_, _01206_);
  nand (_13043_, _13041_, _13037_);
  nand (_13044_, _13043_, _01262_);
  nand (_13045_, _13044_, _13033_);
  nand (_13046_, _13045_, _01275_);
  nor (_13047_, _01296_, _26016_);
  nor (_13048_, _01290_, _25987_);
  nor (_13049_, _13048_, _13047_);
  nand (_13050_, _13049_, _01206_);
  nand (_13051_, _01290_, _26072_);
  nand (_13052_, _01296_, _26044_);
  nand (_13053_, _13052_, _13051_);
  nand (_13054_, _13053_, _01204_);
  nand (_13055_, _13054_, _13050_);
  nand (_13056_, _13055_, _01260_);
  nor (_13057_, _01296_, _25901_);
  nor (_13058_, _01290_, _25873_);
  nor (_13059_, _13058_, _13057_);
  nand (_13060_, _13059_, _01206_);
  nand (_13061_, _01290_, _25959_);
  nand (_13062_, _01296_, _25931_);
  nand (_13063_, _13062_, _13061_);
  nand (_13064_, _13063_, _01204_);
  nand (_13065_, _13064_, _13060_);
  nand (_13066_, _13065_, _01262_);
  nand (_13067_, _13066_, _13056_);
  nand (_13068_, _13067_, _01274_);
  nand (_13069_, _13068_, _13046_);
  nand (_13070_, _13069_, _01308_);
  nand (_13071_, _01290_, _25845_);
  nand (_13072_, _01296_, _25816_);
  nand (_13073_, _13072_, _13071_);
  nand (_13074_, _13073_, _01204_);
  nand (_13075_, _01296_, _25760_);
  nand (_13076_, _01290_, _25788_);
  nand (_13077_, _13076_, _13075_);
  nand (_13078_, _13077_, _01206_);
  nand (_13079_, _13078_, _13074_);
  nand (_13080_, _13079_, _01260_);
  nand (_13081_, _01290_, _25731_);
  nand (_13082_, _01296_, _25703_);
  nand (_13084_, _13082_, _13081_);
  nand (_13085_, _13084_, _01204_);
  nand (_13086_, _01296_, _25646_);
  nand (_13087_, _01290_, _25675_);
  nand (_13088_, _13087_, _13086_);
  nand (_13089_, _13088_, _01206_);
  nand (_13090_, _13089_, _13085_);
  nand (_13091_, _13090_, _01262_);
  nand (_13092_, _13091_, _13080_);
  nand (_13093_, _13092_, _01275_);
  nor (_13095_, _01296_, _25618_);
  nor (_13096_, _01290_, _25589_);
  nor (_13097_, _13096_, _13095_);
  nand (_13098_, _13097_, _01204_);
  nor (_13099_, _01290_, _25560_);
  nor (_13100_, _01296_, _25574_);
  nor (_13101_, _13100_, _13099_);
  nand (_13102_, _13101_, _01206_);
  nand (_13103_, _13102_, _13098_);
  nand (_13104_, _13103_, _01260_);
  nor (_13105_, _01296_, _25545_);
  nor (_13106_, _01290_, _25531_);
  nor (_13107_, _13106_, _13105_);
  nand (_13108_, _13107_, _01204_);
  nor (_13109_, _01290_, _25502_);
  nor (_13110_, _01296_, _25517_);
  nor (_13111_, _13110_, _13109_);
  nand (_13112_, _13111_, _01206_);
  nand (_13113_, _13112_, _13108_);
  nand (_13114_, _13113_, _01262_);
  nand (_13115_, _13114_, _13104_);
  nand (_13116_, _13115_, _01274_);
  nand (_13117_, _13116_, _13093_);
  nand (_13118_, _13117_, _01241_);
  nand (_13119_, _13118_, _13070_);
  nand (_13120_, _13119_, _01245_);
  nor (_13121_, _01296_, _26413_);
  nor (_13122_, _01290_, _26384_);
  nor (_13123_, _13122_, _13121_);
  nand (_13124_, _13123_, _01204_);
  nor (_13126_, _01290_, _26328_);
  nor (_13127_, _01296_, _26356_);
  nor (_13128_, _13127_, _13126_);
  nand (_13129_, _13128_, _01206_);
  nand (_13130_, _13129_, _13124_);
  nand (_13131_, _13130_, _01262_);
  nor (_13132_, _01296_, _26526_);
  nor (_13133_, _01290_, _26498_);
  nor (_13134_, _13133_, _13132_);
  nand (_13135_, _13134_, _01204_);
  nor (_13136_, _01290_, _26441_);
  nor (_13137_, _01296_, _26469_);
  nor (_13138_, _13137_, _13136_);
  nand (_13139_, _13138_, _01206_);
  nand (_13140_, _13139_, _13135_);
  nand (_13141_, _13140_, _01260_);
  nand (_13142_, _13141_, _13131_);
  nand (_13143_, _13142_, _01274_);
  nand (_13144_, _01290_, _26639_);
  nand (_13145_, _01296_, _26611_);
  nand (_13146_, _13145_, _13144_);
  nand (_13147_, _13146_, _01204_);
  nand (_13148_, _01296_, _26554_);
  nand (_13149_, _01290_, _26583_);
  nand (_13150_, _13149_, _13148_);
  nand (_13151_, _13150_, _01206_);
  nand (_13152_, _13151_, _13147_);
  nand (_13153_, _13152_, _01262_);
  nand (_13154_, _01290_, _26754_);
  nand (_13155_, _01296_, _26724_);
  nand (_13156_, _13155_, _13154_);
  nand (_13157_, _13156_, _01204_);
  nand (_13158_, _01296_, _26668_);
  nand (_13159_, _01290_, _26696_);
  nand (_13160_, _13159_, _13158_);
  nand (_13161_, _13160_, _01206_);
  nand (_13162_, _13161_, _13157_);
  nand (_13163_, _13162_, _01260_);
  nand (_13164_, _13163_, _13153_);
  nand (_13165_, _13164_, _01275_);
  nand (_13167_, _13165_, _13143_);
  nand (_13168_, _13167_, _01241_);
  nor (_13169_, _01296_, _26811_);
  nor (_13170_, _01290_, _26782_);
  nor (_13171_, _13170_, _13169_);
  nand (_13172_, _13171_, _01206_);
  nand (_13173_, _01290_, _26867_);
  nand (_13174_, _01296_, _26839_);
  nand (_13175_, _13174_, _13173_);
  nand (_13176_, _13175_, _01204_);
  nand (_13177_, _13176_, _13172_);
  nand (_13178_, _13177_, _01262_);
  nor (_13179_, _01296_, _26924_);
  nor (_13180_, _01290_, _26896_);
  nor (_13181_, _13180_, _13179_);
  nand (_13182_, _13181_, _01206_);
  nand (_13183_, _01290_, _26981_);
  nand (_13184_, _01296_, _26952_);
  nand (_13185_, _13184_, _13183_);
  nand (_13186_, _13185_, _01204_);
  nand (_13187_, _13186_, _13182_);
  nand (_13188_, _13187_, _01260_);
  nand (_13189_, _13188_, _13178_);
  nand (_13190_, _13189_, _01274_);
  nand (_13191_, _01296_, _27066_);
  nand (_13192_, _01290_, _27094_);
  nand (_13193_, _13192_, _13191_);
  nand (_13194_, _13193_, _01204_);
  nand (_13195_, _01290_, _27037_);
  nand (_13196_, _01296_, _27009_);
  nand (_13197_, _13196_, _13195_);
  nand (_13198_, _13197_, _01206_);
  nand (_13199_, _13198_, _13194_);
  nand (_13200_, _13199_, _01262_);
  nand (_13201_, _01296_, _27179_);
  nand (_13202_, _01290_, _27207_);
  nand (_13203_, _13202_, _13201_);
  nand (_13204_, _13203_, _01204_);
  nand (_13205_, _01290_, _27151_);
  nand (_13206_, _01296_, _27122_);
  nand (_13208_, _13206_, _13205_);
  nand (_13209_, _13208_, _01206_);
  nand (_13210_, _13209_, _13204_);
  nand (_13211_, _13210_, _01260_);
  nand (_13212_, _13211_, _13200_);
  nand (_13213_, _13212_, _01275_);
  nand (_13214_, _13213_, _13190_);
  nand (_13215_, _13214_, _01308_);
  nand (_13216_, _13215_, _13168_);
  nand (_13217_, _13216_, _01244_);
  nand (_13218_, _13217_, _13120_);
  nor (_13219_, _13218_, _01235_);
  nor (_13220_, _13219_, _13023_);
  nor (_13221_, _13220_, _28717_);
  nand (_13222_, _01290_, _24855_);
  nand (_13223_, _01296_, _24840_);
  nand (_13224_, _13223_, _13222_);
  nand (_13225_, _13224_, _01204_);
  nand (_13226_, _01296_, _24812_);
  nand (_13227_, _01290_, _24826_);
  nand (_13228_, _13227_, _13226_);
  nand (_13229_, _13228_, _01206_);
  nand (_13230_, _13229_, _13225_);
  nand (_13231_, _13230_, _01260_);
  nand (_13232_, _01290_, _24797_);
  nand (_13233_, _01296_, _24783_);
  nand (_13234_, _13233_, _13232_);
  nand (_13235_, _13234_, _01204_);
  nand (_13236_, _01296_, _24754_);
  nand (_13237_, _01290_, _24769_);
  nand (_13238_, _13237_, _13236_);
  nand (_13239_, _13238_, _01206_);
  nand (_13240_, _13239_, _13235_);
  nand (_13241_, _13240_, _01262_);
  nand (_13242_, _13241_, _13231_);
  nand (_13243_, _13242_, _01275_);
  nor (_13244_, _01296_, _24740_);
  nor (_13245_, _01290_, _24725_);
  nor (_13246_, _13245_, _13244_);
  nand (_13247_, _13246_, _01204_);
  nor (_13249_, _01290_, _24697_);
  nor (_13250_, _01296_, _24711_);
  nor (_13251_, _13250_, _13249_);
  nand (_13252_, _13251_, _01206_);
  nand (_13253_, _13252_, _13247_);
  nand (_13254_, _13253_, _01260_);
  nor (_13255_, _01296_, _24682_);
  nor (_13256_, _01290_, _24668_);
  nor (_13257_, _13256_, _13255_);
  nand (_13258_, _13257_, _01204_);
  nor (_13259_, _01290_, _24639_);
  nor (_13260_, _01296_, _24654_);
  nor (_13261_, _13260_, _13259_);
  nand (_13262_, _13261_, _01206_);
  nand (_13263_, _13262_, _13258_);
  nand (_13264_, _13263_, _01262_);
  nand (_13265_, _13264_, _13254_);
  nand (_13266_, _13265_, _01274_);
  nand (_13267_, _13266_, _13243_);
  nand (_13268_, _13267_, _01241_);
  nand (_13269_, _01296_, _25071_);
  nand (_13270_, _01290_, _25085_);
  nand (_13271_, _13270_, _13269_);
  nand (_13272_, _13271_, _01204_);
  nand (_13273_, _01290_, _25057_);
  nand (_13274_, _01296_, _25042_);
  nand (_13275_, _13274_, _13273_);
  nand (_13276_, _13275_, _01206_);
  nand (_13277_, _13276_, _13272_);
  nand (_13278_, _13277_, _01260_);
  nand (_13279_, _01296_, _25013_);
  nand (_13280_, _01290_, _25028_);
  nand (_13281_, _13280_, _13279_);
  nand (_13282_, _13281_, _01204_);
  nand (_13283_, _01290_, _24999_);
  nand (_13284_, _01296_, _24985_);
  nand (_13285_, _13284_, _13283_);
  nand (_13286_, _13285_, _01206_);
  nand (_13287_, _13286_, _13282_);
  nand (_13288_, _13287_, _01262_);
  nand (_13290_, _13288_, _13278_);
  nand (_13291_, _13290_, _01275_);
  nor (_13292_, _01296_, _24942_);
  nor (_13293_, _01290_, _24926_);
  nor (_13294_, _13293_, _13292_);
  nand (_13295_, _13294_, _01206_);
  nand (_13296_, _01290_, _24970_);
  nand (_13297_, _01296_, _24956_);
  nand (_13298_, _13297_, _13296_);
  nand (_13299_, _13298_, _01204_);
  nand (_13300_, _13299_, _13295_);
  nand (_13301_, _13300_, _01260_);
  nor (_13302_, _01296_, _24883_);
  nor (_13303_, _01290_, _24869_);
  nor (_13304_, _13303_, _13302_);
  nand (_13305_, _13304_, _01206_);
  nand (_13306_, _01290_, _24912_);
  nand (_13307_, _01296_, _24898_);
  nand (_13308_, _13307_, _13306_);
  nand (_13309_, _13308_, _01204_);
  nand (_13310_, _13309_, _13305_);
  nand (_13311_, _13310_, _01262_);
  nand (_13312_, _13311_, _13301_);
  nand (_13313_, _13312_, _01274_);
  nand (_13314_, _13313_, _13291_);
  nand (_13315_, _13314_, _01308_);
  nand (_13316_, _13315_, _13268_);
  nand (_13317_, _13316_, _01245_);
  nand (_13318_, _01296_, _25474_);
  nand (_13319_, _01290_, _25488_);
  nand (_13320_, _13319_, _13318_);
  nand (_13321_, _13320_, _01204_);
  nand (_13322_, _01290_, _25459_);
  nand (_13323_, _01296_, _25445_);
  nand (_13324_, _13323_, _13322_);
  nand (_13325_, _13324_, _01206_);
  nand (_13326_, _13325_, _13321_);
  nand (_13327_, _13326_, _01260_);
  nand (_13328_, _01296_, _25416_);
  nand (_13329_, _01290_, _25431_);
  nand (_13331_, _13329_, _13328_);
  nand (_13332_, _13331_, _01204_);
  nand (_13333_, _01290_, _25402_);
  nand (_13334_, _01296_, _25388_);
  nand (_13335_, _13334_, _13333_);
  nand (_13336_, _13335_, _01206_);
  nand (_13337_, _13336_, _13332_);
  nand (_13338_, _13337_, _01262_);
  nand (_13339_, _13338_, _13327_);
  nand (_13340_, _13339_, _01275_);
  nor (_13341_, _01296_, _25345_);
  nor (_13342_, _01290_, _25329_);
  nor (_13343_, _13342_, _13341_);
  nand (_13344_, _13343_, _01206_);
  nand (_13345_, _01290_, _25373_);
  nand (_13346_, _01296_, _25359_);
  nand (_13347_, _13346_, _13345_);
  nand (_13348_, _13347_, _01204_);
  nand (_13349_, _13348_, _13344_);
  nand (_13350_, _13349_, _01260_);
  nor (_13351_, _01296_, _25286_);
  nor (_13352_, _01290_, _25272_);
  nor (_13353_, _13352_, _13351_);
  nand (_13354_, _13353_, _01206_);
  nand (_13355_, _01290_, _25315_);
  nand (_13356_, _01296_, _25300_);
  nand (_13357_, _13356_, _13355_);
  nand (_13358_, _13357_, _01204_);
  nand (_13359_, _13358_, _13354_);
  nand (_13360_, _13359_, _01262_);
  nand (_13361_, _13360_, _13350_);
  nand (_13362_, _13361_, _01274_);
  nand (_13363_, _13362_, _13340_);
  nand (_13364_, _13363_, _01308_);
  nand (_13365_, _01290_, _25257_);
  nand (_13366_, _01296_, _25243_);
  nand (_13367_, _13366_, _13365_);
  nand (_13368_, _13367_, _01204_);
  nand (_13369_, _01296_, _25214_);
  nand (_13370_, _01290_, _25229_);
  nand (_13372_, _13370_, _13369_);
  nand (_13373_, _13372_, _01206_);
  nand (_13374_, _13373_, _13368_);
  nand (_13375_, _13374_, _01260_);
  nand (_13376_, _01290_, _25200_);
  nand (_13377_, _01296_, _25186_);
  nand (_13378_, _13377_, _13376_);
  nand (_13379_, _13378_, _01204_);
  nand (_13380_, _01296_, _25157_);
  nand (_13381_, _01290_, _25171_);
  nand (_13382_, _13381_, _13380_);
  nand (_13383_, _13382_, _01206_);
  nand (_13384_, _13383_, _13379_);
  nand (_13385_, _13384_, _01262_);
  nand (_13386_, _13385_, _13375_);
  nand (_13387_, _13386_, _01275_);
  nor (_13388_, _01296_, _25143_);
  nor (_13389_, _01290_, _25128_);
  nor (_13390_, _13389_, _13388_);
  nand (_13391_, _13390_, _01204_);
  nor (_13392_, _01290_, _23680_);
  nor (_13393_, _01296_, _25114_);
  nor (_13394_, _13393_, _13392_);
  nand (_13395_, _13394_, _01206_);
  nand (_13396_, _13395_, _13391_);
  nand (_13397_, _13396_, _01260_);
  nor (_13398_, _01296_, _23651_);
  nor (_13399_, _01290_, _23637_);
  nor (_13400_, _13399_, _13398_);
  nand (_13401_, _13400_, _01204_);
  nor (_13402_, _01290_, _25100_);
  nor (_13403_, _01296_, _23666_);
  nor (_13404_, _13403_, _13402_);
  nand (_13405_, _13404_, _01206_);
  nand (_13406_, _13405_, _13401_);
  nand (_13407_, _13406_, _01262_);
  nand (_13408_, _13407_, _13397_);
  nand (_13409_, _13408_, _01274_);
  nand (_13410_, _13409_, _13387_);
  nand (_13411_, _13410_, _01241_);
  nand (_13413_, _13411_, _13364_);
  nand (_13414_, _13413_, _01244_);
  nand (_13415_, _13414_, _13317_);
  nor (_13416_, _13415_, _01231_);
  nand (_13417_, _01296_, _24150_);
  nand (_13418_, _01290_, _24165_);
  nand (_13419_, _13418_, _13417_);
  nand (_13420_, _13419_, _01204_);
  nand (_13421_, _01290_, _24136_);
  nand (_13422_, _01296_, _24122_);
  nand (_13423_, _13422_, _13421_);
  nand (_13424_, _13423_, _01206_);
  nand (_13425_, _13424_, _13420_);
  nand (_13426_, _13425_, _01260_);
  nand (_13427_, _01296_, _24092_);
  nand (_13428_, _01290_, _24106_);
  nand (_13429_, _13428_, _13427_);
  nand (_13430_, _13429_, _01204_);
  nand (_13431_, _01290_, _24078_);
  nand (_13432_, _01296_, _24063_);
  nand (_13433_, _13432_, _13431_);
  nand (_13434_, _13433_, _01206_);
  nand (_13435_, _13434_, _13430_);
  nand (_13436_, _13435_, _01262_);
  nand (_13437_, _13436_, _13426_);
  nand (_13438_, _13437_, _01275_);
  nor (_13439_, _01296_, _24020_);
  nor (_13440_, _01290_, _24006_);
  nor (_13441_, _13440_, _13439_);
  nand (_13442_, _13441_, _01206_);
  nand (_13443_, _01290_, _24049_);
  nand (_13444_, _01296_, _24035_);
  nand (_13445_, _13444_, _13443_);
  nand (_13446_, _13445_, _01204_);
  nand (_13447_, _13446_, _13442_);
  nand (_13448_, _13447_, _01260_);
  nor (_13449_, _01296_, _23963_);
  nor (_13450_, _01290_, _23949_);
  nor (_13451_, _13450_, _13449_);
  nand (_13452_, _13451_, _01206_);
  nand (_13454_, _01290_, _23992_);
  nand (_13455_, _01296_, _23977_);
  nand (_13456_, _13455_, _13454_);
  nand (_13457_, _13456_, _01204_);
  nand (_13458_, _13457_, _13452_);
  nand (_13459_, _13458_, _01262_);
  nand (_13460_, _13459_, _13448_);
  nand (_13461_, _13460_, _01274_);
  nand (_13462_, _13461_, _13438_);
  nand (_13463_, _13462_, _01308_);
  nand (_13464_, _01290_, _23934_);
  nand (_13465_, _01296_, _23920_);
  nand (_13466_, _13465_, _13464_);
  nand (_13467_, _13466_, _01204_);
  nand (_13468_, _01296_, _23891_);
  nand (_13469_, _01290_, _23906_);
  nand (_13470_, _13469_, _13468_);
  nand (_13471_, _13470_, _01206_);
  nand (_13472_, _13471_, _13467_);
  nand (_13473_, _13472_, _01260_);
  nand (_13474_, _01290_, _23877_);
  nand (_13475_, _01296_, _23862_);
  nand (_13476_, _13475_, _13474_);
  nand (_13477_, _13476_, _01204_);
  nand (_13478_, _01296_, _23834_);
  nand (_13479_, _01290_, _23848_);
  nand (_13480_, _13479_, _13478_);
  nand (_13481_, _13480_, _01206_);
  nand (_13482_, _13481_, _13477_);
  nand (_13483_, _13482_, _01262_);
  nand (_13484_, _13483_, _13473_);
  nand (_13485_, _13484_, _01275_);
  nor (_13486_, _01296_, _23819_);
  nor (_13487_, _01290_, _23805_);
  nor (_13488_, _13487_, _13486_);
  nand (_13489_, _13488_, _01204_);
  nor (_13490_, _01290_, _23776_);
  nor (_13491_, _01296_, _23791_);
  nor (_13492_, _13491_, _13490_);
  nand (_13493_, _13492_, _01206_);
  nand (_13495_, _13493_, _13489_);
  nand (_13496_, _13495_, _01260_);
  nor (_13497_, _01296_, _23762_);
  nor (_13498_, _01290_, _23748_);
  nor (_13499_, _13498_, _13497_);
  nand (_13500_, _13499_, _01204_);
  nor (_13501_, _01290_, _23719_);
  nor (_13502_, _01296_, _23733_);
  nor (_13503_, _13502_, _13501_);
  nand (_13504_, _13503_, _01206_);
  nand (_13506_, _13504_, _13500_);
  nand (_13507_, _13506_, _01262_);
  nand (_13508_, _13507_, _13496_);
  nand (_13509_, _13508_, _01274_);
  nand (_13510_, _13509_, _13485_);
  nand (_13511_, _13510_, _01241_);
  nand (_13512_, _13511_, _13463_);
  nand (_13513_, _13512_, _01245_);
  nor (_13514_, _01296_, _24222_);
  nor (_13515_, _01290_, _24208_);
  nor (_13516_, _13515_, _13514_);
  nand (_13517_, _13516_, _01204_);
  nor (_13518_, _01290_, _24179_);
  nor (_13519_, _01296_, _24194_);
  nor (_13520_, _13519_, _13518_);
  nand (_13521_, _13520_, _01206_);
  nand (_13522_, _13521_, _13517_);
  nand (_13523_, _13522_, _01262_);
  nor (_13524_, _01296_, _24280_);
  nor (_13525_, _01290_, _24265_);
  nor (_13526_, _13525_, _13524_);
  nand (_13527_, _13526_, _01204_);
  nor (_13528_, _01290_, _24237_);
  nor (_13529_, _01296_, _24251_);
  nor (_13530_, _13529_, _13528_);
  nand (_13531_, _13530_, _01206_);
  nand (_13532_, _13531_, _13527_);
  nand (_13533_, _13532_, _01260_);
  nand (_13534_, _13533_, _13523_);
  nand (_13535_, _13534_, _01274_);
  nand (_13537_, _01290_, _24337_);
  nand (_13538_, _01296_, _24323_);
  nand (_13539_, _13538_, _13537_);
  nand (_13540_, _13539_, _01204_);
  nand (_13541_, _01296_, _24294_);
  nand (_13542_, _01290_, _24308_);
  nand (_13543_, _13542_, _13541_);
  nand (_13544_, _13543_, _01206_);
  nand (_13545_, _13544_, _13540_);
  nand (_13546_, _13545_, _01262_);
  nand (_13547_, _01290_, _24394_);
  nand (_13548_, _01296_, _24380_);
  nand (_13549_, _13548_, _13547_);
  nand (_13550_, _13549_, _01204_);
  nand (_13551_, _01296_, _24351_);
  nand (_13552_, _01290_, _24366_);
  nand (_13553_, _13552_, _13551_);
  nand (_13554_, _13553_, _01206_);
  nand (_13555_, _13554_, _13550_);
  nand (_13556_, _13555_, _01260_);
  nand (_13557_, _13556_, _13546_);
  nand (_13558_, _13557_, _01275_);
  nand (_13559_, _13558_, _13535_);
  nand (_13560_, _13559_, _01241_);
  nor (_13561_, _01296_, _24423_);
  nor (_13562_, _01290_, _24409_);
  nor (_13563_, _13562_, _13561_);
  nand (_13564_, _13563_, _01206_);
  nand (_13565_, _01290_, _24452_);
  nand (_13566_, _01296_, _24437_);
  nand (_13567_, _13566_, _13565_);
  nand (_13568_, _13567_, _01204_);
  nand (_13569_, _13568_, _13564_);
  nand (_13570_, _13569_, _01262_);
  nor (_13571_, _01296_, _24481_);
  nor (_13572_, _01290_, _24466_);
  nor (_13573_, _13572_, _13571_);
  nand (_13574_, _13573_, _01206_);
  nand (_13575_, _01290_, _24509_);
  nand (_13576_, _01296_, _24495_);
  nand (_13578_, _13576_, _13575_);
  nand (_13579_, _13578_, _01204_);
  nand (_13580_, _13579_, _13574_);
  nand (_13581_, _13580_, _01260_);
  nand (_13582_, _13581_, _13570_);
  nand (_13583_, _13582_, _01274_);
  nand (_13584_, _01296_, _24553_);
  nand (_13585_, _01290_, _24568_);
  nand (_13586_, _13585_, _13584_);
  nand (_13587_, _13586_, _01204_);
  nand (_13588_, _01290_, _24539_);
  nand (_13589_, _01296_, _24525_);
  nand (_13590_, _13589_, _13588_);
  nand (_13591_, _13590_, _01206_);
  nand (_13592_, _13591_, _13587_);
  nand (_13593_, _13592_, _01262_);
  nand (_13594_, _01296_, _24611_);
  nand (_13595_, _01290_, _24625_);
  nand (_13596_, _13595_, _13594_);
  nand (_13597_, _13596_, _01204_);
  nand (_13598_, _01290_, _24596_);
  nand (_13599_, _01296_, _24582_);
  nand (_13600_, _13599_, _13598_);
  nand (_13601_, _13600_, _01206_);
  nand (_13602_, _13601_, _13597_);
  nand (_13603_, _13602_, _01260_);
  nand (_13604_, _13603_, _13593_);
  nand (_13605_, _13604_, _01275_);
  nand (_13606_, _13605_, _13583_);
  nand (_13607_, _13606_, _01308_);
  nand (_13608_, _13607_, _13560_);
  nand (_13609_, _13608_, _01244_);
  nand (_13610_, _13609_, _13513_);
  nor (_13611_, _13610_, _01235_);
  nor (_13612_, _13611_, _13416_);
  nor (_13613_, _13612_, _28718_);
  nor (_13614_, _13613_, _13221_);
  nor (_13615_, _13614_, _06280_);
  nand (_13616_, _06280_, _27140_);
  nand (_13617_, _13616_, _29344_);
  nor (_15271_, _13617_, _13615_);
  not (_13619_, _00891_);
  nor (_13620_, _13619_, _15473_);
  nor (_15488_, _13620_, _01011_);
  nor (_13621_, _01159_, _01304_);
  nor (_13622_, _01240_, _01304_);
  nor (_13623_, _01243_, _01304_);
  nor (_13624_, _13623_, _13622_);
  not (_13625_, _13624_);
  nor (_13626_, _01160_, _27612_);
  not (_13627_, _13626_);
  nor (_13628_, _13627_, _01304_);
  nor (_13629_, _13628_, _13625_);
  not (_13630_, _13629_);
  nor (_13631_, _01255_, _01304_);
  nor (_13632_, _01270_, _01304_);
  nor (_13633_, _13632_, _13631_);
  not (_13634_, _13633_);
  nor (_13635_, _01285_, _01304_);
  not (_13636_, _13635_);
  nor (_13637_, _01164_, _01304_);
  nor (_13638_, _13637_, _13636_);
  not (_13639_, _13638_);
  nor (_13640_, _13639_, _13634_);
  not (_13641_, _13640_);
  nor (_13642_, _13641_, _13630_);
  nand (_13643_, _13642_, _13621_);
  not (_13644_, _13642_);
  nand (_13645_, _13644_, _15535_);
  nand (_15543_, _13645_, _13643_);
  not (_13646_, _13637_);
  nor (_13647_, _13646_, _13635_);
  not (_13648_, _13647_);
  nor (_13649_, _13648_, _13634_);
  not (_13650_, _13649_);
  nor (_13651_, _13650_, _13630_);
  nand (_13652_, _13651_, _13621_);
  not (_13653_, _13651_);
  nand (_13654_, _13653_, _15591_);
  nand (_15598_, _13654_, _13652_);
  nor (_13656_, _13646_, _13636_);
  not (_13657_, _13656_);
  nor (_13658_, _13657_, _13634_);
  not (_13659_, _13658_);
  nor (_13660_, _13659_, _13630_);
  nand (_13661_, _13660_, _13621_);
  not (_13662_, _13660_);
  nand (_13663_, _13662_, _15633_);
  nand (_15640_, _13663_, _13661_);
  nor (_13664_, _13637_, _13635_);
  not (_13665_, _13664_);
  not (_13666_, _13631_);
  nor (_13667_, _13632_, _13666_);
  not (_13668_, _13667_);
  nor (_13669_, _13668_, _13665_);
  not (_13670_, _13669_);
  nor (_13671_, _13670_, _13630_);
  nand (_13672_, _13671_, _13621_);
  not (_13673_, _13671_);
  nand (_13674_, _13673_, _15689_);
  nand (_15697_, _13674_, _13672_);
  nor (_13675_, _13668_, _13639_);
  not (_13676_, _13675_);
  nor (_13677_, _13676_, _13630_);
  nand (_13678_, _13677_, _13621_);
  not (_13679_, _13677_);
  nand (_13680_, _13679_, _15724_);
  nand (_15732_, _13680_, _13678_);
  nor (_13681_, _13668_, _13648_);
  not (_13682_, _13681_);
  nor (_13683_, _13682_, _13630_);
  nand (_13684_, _13683_, _13621_);
  not (_13685_, _13683_);
  nand (_13686_, _13685_, _15760_);
  nand (_15767_, _13686_, _13684_);
  nor (_13687_, _13668_, _13657_);
  not (_13688_, _13687_);
  nor (_13689_, _13688_, _13630_);
  nand (_13690_, _13689_, _13621_);
  not (_13691_, _13689_);
  nand (_13693_, _13691_, _15795_);
  nand (_15803_, _13693_, _13690_);
  not (_13694_, _13632_);
  nor (_13695_, _13694_, _13631_);
  not (_13696_, _13695_);
  nor (_13697_, _13696_, _13665_);
  not (_13698_, _13697_);
  nor (_13699_, _13698_, _13630_);
  nand (_13700_, _13699_, _13621_);
  not (_13701_, _13699_);
  nand (_13702_, _13701_, _15850_);
  nand (_15858_, _13702_, _13700_);
  nor (_13703_, _13696_, _13639_);
  not (_13704_, _13703_);
  nor (_13705_, _13704_, _13630_);
  nand (_13706_, _13705_, _13621_);
  not (_13707_, _13705_);
  nand (_13708_, _13707_, _15886_);
  nand (_15893_, _13708_, _13706_);
  nor (_13709_, _13696_, _13648_);
  not (_13710_, _13709_);
  nor (_13711_, _13710_, _13630_);
  nand (_13712_, _13711_, _13621_);
  not (_13713_, _13711_);
  nand (_13714_, _13713_, _15921_);
  nand (_15929_, _13714_, _13712_);
  nor (_13715_, _13696_, _13657_);
  not (_13716_, _13715_);
  nor (_13717_, _13716_, _13630_);
  nand (_13718_, _13717_, _13621_);
  not (_13719_, _13717_);
  nand (_13720_, _13719_, _15956_);
  nand (_15964_, _13720_, _13718_);
  nor (_13721_, _13694_, _13666_);
  not (_13722_, _13721_);
  nor (_13723_, _13722_, _13665_);
  not (_13724_, _13723_);
  nor (_13725_, _13724_, _13630_);
  nand (_13726_, _13725_, _13621_);
  not (_13727_, _13725_);
  nand (_13729_, _13727_, _15999_);
  nand (_16007_, _13729_, _13726_);
  nor (_13730_, _13722_, _13639_);
  not (_13731_, _13730_);
  nor (_13732_, _13731_, _13630_);
  nand (_13733_, _13732_, _13621_);
  not (_13734_, _13732_);
  nand (_13735_, _13734_, _16035_);
  nand (_16042_, _13735_, _13733_);
  nor (_13736_, _13722_, _13648_);
  not (_13737_, _13736_);
  nor (_13738_, _13737_, _13630_);
  nand (_13739_, _13738_, _13621_);
  not (_13740_, _13738_);
  nand (_13741_, _13740_, _16070_);
  nand (_16078_, _13741_, _13739_);
  nor (_13742_, _13722_, _13657_);
  not (_13743_, _13742_);
  nor (_13744_, _13743_, _13630_);
  nand (_13745_, _13744_, _13621_);
  not (_13746_, _13744_);
  nand (_13747_, _13746_, _16105_);
  nand (_16113_, _13747_, _13745_);
  nor (_13748_, _13634_, _13665_);
  not (_13749_, _13748_);
  not (_13750_, _13622_);
  nor (_13751_, _13623_, _13750_);
  not (_13752_, _13751_);
  nor (_13753_, _13752_, _13626_);
  not (_13754_, _13753_);
  nor (_13755_, _13754_, _13749_);
  nand (_13756_, _13755_, _13621_);
  not (_13757_, _13755_);
  nand (_13758_, _13757_, _16161_);
  nand (_16168_, _13758_, _13756_);
  nor (_13759_, _13754_, _13641_);
  nand (_13760_, _13759_, _13621_);
  not (_13761_, _13759_);
  nand (_13762_, _13761_, _16189_);
  nand (_16197_, _13762_, _13760_);
  nor (_13764_, _13754_, _13650_);
  nand (_13765_, _13764_, _13621_);
  not (_13766_, _13764_);
  nand (_13767_, _13766_, _16218_);
  nand (_16226_, _13767_, _13765_);
  nor (_13768_, _13754_, _13659_);
  nand (_13769_, _13768_, _13621_);
  not (_13770_, _13768_);
  nand (_13771_, _13770_, _16247_);
  nand (_16255_, _13771_, _13769_);
  nor (_13772_, _13754_, _13670_);
  nand (_13773_, _13772_, _13621_);
  not (_13774_, _13772_);
  nand (_13775_, _13774_, _16276_);
  nand (_16284_, _13775_, _13773_);
  nor (_13776_, _13754_, _13676_);
  nand (_13777_, _13776_, _13621_);
  not (_13778_, _13776_);
  nand (_13779_, _13778_, _16305_);
  nand (_16313_, _13779_, _13777_);
  nor (_13780_, _13754_, _13682_);
  nand (_13781_, _13780_, _13621_);
  not (_13782_, _13780_);
  nand (_13783_, _13782_, _16334_);
  nand (_16341_, _13783_, _13781_);
  nor (_13784_, _13754_, _13688_);
  nand (_13785_, _13784_, _13621_);
  not (_13786_, _13784_);
  nand (_13787_, _13786_, _16362_);
  nand (_16370_, _13787_, _13785_);
  nor (_13788_, _13754_, _13698_);
  nand (_13789_, _13788_, _13621_);
  not (_13790_, _13788_);
  nand (_13791_, _13790_, _16391_);
  nand (_16399_, _13791_, _13789_);
  nor (_13792_, _13754_, _13704_);
  nand (_13793_, _13792_, _13621_);
  not (_13794_, _13792_);
  nand (_13795_, _13794_, _16420_);
  nand (_16427_, _13795_, _13793_);
  nor (_13797_, _13754_, _13710_);
  nand (_13798_, _13797_, _13621_);
  not (_13799_, _13797_);
  nand (_13800_, _13799_, _16448_);
  nand (_16456_, _13800_, _13798_);
  nor (_13801_, _13754_, _13716_);
  nand (_13802_, _13801_, _13621_);
  not (_13803_, _13801_);
  nand (_13804_, _13803_, _16477_);
  nand (_16485_, _13804_, _13802_);
  nor (_13805_, _13754_, _13724_);
  nand (_13806_, _13805_, _13621_);
  not (_13807_, _13805_);
  nand (_13808_, _13807_, _16506_);
  nand (_16513_, _13808_, _13806_);
  nor (_13809_, _13754_, _13731_);
  nand (_13810_, _13809_, _13621_);
  not (_13811_, _13809_);
  nand (_13812_, _13811_, _16534_);
  nand (_16543_, _13812_, _13810_);
  nor (_13813_, _13754_, _13737_);
  nand (_13814_, _13813_, _13621_);
  not (_13815_, _13813_);
  nand (_13816_, _13815_, _16564_);
  nand (_16572_, _13816_, _13814_);
  nor (_13817_, _13754_, _13743_);
  nand (_13818_, _13817_, _13621_);
  not (_13819_, _13817_);
  nand (_13820_, _13819_, _16593_);
  nand (_16600_, _13820_, _13818_);
  not (_13821_, _13623_);
  nor (_13822_, _13821_, _13622_);
  not (_13823_, _13822_);
  nor (_13824_, _13823_, _13626_);
  not (_13825_, _13824_);
  nor (_13826_, _13825_, _13749_);
  nand (_13827_, _13826_, _13621_);
  not (_13828_, _13826_);
  nand (_13829_, _13828_, _16648_);
  nand (_16656_, _13829_, _13827_);
  nor (_13831_, _13825_, _13641_);
  nand (_13832_, _13831_, _13621_);
  not (_13833_, _13831_);
  nand (_13834_, _13833_, _16677_);
  nand (_16684_, _13834_, _13832_);
  nor (_13835_, _13825_, _13650_);
  nand (_13836_, _13835_, _13621_);
  not (_13837_, _13835_);
  nand (_13838_, _13837_, _16705_);
  nand (_16713_, _13838_, _13836_);
  nor (_13839_, _13825_, _13659_);
  nand (_13840_, _13839_, _13621_);
  not (_13841_, _13839_);
  nand (_13842_, _13841_, _16734_);
  nand (_16742_, _13842_, _13840_);
  nor (_13843_, _13825_, _13670_);
  nand (_13844_, _13843_, _13621_);
  not (_13845_, _13843_);
  nand (_13846_, _13845_, _16763_);
  nand (_16770_, _13846_, _13844_);
  nor (_13847_, _13825_, _13676_);
  nand (_13848_, _13847_, _13621_);
  not (_13849_, _13847_);
  nand (_13850_, _13849_, _16791_);
  nand (_16799_, _13850_, _13848_);
  nor (_13851_, _13825_, _13682_);
  nand (_13852_, _13851_, _13621_);
  not (_13853_, _13851_);
  nand (_13854_, _13853_, _16820_);
  nand (_16829_, _13854_, _13852_);
  nor (_13855_, _13825_, _13688_);
  nand (_13856_, _13855_, _13621_);
  not (_13857_, _13855_);
  nand (_13858_, _13857_, _16850_);
  nand (_16857_, _13858_, _13856_);
  nor (_13859_, _13825_, _13698_);
  nand (_13860_, _13859_, _13621_);
  not (_13861_, _13859_);
  nand (_13862_, _13861_, _16878_);
  nand (_16886_, _13862_, _13860_);
  nor (_13864_, _13825_, _13704_);
  nand (_13865_, _13864_, _13621_);
  not (_13866_, _13864_);
  nand (_13867_, _13866_, _16907_);
  nand (_16915_, _13867_, _13865_);
  nor (_13868_, _13825_, _13710_);
  nand (_13869_, _13868_, _13621_);
  not (_13870_, _13868_);
  nand (_13871_, _13870_, _16936_);
  nand (_16943_, _13871_, _13869_);
  nor (_13873_, _13825_, _13716_);
  nand (_13874_, _13873_, _13621_);
  not (_13875_, _13873_);
  nand (_13876_, _13875_, _16964_);
  nand (_16972_, _13876_, _13874_);
  nor (_13877_, _13825_, _13724_);
  nand (_13878_, _13877_, _13621_);
  not (_13879_, _13877_);
  nand (_13880_, _13879_, _16993_);
  nand (_17001_, _13880_, _13878_);
  nor (_13881_, _13825_, _13731_);
  nand (_13882_, _13881_, _13621_);
  not (_13883_, _13881_);
  nand (_13884_, _13883_, _17022_);
  nand (_17029_, _13884_, _13882_);
  nor (_13885_, _13825_, _13737_);
  nand (_13886_, _13885_, _13621_);
  not (_13887_, _13885_);
  nand (_13888_, _13887_, _17050_);
  nand (_17058_, _13888_, _13886_);
  nor (_13889_, _13825_, _13743_);
  nand (_13890_, _13889_, _13621_);
  not (_13891_, _13889_);
  nand (_13892_, _13891_, _17079_);
  nand (_17087_, _13892_, _13890_);
  nor (_13893_, _13821_, _01240_);
  not (_13894_, _13893_);
  nor (_13895_, _13894_, _13626_);
  not (_13896_, _13895_);
  nor (_13897_, _13896_, _13749_);
  nand (_13899_, _13897_, _13621_);
  not (_13900_, _13897_);
  nand (_13901_, _13900_, _17122_);
  nand (_17130_, _13901_, _13899_);
  nor (_13902_, _13896_, _13641_);
  nand (_13903_, _13902_, _13621_);
  not (_13904_, _13902_);
  nand (_13905_, _13904_, _17151_);
  nand (_17158_, _13905_, _13903_);
  nor (_13906_, _13896_, _13650_);
  nand (_13907_, _13906_, _13621_);
  not (_13908_, _13906_);
  nand (_13909_, _13908_, _17179_);
  nand (_17187_, _13909_, _13907_);
  nor (_13910_, _13896_, _13659_);
  nand (_13911_, _13910_, _13621_);
  not (_13912_, _13910_);
  nand (_13913_, _13912_, _17208_);
  nand (_17216_, _13913_, _13911_);
  nor (_13914_, _13896_, _13670_);
  nand (_13915_, _13914_, _13621_);
  not (_13916_, _13914_);
  nand (_13917_, _13916_, _17237_);
  nand (_17244_, _13917_, _13915_);
  nor (_13918_, _13896_, _13676_);
  nand (_13919_, _13918_, _13621_);
  not (_13920_, _13918_);
  nand (_13921_, _13920_, _17265_);
  nand (_17273_, _13921_, _13919_);
  nor (_13922_, _13896_, _13682_);
  nand (_13923_, _13922_, _13621_);
  not (_13924_, _13922_);
  nand (_13925_, _13924_, _17294_);
  nand (_17302_, _13925_, _13923_);
  nor (_13926_, _13896_, _13688_);
  nand (_13927_, _13926_, _13621_);
  not (_13928_, _13926_);
  nand (_13929_, _13928_, _17323_);
  nand (_17330_, _13929_, _13927_);
  nor (_13930_, _13896_, _13698_);
  nand (_13932_, _13930_, _13621_);
  not (_13933_, _13930_);
  nand (_13934_, _13933_, _17351_);
  nand (_17359_, _13934_, _13932_);
  nor (_13935_, _13896_, _13704_);
  nand (_13936_, _13935_, _13621_);
  not (_13937_, _13935_);
  nand (_13938_, _13937_, _17380_);
  nand (_17388_, _13938_, _13936_);
  nor (_13939_, _13896_, _13710_);
  nand (_13940_, _13939_, _13621_);
  not (_13941_, _13939_);
  nand (_13942_, _13941_, _17411_);
  nand (_17418_, _13942_, _13940_);
  nor (_13943_, _13896_, _13716_);
  nand (_13944_, _13943_, _13621_);
  not (_13945_, _13943_);
  nand (_13946_, _13945_, _17439_);
  nand (_17447_, _13946_, _13944_);
  nor (_13947_, _13896_, _13724_);
  nand (_13948_, _13947_, _13621_);
  not (_13949_, _13947_);
  nand (_13950_, _13949_, _17468_);
  nand (_17476_, _13950_, _13948_);
  nor (_13951_, _13896_, _13731_);
  nand (_13952_, _13951_, _13621_);
  not (_13953_, _13951_);
  nand (_13954_, _13953_, _17497_);
  nand (_17504_, _13954_, _13952_);
  nor (_13955_, _13896_, _13737_);
  nand (_13956_, _13955_, _13621_);
  not (_13957_, _13955_);
  nand (_13958_, _13957_, _17525_);
  nand (_17533_, _13958_, _13956_);
  nor (_13959_, _13896_, _13743_);
  nand (_13960_, _13959_, _13621_);
  not (_13961_, _13959_);
  nand (_13962_, _13961_, _17554_);
  nand (_17562_, _13962_, _13960_);
  nor (_13963_, _26781_, _27608_);
  nand (_13965_, _13963_, _01210_);
  nor (_13966_, _13965_, _13625_);
  not (_13967_, _13966_);
  nor (_13968_, _13967_, _13749_);
  nand (_13969_, _13968_, _13621_);
  not (_13970_, _13968_);
  nand (_13971_, _13970_, _17609_);
  nand (_17617_, _13971_, _13969_);
  nor (_13972_, _13967_, _13641_);
  nand (_13973_, _13972_, _13621_);
  not (_13974_, _13972_);
  nand (_13975_, _13974_, _17638_);
  nand (_17646_, _13975_, _13973_);
  nor (_13976_, _13967_, _13650_);
  nand (_13977_, _13976_, _13621_);
  not (_13978_, _13976_);
  nand (_13979_, _13978_, _17667_);
  nand (_17674_, _13979_, _13977_);
  nor (_13980_, _13967_, _13659_);
  nand (_13981_, _13980_, _13621_);
  not (_13982_, _13980_);
  nand (_13983_, _13982_, _17696_);
  nand (_17704_, _13983_, _13981_);
  nor (_13984_, _13967_, _13670_);
  nand (_13985_, _13984_, _13621_);
  not (_13986_, _13984_);
  nand (_13987_, _13986_, _17725_);
  nand (_17733_, _13987_, _13985_);
  nor (_13988_, _13967_, _13676_);
  nand (_13989_, _13988_, _13621_);
  not (_13990_, _13988_);
  nand (_13991_, _13990_, _17754_);
  nand (_17761_, _13991_, _13989_);
  nor (_13992_, _13967_, _13682_);
  nand (_13993_, _13992_, _13621_);
  not (_13994_, _13992_);
  nand (_13995_, _13994_, _17782_);
  nand (_17790_, _13995_, _13993_);
  nor (_13996_, _13967_, _13688_);
  nand (_13997_, _13996_, _13621_);
  not (_13999_, _13996_);
  nand (_14000_, _13999_, _17811_);
  nand (_17819_, _14000_, _13997_);
  nor (_14001_, _13967_, _13698_);
  nand (_14002_, _14001_, _13621_);
  not (_14003_, _14001_);
  nand (_14004_, _14003_, _17840_);
  nand (_17847_, _14004_, _14002_);
  nor (_14005_, _13967_, _13704_);
  nand (_14006_, _14005_, _13621_);
  not (_14007_, _14005_);
  nand (_14008_, _14007_, _17868_);
  nand (_17876_, _14008_, _14006_);
  nor (_14009_, _13967_, _13710_);
  nand (_14010_, _14009_, _13621_);
  not (_14011_, _14009_);
  nand (_14012_, _14011_, _17897_);
  nand (_17905_, _14012_, _14010_);
  nor (_14013_, _13967_, _13716_);
  nand (_14014_, _14013_, _13621_);
  not (_14015_, _14013_);
  nand (_14016_, _14015_, _17926_);
  nand (_17933_, _14016_, _14014_);
  nor (_14017_, _13967_, _13724_);
  nand (_14018_, _14017_, _13621_);
  not (_14019_, _14017_);
  nand (_14020_, _14019_, _17954_);
  nand (_17962_, _14020_, _14018_);
  nor (_14021_, _13967_, _13731_);
  nand (_14022_, _14021_, _13621_);
  not (_14023_, _14021_);
  nand (_14024_, _14023_, _17984_);
  nand (_17992_, _14024_, _14022_);
  nor (_14025_, _13967_, _13737_);
  nand (_14026_, _14025_, _13621_);
  not (_14027_, _14025_);
  nand (_14028_, _14027_, _18013_);
  nand (_18020_, _14028_, _14026_);
  nor (_14029_, _13967_, _13743_);
  nand (_14030_, _14029_, _13621_);
  not (_14032_, _14029_);
  nand (_14033_, _14032_, _18041_);
  nand (_18049_, _14033_, _14030_);
  nor (_14034_, _13965_, _13752_);
  not (_14035_, _14034_);
  nor (_14036_, _14035_, _13749_);
  nand (_14037_, _14036_, _13621_);
  not (_14038_, _14036_);
  nand (_14039_, _14038_, _18077_);
  nand (_18084_, _14039_, _14037_);
  nor (_14040_, _14035_, _13641_);
  nand (_14041_, _14040_, _13621_);
  not (_14042_, _14040_);
  nand (_14043_, _14042_, _18105_);
  nand (_18113_, _14043_, _14041_);
  nor (_14044_, _14035_, _13650_);
  nand (_14045_, _14044_, _13621_);
  not (_14046_, _14044_);
  nand (_14047_, _14046_, _18134_);
  nand (_18142_, _14047_, _14045_);
  nor (_14048_, _14035_, _13659_);
  nand (_14049_, _14048_, _13621_);
  not (_14050_, _14048_);
  nand (_14051_, _14050_, _18163_);
  nand (_18170_, _14051_, _14049_);
  nor (_14052_, _14035_, _13670_);
  nand (_14053_, _14052_, _13621_);
  not (_14054_, _14052_);
  nand (_14055_, _14054_, _18191_);
  nand (_18199_, _14055_, _14053_);
  nor (_14056_, _14035_, _13676_);
  nand (_14057_, _14056_, _13621_);
  not (_14058_, _14056_);
  nand (_14059_, _14058_, _18220_);
  nand (_18228_, _14059_, _14057_);
  nor (_14060_, _14035_, _13682_);
  nand (_14061_, _14060_, _13621_);
  not (_14062_, _14060_);
  nand (_14063_, _14062_, _18249_);
  nand (_18256_, _14063_, _14061_);
  nor (_14065_, _14035_, _13688_);
  nand (_14066_, _14065_, _13621_);
  not (_14067_, _14065_);
  nand (_14068_, _14067_, _18278_);
  nand (_18286_, _14068_, _14066_);
  nor (_14069_, _14035_, _13698_);
  nand (_14070_, _14069_, _13621_);
  not (_14071_, _14069_);
  nand (_14072_, _14071_, _18307_);
  nand (_18315_, _14072_, _14070_);
  nor (_14073_, _14035_, _13704_);
  nand (_14074_, _14073_, _13621_);
  not (_14075_, _14073_);
  nand (_14076_, _14075_, _18336_);
  nand (_18343_, _14076_, _14074_);
  nor (_14077_, _14035_, _13710_);
  nand (_14078_, _14077_, _13621_);
  not (_14079_, _14077_);
  nand (_14080_, _14079_, _18364_);
  nand (_18372_, _14080_, _14078_);
  nor (_14081_, _14035_, _13716_);
  nand (_14082_, _14081_, _13621_);
  not (_14083_, _14081_);
  nand (_14084_, _14083_, _18393_);
  nand (_18401_, _14084_, _14082_);
  nor (_14085_, _14035_, _13724_);
  nand (_14086_, _14085_, _13621_);
  not (_14087_, _14085_);
  nand (_14088_, _14087_, _18422_);
  nand (_18429_, _14088_, _14086_);
  nor (_14089_, _14035_, _13731_);
  nand (_14090_, _14089_, _13621_);
  not (_14091_, _14089_);
  nand (_14092_, _14091_, _18450_);
  nand (_18458_, _14092_, _14090_);
  nor (_14093_, _14035_, _13737_);
  nand (_14094_, _14093_, _13621_);
  not (_14095_, _14093_);
  nand (_14096_, _14095_, _18479_);
  nand (_18487_, _14096_, _14094_);
  nor (_14098_, _14035_, _13743_);
  nand (_14099_, _14098_, _13621_);
  not (_14100_, _14098_);
  nand (_14101_, _14100_, _18508_);
  nand (_18515_, _14101_, _14099_);
  nor (_14102_, _13965_, _13823_);
  not (_14103_, _14102_);
  nor (_14104_, _14103_, _13749_);
  nand (_14105_, _14104_, _13621_);
  not (_14106_, _14104_);
  nand (_14107_, _14106_, _18543_);
  nand (_18552_, _14107_, _14105_);
  nor (_14108_, _14103_, _13641_);
  nand (_14109_, _14108_, _13621_);
  not (_14110_, _14108_);
  nand (_14111_, _14110_, _18573_);
  nand (_18580_, _14111_, _14109_);
  nor (_14112_, _14103_, _13650_);
  nand (_14113_, _14112_, _13621_);
  not (_14114_, _14112_);
  nand (_14115_, _14114_, _18599_);
  nand (_18608_, _14115_, _14113_);
  nor (_14116_, _14103_, _13659_);
  nand (_14117_, _14116_, _13621_);
  not (_14118_, _14116_);
  nand (_14119_, _14118_, _18633_);
  nand (_18642_, _14119_, _14117_);
  nor (_14120_, _14103_, _13670_);
  nand (_14121_, _14120_, _13621_);
  not (_14122_, _14120_);
  nand (_14123_, _14122_, _18667_);
  nand (_18676_, _14123_, _14121_);
  nor (_14124_, _14103_, _13676_);
  nand (_14125_, _14124_, _13621_);
  not (_14126_, _14124_);
  nand (_14127_, _14126_, _18701_);
  nand (_18710_, _14127_, _14125_);
  nor (_14128_, _14103_, _13682_);
  nand (_14129_, _14128_, _13621_);
  not (_14130_, _14128_);
  nand (_14132_, _14130_, _18735_);
  nand (_18744_, _14132_, _14129_);
  nor (_14133_, _14103_, _13688_);
  nand (_14134_, _14133_, _13621_);
  not (_14135_, _14133_);
  nand (_14136_, _14135_, _18775_);
  nand (_18786_, _14136_, _14134_);
  nor (_14137_, _14103_, _13698_);
  nand (_14138_, _14137_, _13621_);
  not (_14139_, _14137_);
  nand (_14140_, _14139_, _18817_);
  nand (_18828_, _14140_, _14138_);
  nor (_14141_, _14103_, _13704_);
  nand (_14142_, _14141_, _13621_);
  not (_14143_, _14141_);
  nand (_14144_, _14143_, _18859_);
  nand (_18870_, _14144_, _14142_);
  nor (_14145_, _14103_, _13710_);
  nand (_14146_, _14145_, _13621_);
  not (_14147_, _14145_);
  nand (_14148_, _14147_, _18900_);
  nand (_18912_, _14148_, _14146_);
  nor (_14149_, _14103_, _13716_);
  nand (_14150_, _14149_, _13621_);
  not (_14151_, _14149_);
  nand (_14152_, _14151_, _18943_);
  nand (_18954_, _14152_, _14150_);
  nor (_14153_, _14103_, _13724_);
  nand (_14154_, _14153_, _13621_);
  not (_14155_, _14153_);
  nand (_14156_, _14155_, _18985_);
  nand (_18996_, _14156_, _14154_);
  nor (_14157_, _14103_, _13731_);
  nand (_14158_, _14157_, _13621_);
  not (_14159_, _14157_);
  nand (_14160_, _14159_, _19026_);
  nand (_19037_, _14160_, _14158_);
  nor (_14161_, _14103_, _13737_);
  nand (_14162_, _14161_, _13621_);
  not (_14163_, _14161_);
  nand (_14165_, _14163_, _19068_);
  nand (_19079_, _14165_, _14162_);
  nor (_14166_, _14103_, _13743_);
  nand (_14167_, _14166_, _13621_);
  not (_14168_, _14166_);
  nand (_14169_, _14168_, _19109_);
  nand (_19120_, _14169_, _14167_);
  nor (_14170_, _13965_, _13894_);
  not (_14171_, _14170_);
  nor (_14172_, _14171_, _13749_);
  nand (_14173_, _14172_, _13621_);
  not (_14174_, _14172_);
  nand (_14175_, _14174_, _19161_);
  nand (_19171_, _14175_, _14173_);
  nor (_14176_, _14171_, _13641_);
  nand (_14177_, _14176_, _13621_);
  not (_14178_, _14176_);
  nand (_14179_, _14178_, _19202_);
  nand (_19213_, _14179_, _14177_);
  nor (_14180_, _14171_, _13650_);
  nand (_14181_, _14180_, _13621_);
  not (_14182_, _14180_);
  nand (_14183_, _14182_, _19236_);
  nand (_19246_, _14183_, _14181_);
  nor (_14184_, _14171_, _13659_);
  nand (_14185_, _14184_, _13621_);
  not (_14186_, _14184_);
  nand (_14187_, _14186_, _19272_);
  nand (_19281_, _14187_, _14185_);
  nor (_14188_, _14171_, _13670_);
  nand (_14189_, _14188_, _13621_);
  not (_14190_, _14188_);
  nand (_14191_, _14190_, _19311_);
  nand (_19322_, _14191_, _14189_);
  nor (_14192_, _14171_, _13676_);
  nand (_14193_, _14192_, _13621_);
  not (_14194_, _14192_);
  nand (_14195_, _14194_, _19352_);
  nand (_19363_, _14195_, _14193_);
  nor (_14196_, _14171_, _13682_);
  nand (_14198_, _14196_, _13621_);
  not (_14199_, _14196_);
  nand (_14200_, _14199_, _19392_);
  nand (_19403_, _14200_, _14198_);
  nor (_14201_, _14171_, _13688_);
  nand (_14202_, _14201_, _13621_);
  not (_14203_, _14201_);
  nand (_14204_, _14203_, _19432_);
  nand (_19443_, _14204_, _14202_);
  nor (_14205_, _14171_, _13698_);
  nand (_14207_, _14205_, _13621_);
  not (_14208_, _14205_);
  nand (_14209_, _14208_, _19472_);
  nand (_19483_, _14209_, _14207_);
  nor (_14210_, _14171_, _13704_);
  nand (_14211_, _14210_, _13621_);
  not (_14212_, _14210_);
  nand (_14213_, _14212_, _19512_);
  nand (_19523_, _14213_, _14211_);
  nor (_14214_, _14171_, _13710_);
  nand (_14215_, _14214_, _13621_);
  not (_14216_, _14214_);
  nand (_14217_, _14216_, _19552_);
  nand (_19563_, _14217_, _14215_);
  nor (_14218_, _14171_, _13716_);
  nand (_14219_, _14218_, _13621_);
  not (_14220_, _14218_);
  nand (_14221_, _14220_, _19592_);
  nand (_19603_, _14221_, _14219_);
  nor (_14222_, _14171_, _13724_);
  nand (_14223_, _14222_, _13621_);
  not (_14224_, _14222_);
  nand (_14225_, _14224_, _19632_);
  nand (_19643_, _14225_, _14223_);
  nor (_14226_, _14171_, _13731_);
  nand (_14227_, _14226_, _13621_);
  not (_14228_, _14226_);
  nand (_14229_, _14228_, _19672_);
  nand (_19683_, _14229_, _14227_);
  nor (_14230_, _14171_, _13737_);
  nand (_14232_, _14230_, _13621_);
  not (_14233_, _14230_);
  nand (_14234_, _14233_, _19713_);
  nand (_19724_, _14234_, _14232_);
  nor (_14235_, _14171_, _13743_);
  nand (_14236_, _14235_, _13621_);
  not (_14237_, _14235_);
  nand (_14238_, _14237_, _19754_);
  nand (_19764_, _14238_, _14236_);
  nor (_14239_, _01304_, _04274_);
  not (_14240_, _14239_);
  nor (_14241_, _14240_, _13625_);
  not (_14242_, _14241_);
  nor (_14243_, _14242_, _13749_);
  nand (_14244_, _14243_, _13621_);
  not (_14245_, _14243_);
  nand (_14246_, _14245_, _19844_);
  nand (_19854_, _14246_, _14244_);
  nor (_14247_, _14242_, _13641_);
  nand (_14248_, _14247_, _13621_);
  not (_14249_, _14247_);
  nand (_14250_, _14249_, _19885_);
  nand (_19896_, _14250_, _14248_);
  nor (_14251_, _14242_, _13650_);
  nand (_14252_, _14251_, _13621_);
  not (_14253_, _14251_);
  nand (_14254_, _14253_, _19926_);
  nand (_19937_, _14254_, _14252_);
  nor (_14255_, _14242_, _13659_);
  nand (_14256_, _14255_, _13621_);
  not (_14257_, _14255_);
  nand (_14258_, _14257_, _19967_);
  nand (_19978_, _14258_, _14256_);
  nor (_14259_, _14242_, _13670_);
  nand (_14260_, _14259_, _13621_);
  not (_14261_, _14259_);
  nand (_14262_, _14261_, _20008_);
  nand (_20019_, _14262_, _14260_);
  nor (_14263_, _14242_, _13676_);
  nand (_14264_, _14263_, _13621_);
  not (_14266_, _14263_);
  nand (_14267_, _14266_, _20050_);
  nand (_20060_, _14267_, _14264_);
  nor (_14268_, _14242_, _13682_);
  nand (_14269_, _14268_, _13621_);
  not (_14270_, _14268_);
  nand (_14271_, _14270_, _20091_);
  nand (_20102_, _14271_, _14269_);
  nor (_14272_, _14242_, _13688_);
  nand (_14273_, _14272_, _13621_);
  not (_14274_, _14272_);
  nand (_14275_, _14274_, _20133_);
  nand (_20144_, _14275_, _14273_);
  nor (_14276_, _14242_, _13698_);
  nand (_14277_, _14276_, _13621_);
  not (_14278_, _14276_);
  nand (_14279_, _14278_, _20174_);
  nand (_20185_, _14279_, _14277_);
  nor (_14280_, _14242_, _13704_);
  nand (_14281_, _14280_, _13621_);
  not (_14282_, _14280_);
  nand (_14283_, _14282_, _20215_);
  nand (_20226_, _14283_, _14281_);
  nor (_14284_, _14242_, _13710_);
  nand (_14285_, _14284_, _13621_);
  not (_14286_, _14284_);
  nand (_14287_, _14286_, _20256_);
  nand (_20267_, _14287_, _14285_);
  nor (_14288_, _14242_, _13716_);
  nand (_14289_, _14288_, _13621_);
  not (_14290_, _14288_);
  nand (_14291_, _14290_, _20298_);
  nand (_20308_, _14291_, _14289_);
  nor (_14292_, _14242_, _13724_);
  nand (_14293_, _14292_, _13621_);
  not (_14294_, _14292_);
  nand (_14295_, _14294_, _20339_);
  nand (_20350_, _14295_, _14293_);
  nor (_14296_, _14242_, _13731_);
  nand (_14297_, _14296_, _13621_);
  not (_14299_, _14296_);
  nand (_14300_, _14299_, _20380_);
  nand (_20391_, _14300_, _14297_);
  nor (_14301_, _14242_, _13737_);
  nand (_14302_, _14301_, _13621_);
  not (_14303_, _14301_);
  nand (_14304_, _14303_, _20421_);
  nand (_20432_, _14304_, _14302_);
  nor (_14305_, _14242_, _13743_);
  nand (_14306_, _14305_, _13621_);
  not (_14307_, _14305_);
  nand (_14308_, _14307_, _20462_);
  nand (_20473_, _14308_, _14306_);
  nor (_14309_, _13752_, _04274_);
  not (_14310_, _14309_);
  nor (_14311_, _14310_, _13749_);
  nand (_14312_, _14311_, _13621_);
  not (_14313_, _14311_);
  nand (_14314_, _14313_, _20512_);
  nand (_20522_, _14314_, _14312_);
  nor (_14315_, _14310_, _13641_);
  nand (_14316_, _14315_, _13621_);
  not (_14317_, _14315_);
  nand (_14318_, _14317_, _20553_);
  nand (_20563_, _14318_, _14316_);
  nor (_14319_, _14310_, _13650_);
  nand (_14320_, _14319_, _13621_);
  not (_14321_, _14319_);
  nand (_14322_, _14321_, _20593_);
  nand (_20604_, _14322_, _14320_);
  nor (_14323_, _14310_, _13659_);
  nand (_14324_, _14323_, _13621_);
  not (_14325_, _14323_);
  nand (_14326_, _14325_, _20633_);
  nand (_20644_, _14326_, _14324_);
  nor (_14327_, _14310_, _13670_);
  nand (_14328_, _14327_, _13621_);
  not (_14329_, _14327_);
  nand (_14330_, _14329_, _20674_);
  nand (_20684_, _14330_, _14328_);
  nor (_14332_, _14310_, _13676_);
  nand (_14333_, _14332_, _13621_);
  not (_14334_, _14332_);
  nand (_14335_, _14334_, _20714_);
  nand (_20724_, _14335_, _14333_);
  nor (_14336_, _14310_, _13682_);
  nand (_14337_, _14336_, _13621_);
  not (_14338_, _14336_);
  nand (_14339_, _14338_, _20754_);
  nand (_20765_, _14339_, _14337_);
  nor (_14340_, _14310_, _13688_);
  nand (_14341_, _14340_, _13621_);
  not (_14342_, _14340_);
  nand (_14343_, _14342_, _20793_);
  nand (_20804_, _14343_, _14341_);
  nor (_14344_, _14310_, _13698_);
  nand (_14345_, _14344_, _13621_);
  not (_14346_, _14344_);
  nand (_14347_, _14346_, _20832_);
  nand (_20842_, _14347_, _14345_);
  nor (_14348_, _14310_, _13704_);
  nand (_14349_, _14348_, _13621_);
  not (_14350_, _14348_);
  nand (_14351_, _14350_, _20871_);
  nand (_20881_, _14351_, _14349_);
  nor (_14352_, _14310_, _13710_);
  nand (_14353_, _14352_, _13621_);
  not (_14354_, _14352_);
  nand (_14355_, _14354_, _20909_);
  nand (_20920_, _14355_, _14353_);
  nor (_14356_, _14310_, _13716_);
  nand (_14357_, _14356_, _13621_);
  not (_14358_, _14356_);
  nand (_14359_, _14358_, _20950_);
  nand (_20960_, _14359_, _14357_);
  nor (_14360_, _14310_, _13724_);
  nand (_14361_, _14360_, _13621_);
  not (_14362_, _14360_);
  nand (_14363_, _14362_, _20989_);
  nand (_20999_, _14363_, _14361_);
  nor (_14365_, _14310_, _13731_);
  nand (_14366_, _14365_, _13621_);
  not (_14367_, _14365_);
  nand (_14368_, _14367_, _21028_);
  nand (_21038_, _14368_, _14366_);
  nor (_14369_, _14310_, _13737_);
  nand (_14370_, _14369_, _13621_);
  not (_14371_, _14369_);
  nand (_14372_, _14371_, _21067_);
  nand (_21077_, _14372_, _14370_);
  nor (_14373_, _14310_, _13743_);
  nand (_14374_, _14373_, _13621_);
  not (_14375_, _14373_);
  nand (_14376_, _14375_, _21106_);
  nand (_21116_, _14376_, _14374_);
  nor (_14377_, _14240_, _13823_);
  not (_14378_, _14377_);
  nor (_14379_, _14378_, _13749_);
  not (_14380_, _14379_);
  nand (_14381_, _14380_, _21154_);
  nand (_14382_, _14379_, _13621_);
  nand (_21164_, _14382_, _14381_);
  nor (_14383_, _14378_, _13641_);
  not (_14384_, _14383_);
  nand (_14385_, _14384_, _21193_);
  nand (_14386_, _14383_, _13621_);
  nand (_21203_, _14386_, _14385_);
  nor (_14387_, _14378_, _13650_);
  not (_14388_, _14387_);
  nand (_14389_, _14388_, _21232_);
  nand (_14390_, _14387_, _13621_);
  nand (_21242_, _14390_, _14389_);
  nor (_14391_, _14378_, _13659_);
  not (_14392_, _14391_);
  nand (_14393_, _14392_, _21271_);
  nand (_14394_, _14391_, _13621_);
  nand (_21281_, _14394_, _14393_);
  nor (_14395_, _14378_, _13670_);
  not (_14396_, _14395_);
  nand (_14397_, _14396_, _21310_);
  nand (_14399_, _14395_, _13621_);
  nand (_21321_, _14399_, _14397_);
  nor (_14400_, _14378_, _13676_);
  not (_14401_, _14400_);
  nand (_14402_, _14401_, _21350_);
  nand (_14403_, _14400_, _13621_);
  nand (_21360_, _14403_, _14402_);
  nor (_14404_, _14378_, _13682_);
  not (_14405_, _14404_);
  nand (_14406_, _14405_, _21388_);
  nand (_14407_, _14404_, _13621_);
  nand (_21399_, _14407_, _14406_);
  nor (_14408_, _14378_, _13688_);
  not (_14409_, _14408_);
  nand (_14410_, _14409_, _21427_);
  nand (_14411_, _14408_, _13621_);
  nand (_21437_, _14411_, _14410_);
  nor (_14412_, _14378_, _13698_);
  not (_14413_, _14412_);
  nand (_14414_, _14413_, _21466_);
  nand (_14415_, _14412_, _13621_);
  nand (_21476_, _14415_, _14414_);
  nor (_14416_, _14378_, _13704_);
  not (_14417_, _14416_);
  nand (_14418_, _14417_, _21504_);
  nand (_14419_, _14416_, _13621_);
  nand (_21515_, _14419_, _14418_);
  nor (_14420_, _14378_, _13710_);
  not (_14421_, _14420_);
  nand (_14422_, _14421_, _21543_);
  nand (_14423_, _14420_, _13621_);
  nand (_21553_, _14423_, _14422_);
  nor (_14424_, _14378_, _13716_);
  not (_14425_, _14424_);
  nand (_14426_, _14425_, _21582_);
  nand (_14427_, _14424_, _13621_);
  nand (_21592_, _14427_, _14426_);
  nor (_14428_, _14378_, _13724_);
  not (_14429_, _14428_);
  nand (_14430_, _14429_, _21620_);
  nand (_14432_, _14428_, _13621_);
  nand (_21631_, _14432_, _14430_);
  nor (_14433_, _14378_, _13731_);
  not (_14434_, _14433_);
  nand (_14435_, _14434_, _21659_);
  nand (_14436_, _14433_, _13621_);
  nand (_21669_, _14436_, _14435_);
  nor (_14437_, _14378_, _13737_);
  not (_14438_, _14437_);
  nand (_14439_, _14438_, _21698_);
  nand (_14440_, _14437_, _13621_);
  nand (_21709_, _14440_, _14439_);
  nor (_14441_, _14378_, _13743_);
  not (_14442_, _14441_);
  nand (_14443_, _14442_, _21737_);
  nand (_14444_, _14441_, _13621_);
  nand (_21748_, _14444_, _14443_);
  nor (_14445_, _13894_, _04274_);
  not (_14446_, _14445_);
  nor (_14447_, _14446_, _13749_);
  not (_14448_, _14447_);
  nand (_14449_, _14448_, _21786_);
  nand (_14450_, _14447_, _13621_);
  nand (_21796_, _14450_, _14449_);
  nor (_14451_, _14446_, _13641_);
  not (_14452_, _14451_);
  nand (_14453_, _14452_, _21825_);
  nand (_14454_, _14451_, _13621_);
  nand (_21835_, _14454_, _14453_);
  nor (_14455_, _14446_, _13650_);
  not (_14456_, _14455_);
  nand (_14457_, _14456_, _21863_);
  nand (_14458_, _14455_, _13621_);
  nand (_21874_, _14458_, _14457_);
  nor (_14459_, _14446_, _13659_);
  not (_14460_, _14459_);
  nand (_14461_, _14460_, _21902_);
  nand (_14462_, _14459_, _13621_);
  nand (_21912_, _14462_, _14461_);
  nor (_14463_, _14446_, _13670_);
  not (_14465_, _14463_);
  nand (_14466_, _14465_, _21941_);
  nand (_14467_, _14463_, _13621_);
  nand (_21951_, _14467_, _14466_);
  nor (_14468_, _14446_, _13676_);
  not (_14469_, _14468_);
  nand (_14470_, _14469_, _21980_);
  nand (_14471_, _14468_, _13621_);
  nand (_21990_, _14471_, _14470_);
  nor (_14472_, _14446_, _13682_);
  not (_14473_, _14472_);
  nand (_14474_, _14473_, _22018_);
  nand (_14475_, _14472_, _13621_);
  nand (_22029_, _14475_, _14474_);
  nor (_14476_, _14446_, _13688_);
  not (_14477_, _14476_);
  nand (_14478_, _14477_, _22058_);
  nand (_14479_, _14476_, _13621_);
  nand (_22069_, _14479_, _14478_);
  nor (_14480_, _14446_, _13698_);
  not (_14481_, _14480_);
  nand (_14482_, _14481_, _22101_);
  nand (_14483_, _14480_, _13621_);
  nand (_22112_, _14483_, _14482_);
  nor (_14484_, _14446_, _13704_);
  not (_14485_, _14484_);
  nand (_14486_, _14485_, _22143_);
  nand (_14487_, _14484_, _13621_);
  nand (_22154_, _14487_, _14486_);
  nor (_14488_, _14446_, _13710_);
  not (_14489_, _14488_);
  nand (_14490_, _14489_, _22185_);
  nand (_14491_, _14488_, _13621_);
  nand (_22196_, _14491_, _14490_);
  nor (_14492_, _14446_, _13716_);
  not (_14493_, _14492_);
  nand (_14494_, _14493_, _22227_);
  nand (_14495_, _14492_, _13621_);
  nand (_22238_, _14495_, _14494_);
  nor (_14496_, _14446_, _13724_);
  not (_14498_, _14496_);
  nand (_14499_, _14498_, _22269_);
  nand (_14500_, _14496_, _13621_);
  nand (_22280_, _14500_, _14499_);
  nor (_14501_, _14446_, _13731_);
  not (_14502_, _14501_);
  nand (_14503_, _14502_, _22311_);
  nand (_14504_, _14501_, _13621_);
  nand (_22322_, _14504_, _14503_);
  nor (_14505_, _14446_, _13737_);
  not (_14506_, _14505_);
  nand (_14507_, _14506_, _22353_);
  nand (_14508_, _14505_, _13621_);
  nand (_22364_, _14508_, _14507_);
  nor (_14509_, _14446_, _13743_);
  not (_14510_, _14509_);
  nand (_14511_, _14510_, _22395_);
  nand (_14512_, _14509_, _13621_);
  nand (_22406_, _14512_, _14511_);
  nor (_14513_, _01304_, _30882_);
  not (_14514_, _14513_);
  nor (_14515_, _14514_, _13625_);
  not (_14516_, _14515_);
  nor (_14517_, _14516_, _13749_);
  nand (_14518_, _14517_, _13621_);
  not (_14519_, _14517_);
  nand (_14520_, _14519_, _22457_);
  nand (_22468_, _14520_, _14518_);
  nor (_14521_, _14516_, _13641_);
  nand (_14522_, _14521_, _13621_);
  not (_14523_, _14521_);
  nand (_14524_, _14523_, _22499_);
  nand (_22510_, _14524_, _14522_);
  nor (_14525_, _14516_, _13650_);
  nand (_14526_, _14525_, _13621_);
  not (_14527_, _14525_);
  nand (_14528_, _14527_, _22542_);
  nand (_22553_, _14528_, _14526_);
  nor (_14529_, _14516_, _13659_);
  nand (_14530_, _14529_, _13621_);
  not (_14532_, _14529_);
  nand (_14533_, _14532_, _22584_);
  nand (_22595_, _14533_, _14530_);
  nor (_14534_, _14516_, _13670_);
  nand (_14535_, _14534_, _13621_);
  not (_14536_, _14534_);
  nand (_14537_, _14536_, _22626_);
  nand (_22637_, _14537_, _14535_);
  nor (_14538_, _14516_, _13676_);
  nand (_14539_, _14538_, _13621_);
  not (_14542_, _14538_);
  nand (_14543_, _14542_, _22668_);
  nand (_22679_, _14543_, _14539_);
  nor (_14544_, _14516_, _13682_);
  nand (_14545_, _14544_, _13621_);
  not (_14546_, _14544_);
  nand (_14547_, _14546_, _22710_);
  nand (_22721_, _14547_, _14545_);
  nor (_14548_, _14516_, _13688_);
  nand (_14549_, _14548_, _13621_);
  not (_14550_, _14548_);
  nand (_14551_, _14550_, _22752_);
  nand (_22763_, _14551_, _14549_);
  nor (_14552_, _14516_, _13698_);
  nand (_14553_, _14552_, _13621_);
  not (_14554_, _14552_);
  nand (_14555_, _14554_, _22794_);
  nand (_22805_, _14555_, _14553_);
  nor (_14556_, _14516_, _13704_);
  nand (_14557_, _14556_, _13621_);
  not (_14558_, _14556_);
  nand (_14559_, _14558_, _22836_);
  nand (_22847_, _14559_, _14557_);
  nor (_14560_, _14516_, _13710_);
  nand (_14561_, _14560_, _13621_);
  not (_14562_, _14560_);
  nand (_14563_, _14562_, _22878_);
  nand (_22889_, _14563_, _14561_);
  nor (_14564_, _14516_, _13716_);
  nand (_14565_, _14564_, _13621_);
  not (_14567_, _14564_);
  nand (_14568_, _14567_, _22920_);
  nand (_22931_, _14568_, _14565_);
  nor (_14569_, _14516_, _13724_);
  nand (_14570_, _14569_, _13621_);
  not (_14571_, _14569_);
  nand (_14572_, _14571_, _22963_);
  nand (_22974_, _14572_, _14570_);
  nor (_14573_, _14516_, _13731_);
  nand (_14574_, _14573_, _13621_);
  not (_14575_, _14573_);
  nand (_14576_, _14575_, _23005_);
  nand (_23016_, _14576_, _14574_);
  nor (_14577_, _14516_, _13737_);
  nand (_14578_, _14577_, _13621_);
  not (_14579_, _14577_);
  nand (_14580_, _14579_, _23047_);
  nand (_23058_, _14580_, _14578_);
  nor (_14581_, _14516_, _13743_);
  nand (_14582_, _14581_, _13621_);
  not (_14583_, _14581_);
  nand (_14584_, _14583_, _23089_);
  nand (_23100_, _14584_, _14582_);
  nor (_14585_, _13752_, _30882_);
  not (_14586_, _14585_);
  nor (_14587_, _14586_, _13749_);
  nand (_14588_, _14587_, _13621_);
  not (_14589_, _14587_);
  nand (_14590_, _14589_, _23141_);
  nand (_23152_, _14590_, _14588_);
  nor (_14591_, _14586_, _13641_);
  nand (_14592_, _14591_, _13621_);
  not (_14593_, _14591_);
  nand (_14594_, _14593_, _23183_);
  nand (_23194_, _14594_, _14592_);
  nor (_14595_, _14586_, _13650_);
  nand (_14596_, _14595_, _13621_);
  not (_14597_, _14595_);
  nand (_14598_, _14597_, _23225_);
  nand (_23236_, _14598_, _14596_);
  nor (_14600_, _14586_, _13659_);
  nand (_14601_, _14600_, _13621_);
  not (_14602_, _14600_);
  nand (_14603_, _14602_, _23258_);
  nand (_23259_, _14603_, _14601_);
  nor (_14604_, _14586_, _13670_);
  nand (_14605_, _14604_, _13621_);
  not (_14606_, _14604_);
  nand (_14607_, _14606_, _23260_);
  nand (_23261_, _14607_, _14605_);
  nor (_14608_, _14586_, _13676_);
  nand (_14609_, _14608_, _13621_);
  not (_14610_, _14608_);
  nand (_14611_, _14610_, _23262_);
  nand (_23264_, _14611_, _14609_);
  nor (_14612_, _14586_, _13682_);
  nand (_14613_, _14612_, _13621_);
  not (_14614_, _14612_);
  nand (_14615_, _14614_, _23265_);
  nand (_23266_, _14615_, _14613_);
  nor (_14616_, _14586_, _13688_);
  nand (_14617_, _14616_, _13621_);
  not (_14618_, _14616_);
  nand (_14619_, _14618_, _23267_);
  nand (_23268_, _14619_, _14617_);
  nor (_14620_, _14586_, _13698_);
  nand (_14621_, _14620_, _13621_);
  not (_14622_, _14620_);
  nand (_14623_, _14622_, _23269_);
  nand (_23270_, _14623_, _14621_);
  nor (_14624_, _14586_, _13704_);
  nand (_14625_, _14624_, _13621_);
  not (_14626_, _14624_);
  nand (_14627_, _14626_, _23271_);
  nand (_23272_, _14627_, _14625_);
  nor (_14628_, _14586_, _13710_);
  nand (_14629_, _14628_, _13621_);
  not (_14630_, _14628_);
  nand (_14631_, _14630_, _23273_);
  nand (_23274_, _14631_, _14629_);
  nor (_14633_, _14586_, _13716_);
  nand (_14634_, _14633_, _13621_);
  not (_14635_, _14633_);
  nand (_14636_, _14635_, _23275_);
  nand (_23276_, _14636_, _14634_);
  nor (_14637_, _14586_, _13724_);
  nand (_14638_, _14637_, _13621_);
  not (_14639_, _14637_);
  nand (_14640_, _14639_, _23277_);
  nand (_23278_, _14640_, _14638_);
  nor (_14641_, _14586_, _13731_);
  nand (_14642_, _14641_, _13621_);
  not (_14643_, _14641_);
  nand (_14644_, _14643_, _23279_);
  nand (_23280_, _14644_, _14642_);
  nor (_14645_, _14586_, _13737_);
  nand (_14646_, _14645_, _13621_);
  not (_14647_, _14645_);
  nand (_14648_, _14647_, _23281_);
  nand (_23282_, _14648_, _14646_);
  nor (_14649_, _14586_, _13743_);
  nand (_14650_, _14649_, _13621_);
  not (_14651_, _14649_);
  nand (_14652_, _14651_, _23283_);
  nand (_23285_, _14652_, _14650_);
  nor (_14653_, _14514_, _13823_);
  not (_14654_, _14653_);
  nor (_14655_, _14654_, _13749_);
  not (_14656_, _14655_);
  nand (_14657_, _14656_, _23286_);
  nand (_14658_, _14655_, _13621_);
  nand (_23287_, _14658_, _14657_);
  nor (_14659_, _14654_, _13641_);
  not (_14660_, _14659_);
  nand (_14661_, _14660_, _23288_);
  nand (_14662_, _14659_, _13621_);
  nand (_23289_, _14662_, _14661_);
  nor (_14663_, _14654_, _13650_);
  not (_14664_, _14663_);
  nand (_14665_, _14664_, _23290_);
  nand (_14667_, _14663_, _13621_);
  nand (_23291_, _14667_, _14665_);
  nor (_14668_, _14654_, _13659_);
  not (_14669_, _14668_);
  nand (_14670_, _14669_, _23292_);
  nand (_14671_, _14668_, _13621_);
  nand (_23293_, _14671_, _14670_);
  nor (_14672_, _14654_, _13670_);
  not (_14673_, _14672_);
  nand (_14674_, _14673_, _23294_);
  nand (_14675_, _14672_, _13621_);
  nand (_23295_, _14675_, _14674_);
  nor (_14676_, _14654_, _13676_);
  not (_14677_, _14676_);
  nand (_14678_, _14677_, _23296_);
  nand (_14679_, _14676_, _13621_);
  nand (_23297_, _14679_, _14678_);
  nor (_14680_, _14654_, _13682_);
  not (_14681_, _14680_);
  nand (_14682_, _14681_, _23298_);
  nand (_14683_, _14680_, _13621_);
  nand (_23299_, _14683_, _14682_);
  nor (_14684_, _14654_, _13688_);
  not (_14685_, _14684_);
  nand (_14686_, _14685_, _23300_);
  nand (_14687_, _14684_, _13621_);
  nand (_23301_, _14687_, _14686_);
  nor (_14688_, _14654_, _13698_);
  not (_14689_, _14688_);
  nand (_14690_, _14689_, _23302_);
  nand (_14691_, _14688_, _13621_);
  nand (_23303_, _14691_, _14690_);
  nor (_14692_, _14654_, _13704_);
  not (_14693_, _14692_);
  nand (_14694_, _14693_, _23305_);
  nand (_14695_, _14692_, _13621_);
  nand (_23306_, _14695_, _14694_);
  nor (_14696_, _14654_, _13710_);
  not (_14697_, _14696_);
  nand (_14698_, _14697_, _23307_);
  nand (_14700_, _14696_, _13621_);
  nand (_23308_, _14700_, _14698_);
  nor (_14701_, _14654_, _13716_);
  not (_14702_, _14701_);
  nand (_14703_, _14702_, _23309_);
  nand (_14704_, _14701_, _13621_);
  nand (_23310_, _14704_, _14703_);
  nor (_14705_, _14654_, _13724_);
  not (_14706_, _14705_);
  nand (_14707_, _14706_, _23311_);
  nand (_14708_, _14705_, _13621_);
  nand (_23312_, _14708_, _14707_);
  nor (_14709_, _14654_, _13731_);
  not (_14710_, _14709_);
  nand (_14711_, _14710_, _23313_);
  nand (_14712_, _14709_, _13621_);
  nand (_23314_, _14712_, _14711_);
  nor (_14713_, _14654_, _13737_);
  not (_14714_, _14713_);
  nand (_14715_, _14714_, _23315_);
  nand (_14716_, _14713_, _13621_);
  nand (_23316_, _14716_, _14715_);
  nor (_14717_, _14654_, _13743_);
  not (_14718_, _14717_);
  nand (_14719_, _14718_, _23317_);
  nand (_14720_, _14717_, _13621_);
  nand (_23318_, _14720_, _14719_);
  nor (_14721_, _13894_, _30882_);
  not (_14722_, _14721_);
  nor (_14723_, _14722_, _13749_);
  nand (_14724_, _14723_, _13621_);
  not (_14725_, _14723_);
  nand (_14726_, _14725_, _23319_);
  nand (_23320_, _14726_, _14724_);
  nor (_14727_, _14722_, _13641_);
  nand (_14728_, _14727_, _13621_);
  not (_14729_, _14727_);
  nand (_14730_, _14729_, _23321_);
  nand (_23322_, _14730_, _14728_);
  nor (_14731_, _14722_, _13650_);
  nand (_14733_, _14731_, _13621_);
  not (_14734_, _14731_);
  nand (_14735_, _14734_, _23323_);
  nand (_23324_, _14735_, _14733_);
  nor (_14736_, _14722_, _13659_);
  nand (_14737_, _14736_, _13621_);
  not (_14738_, _14736_);
  nand (_14739_, _14738_, _23326_);
  nand (_23327_, _14739_, _14737_);
  nor (_14740_, _14722_, _13670_);
  nand (_14741_, _14740_, _13621_);
  not (_14742_, _14740_);
  nand (_14743_, _14742_, _23328_);
  nand (_23329_, _14743_, _14741_);
  nor (_14744_, _14722_, _13676_);
  nand (_14745_, _14744_, _13621_);
  not (_14746_, _14744_);
  nand (_14747_, _14746_, _23330_);
  nand (_23331_, _14747_, _14745_);
  nor (_14748_, _14722_, _13682_);
  nand (_14749_, _14748_, _13621_);
  not (_14750_, _14748_);
  nand (_14751_, _14750_, _23332_);
  nand (_23333_, _14751_, _14749_);
  nor (_14752_, _14722_, _13688_);
  nand (_14753_, _14752_, _13621_);
  not (_14754_, _14752_);
  nand (_14755_, _14754_, _23334_);
  nand (_23335_, _14755_, _14753_);
  nor (_14756_, _14722_, _13698_);
  nand (_14757_, _14756_, _13621_);
  not (_14758_, _14756_);
  nand (_14759_, _14758_, _23336_);
  nand (_23337_, _14759_, _14757_);
  nor (_14760_, _14722_, _13704_);
  nand (_14761_, _14760_, _13621_);
  not (_14762_, _14760_);
  nand (_14763_, _14762_, _23338_);
  nand (_23339_, _14763_, _14761_);
  nor (_14764_, _14722_, _13710_);
  nand (_14766_, _14764_, _13621_);
  not (_14767_, _14764_);
  nand (_14768_, _14767_, _23340_);
  nand (_23341_, _14768_, _14766_);
  nor (_14769_, _14722_, _13716_);
  nand (_14770_, _14769_, _13621_);
  not (_14771_, _14769_);
  nand (_14772_, _14771_, _23342_);
  nand (_23343_, _14772_, _14770_);
  nor (_14773_, _14722_, _13724_);
  nand (_14774_, _14773_, _13621_);
  not (_14775_, _14773_);
  nand (_14776_, _14775_, _23344_);
  nand (_23345_, _14776_, _14774_);
  nor (_14777_, _14722_, _13731_);
  nand (_14778_, _14777_, _13621_);
  not (_14779_, _14777_);
  nand (_14780_, _14779_, _23348_);
  nand (_23349_, _14780_, _14778_);
  nor (_14781_, _14722_, _13737_);
  nand (_14782_, _14781_, _13621_);
  not (_14783_, _14781_);
  nand (_14784_, _14783_, _23350_);
  nand (_23351_, _14784_, _14782_);
  nor (_14785_, _14722_, _13743_);
  nand (_14786_, _14785_, _13621_);
  not (_14787_, _14785_);
  nand (_14788_, _14787_, _23352_);
  nand (_23353_, _14788_, _14786_);
  nor (_14789_, _01136_, _01304_);
  nand (_14790_, _13776_, _14789_);
  nand (_14791_, _13778_, _23354_);
  nand (_23355_, _14791_, _14790_);
  nor (_14792_, _01128_, _01304_);
  nand (_14793_, _14792_, _13776_);
  nand (_14794_, _13778_, _23356_);
  nand (_23357_, _14794_, _14793_);
  nor (_14795_, _01120_, _01304_);
  nand (_14796_, _14795_, _13776_);
  nand (_14797_, _13778_, _23358_);
  nand (_23359_, _14797_, _14796_);
  nor (_14799_, _01110_, _01304_);
  nand (_14800_, _14799_, _13776_);
  nand (_14801_, _13778_, _23360_);
  nand (_23361_, _14801_, _14800_);
  nor (_14802_, _01100_, _01304_);
  nand (_14803_, _14802_, _13776_);
  nand (_14804_, _13778_, _23362_);
  nand (_23363_, _14804_, _14803_);
  nor (_14805_, _01093_, _01304_);
  nand (_14806_, _14805_, _13776_);
  nand (_14807_, _13778_, _23364_);
  nand (_23365_, _14807_, _14806_);
  nor (_14808_, _01085_, _01304_);
  nand (_14809_, _14808_, _13776_);
  nand (_14810_, _13778_, _23366_);
  nand (_23367_, _14810_, _14809_);
  nand (_14811_, _13772_, _14789_);
  nand (_14812_, _13774_, _23368_);
  nand (_23369_, _14812_, _14811_);
  nand (_14813_, _14792_, _13772_);
  nand (_14814_, _13774_, _23370_);
  nand (_23371_, _14814_, _14813_);
  nand (_14815_, _14795_, _13772_);
  nand (_14816_, _13774_, _23372_);
  nand (_23373_, _14816_, _14815_);
  nand (_14817_, _14799_, _13772_);
  nand (_14818_, _13774_, _23374_);
  nand (_23375_, _14818_, _14817_);
  nand (_14819_, _14802_, _13772_);
  nand (_14820_, _13774_, _23377_);
  nand (_23378_, _14820_, _14819_);
  nand (_14821_, _14805_, _13772_);
  nand (_14822_, _13774_, _23379_);
  nand (_23380_, _14822_, _14821_);
  nand (_14823_, _14808_, _13772_);
  nand (_14824_, _13774_, _23381_);
  nand (_23382_, _14824_, _14823_);
  nand (_14825_, _13768_, _14789_);
  nand (_14826_, _13770_, _23383_);
  nand (_23384_, _14826_, _14825_);
  nand (_14828_, _14792_, _13768_);
  nand (_14829_, _13770_, _23385_);
  nand (_23386_, _14829_, _14828_);
  nand (_14830_, _14795_, _13768_);
  nand (_14831_, _13770_, _23387_);
  nand (_23388_, _14831_, _14830_);
  nand (_14832_, _14799_, _13768_);
  nand (_14833_, _13770_, _23389_);
  nand (_23390_, _14833_, _14832_);
  nand (_14834_, _14802_, _13768_);
  nand (_14835_, _13770_, _23391_);
  nand (_23392_, _14835_, _14834_);
  nand (_14836_, _14805_, _13768_);
  nand (_14837_, _13770_, _23393_);
  nand (_23394_, _14837_, _14836_);
  nand (_14838_, _14808_, _13768_);
  nand (_14839_, _13770_, _23395_);
  nand (_23396_, _14839_, _14838_);
  nand (_14840_, _13764_, _14789_);
  nand (_14841_, _13766_, _23397_);
  nand (_23398_, _14841_, _14840_);
  nand (_14842_, _14792_, _13764_);
  nand (_14843_, _13766_, _23399_);
  nand (_23400_, _14843_, _14842_);
  nand (_14844_, _14795_, _13764_);
  nand (_14845_, _13766_, _23401_);
  nand (_23402_, _14845_, _14844_);
  nand (_14846_, _14799_, _13764_);
  nand (_14847_, _13766_, _23403_);
  nand (_23404_, _14847_, _14846_);
  nand (_14848_, _14802_, _13764_);
  nand (_14849_, _13766_, _23405_);
  nand (_23406_, _14849_, _14848_);
  nand (_14850_, _14805_, _13764_);
  nand (_14851_, _13766_, _23407_);
  nand (_23408_, _14851_, _14850_);
  nand (_14852_, _14808_, _13764_);
  nand (_14853_, _13766_, _23409_);
  nand (_23410_, _14853_, _14852_);
  nand (_14855_, _13759_, _14789_);
  nand (_14856_, _13761_, _23411_);
  nand (_23412_, _14856_, _14855_);
  nand (_14857_, _14792_, _13759_);
  nand (_14858_, _13761_, _23413_);
  nand (_23414_, _14858_, _14857_);
  nand (_14859_, _14795_, _13759_);
  nand (_14860_, _13761_, _23415_);
  nand (_23416_, _14860_, _14859_);
  nand (_14861_, _14799_, _13759_);
  nand (_14863_, _13761_, _23418_);
  nand (_23419_, _14863_, _14861_);
  nand (_14864_, _14802_, _13759_);
  nand (_14865_, _13761_, _23420_);
  nand (_23421_, _14865_, _14864_);
  nand (_14866_, _14805_, _13759_);
  nand (_14867_, _13761_, _23422_);
  nand (_23423_, _14867_, _14866_);
  nand (_14868_, _14808_, _13759_);
  nand (_14869_, _13761_, _23424_);
  nand (_23425_, _14869_, _14868_);
  nand (_14870_, _13755_, _14789_);
  nand (_14871_, _13757_, _23426_);
  nand (_23427_, _14871_, _14870_);
  nand (_14872_, _14792_, _13755_);
  nand (_14873_, _13757_, _23428_);
  nand (_23429_, _14873_, _14872_);
  nand (_14874_, _14795_, _13755_);
  nand (_14875_, _13757_, _23430_);
  nand (_23431_, _14875_, _14874_);
  nand (_14876_, _14799_, _13755_);
  nand (_14877_, _13757_, _23432_);
  nand (_23433_, _14877_, _14876_);
  nand (_14878_, _14802_, _13755_);
  nand (_14879_, _13757_, _23434_);
  nand (_23435_, _14879_, _14878_);
  nand (_14880_, _14805_, _13755_);
  nand (_14881_, _13757_, _23436_);
  nand (_23437_, _14881_, _14880_);
  nand (_14882_, _14808_, _13755_);
  nand (_14884_, _13757_, _23438_);
  nand (_23439_, _14884_, _14882_);
  nand (_14885_, _13744_, _14789_);
  nand (_14886_, _13746_, _23440_);
  nand (_23441_, _14886_, _14885_);
  nand (_14887_, _14792_, _13744_);
  nand (_14888_, _13746_, _23442_);
  nand (_23443_, _14888_, _14887_);
  nand (_14889_, _14795_, _13744_);
  nand (_14890_, _13746_, _23444_);
  nand (_23445_, _14890_, _14889_);
  nand (_14891_, _14799_, _13744_);
  nand (_14892_, _13746_, _23446_);
  nand (_23447_, _14892_, _14891_);
  nand (_14893_, _14802_, _13744_);
  nand (_14894_, _13746_, _23448_);
  nand (_23449_, _14894_, _14893_);
  nand (_14895_, _14805_, _13744_);
  nand (_14896_, _13746_, _23450_);
  nand (_23451_, _14896_, _14895_);
  nand (_14897_, _14808_, _13744_);
  nand (_14898_, _13746_, _23452_);
  nand (_23453_, _14898_, _14897_);
  nand (_14899_, _13738_, _14789_);
  nand (_14900_, _13740_, _23454_);
  nand (_23455_, _14900_, _14899_);
  nand (_14901_, _14792_, _13738_);
  nand (_14902_, _13740_, _23456_);
  nand (_23457_, _14902_, _14901_);
  nand (_14903_, _14795_, _13738_);
  nand (_14904_, _13740_, _23459_);
  nand (_23460_, _14904_, _14903_);
  nand (_14905_, _14799_, _13738_);
  nand (_14906_, _13740_, _23461_);
  nand (_23462_, _14906_, _14905_);
  nand (_14907_, _14802_, _13738_);
  nand (_14908_, _13740_, _23463_);
  nand (_23464_, _14908_, _14907_);
  nand (_14909_, _14805_, _13738_);
  nand (_14910_, _13740_, _23465_);
  nand (_23466_, _14910_, _14909_);
  nand (_14912_, _14808_, _13738_);
  nand (_14913_, _13740_, _23467_);
  nand (_23468_, _14913_, _14912_);
  nand (_14914_, _13732_, _14789_);
  nand (_14915_, _13734_, _23469_);
  nand (_23470_, _14915_, _14914_);
  nand (_14916_, _14792_, _13732_);
  nand (_14917_, _13734_, _23471_);
  nand (_23472_, _14917_, _14916_);
  nand (_14918_, _14795_, _13732_);
  nand (_14919_, _13734_, _23473_);
  nand (_23474_, _14919_, _14918_);
  nand (_14920_, _14799_, _13732_);
  nand (_14921_, _13734_, _23475_);
  nand (_23476_, _14921_, _14920_);
  nand (_14922_, _14802_, _13732_);
  nand (_14923_, _13734_, _23477_);
  nand (_23478_, _14923_, _14922_);
  nand (_14924_, _14805_, _13732_);
  nand (_14925_, _13734_, _23479_);
  nand (_23480_, _14925_, _14924_);
  nand (_14926_, _14808_, _13732_);
  nand (_14927_, _13734_, _23481_);
  nand (_23482_, _14927_, _14926_);
  nand (_14928_, _13725_, _14789_);
  nand (_14929_, _13727_, _23483_);
  nand (_23484_, _14929_, _14928_);
  nand (_14930_, _14792_, _13725_);
  nand (_14931_, _13727_, _23485_);
  nand (_23486_, _14931_, _14930_);
  nand (_14932_, _14795_, _13725_);
  nand (_14933_, _13727_, _23487_);
  nand (_23488_, _14933_, _14932_);
  nand (_14934_, _14799_, _13725_);
  nand (_14935_, _13727_, _23489_);
  nand (_23490_, _14935_, _14934_);
  nand (_14936_, _14802_, _13725_);
  nand (_14937_, _13727_, _23491_);
  nand (_23492_, _14937_, _14936_);
  nand (_14939_, _14805_, _13725_);
  nand (_14940_, _13727_, _23493_);
  nand (_23494_, _14940_, _14939_);
  nand (_14941_, _14808_, _13725_);
  nand (_14942_, _13727_, _23495_);
  nand (_23496_, _14942_, _14941_);
  nand (_14943_, _13717_, _14789_);
  nand (_14944_, _13719_, _23497_);
  nand (_23498_, _14944_, _14943_);
  nand (_14945_, _14792_, _13717_);
  nand (_14946_, _13719_, _23500_);
  nand (_23501_, _14946_, _14945_);
  nand (_14947_, _14795_, _13717_);
  nand (_14948_, _13719_, _23502_);
  nand (_23503_, _14948_, _14947_);
  nand (_14949_, _14799_, _13717_);
  nand (_14950_, _13719_, _23504_);
  nand (_23505_, _14950_, _14949_);
  nand (_14951_, _14802_, _13717_);
  nand (_14952_, _13719_, _23506_);
  nand (_23507_, _14952_, _14951_);
  nand (_14953_, _14805_, _13717_);
  nand (_14954_, _13719_, _23508_);
  nand (_23509_, _14954_, _14953_);
  nand (_14955_, _14808_, _13717_);
  nand (_14956_, _13719_, _23510_);
  nand (_23511_, _14956_, _14955_);
  nand (_14957_, _13797_, _14789_);
  nand (_14958_, _13799_, _23512_);
  nand (_23513_, _14958_, _14957_);
  nand (_14959_, _14792_, _13797_);
  nand (_14960_, _13799_, _23514_);
  nand (_23515_, _14960_, _14959_);
  nand (_14961_, _14795_, _13797_);
  nand (_14962_, _13799_, _23516_);
  nand (_23517_, _14962_, _14961_);
  nand (_14963_, _14799_, _13797_);
  nand (_14964_, _13799_, _23518_);
  nand (_23519_, _14964_, _14963_);
  nand (_14965_, _14802_, _13797_);
  nand (_14967_, _13799_, _23520_);
  nand (_23521_, _14967_, _14965_);
  nand (_14968_, _14805_, _13797_);
  nand (_14969_, _13799_, _23522_);
  nand (_23523_, _14969_, _14968_);
  nand (_14970_, _14808_, _13797_);
  nand (_14971_, _13799_, _23524_);
  nand (_23525_, _14971_, _14970_);
  nand (_14972_, _13792_, _14789_);
  nand (_14973_, _13794_, _23526_);
  nand (_23527_, _14973_, _14972_);
  nand (_14974_, _14792_, _13792_);
  nand (_14975_, _13794_, _23528_);
  nand (_23529_, _14975_, _14974_);
  nand (_14976_, _14795_, _13792_);
  nand (_14977_, _13794_, _23530_);
  nand (_23531_, _14977_, _14976_);
  nand (_14978_, _14799_, _13792_);
  nand (_14979_, _13794_, _23532_);
  nand (_23533_, _14979_, _14978_);
  nand (_14980_, _14802_, _13792_);
  nand (_14981_, _13794_, _23534_);
  nand (_23535_, _14981_, _14980_);
  nand (_14982_, _14805_, _13792_);
  nand (_14983_, _13794_, _23536_);
  nand (_23537_, _14983_, _14982_);
  nand (_14984_, _14808_, _13792_);
  nand (_14985_, _13794_, _23538_);
  nand (_23539_, _14985_, _14984_);
  nand (_14986_, _13817_, _14789_);
  nand (_14987_, _13819_, _23541_);
  nand (_23542_, _14987_, _14986_);
  nand (_14988_, _14792_, _13817_);
  nand (_14989_, _13819_, _23543_);
  nand (_23544_, _14989_, _14988_);
  nand (_14990_, _14795_, _13817_);
  nand (_14991_, _13819_, _23545_);
  nand (_23546_, _14991_, _14990_);
  nand (_14992_, _14799_, _13817_);
  nand (_14993_, _13819_, _23547_);
  nand (_23548_, _14993_, _14992_);
  nand (_14995_, _14802_, _13817_);
  nand (_14996_, _13819_, _23549_);
  nand (_23550_, _14996_, _14995_);
  nand (_14997_, _14805_, _13817_);
  nand (_14998_, _13819_, _23551_);
  nand (_23552_, _14998_, _14997_);
  nand (_14999_, _14808_, _13817_);
  nand (_15000_, _13819_, _23553_);
  nand (_23554_, _15000_, _14999_);
  nand (_15001_, _13831_, _14789_);
  nand (_15002_, _13833_, _23555_);
  nand (_23556_, _15002_, _15001_);
  nand (_15003_, _14792_, _13831_);
  nand (_15004_, _13833_, _23557_);
  nand (_23558_, _15004_, _15003_);
  nand (_15005_, _14795_, _13831_);
  nand (_15006_, _13833_, _23559_);
  nand (_23560_, _15006_, _15005_);
  nand (_15007_, _14799_, _13831_);
  nand (_15008_, _13833_, _23561_);
  nand (_23562_, _15008_, _15007_);
  nand (_15009_, _14802_, _13831_);
  nand (_15010_, _13833_, _23563_);
  nand (_23564_, _15010_, _15009_);
  nand (_15011_, _14805_, _13831_);
  nand (_15012_, _13833_, _23565_);
  nand (_23566_, _15012_, _15011_);
  nand (_15013_, _14808_, _13831_);
  nand (_15014_, _13833_, _23567_);
  nand (_23568_, _15014_, _15013_);
  nand (_15015_, _13839_, _14789_);
  nand (_15016_, _13841_, _23569_);
  nand (_23570_, _15016_, _15015_);
  nand (_15017_, _14792_, _13839_);
  nand (_15018_, _13841_, _23571_);
  nand (_23572_, _15018_, _15017_);
  nand (_15019_, _14795_, _13839_);
  nand (_15020_, _13841_, _23573_);
  nand (_23574_, _15020_, _15019_);
  nand (_15022_, _14799_, _13839_);
  nand (_15023_, _13841_, _23575_);
  nand (_23576_, _15023_, _15022_);
  nand (_15024_, _14802_, _13839_);
  nand (_15025_, _13841_, _23577_);
  nand (_23578_, _15025_, _15024_);
  nand (_15026_, _14805_, _13839_);
  nand (_15027_, _13841_, _23579_);
  nand (_23580_, _15027_, _15026_);
  nand (_15028_, _14808_, _13839_);
  nand (_15029_, _13841_, _23582_);
  nand (_23583_, _15029_, _15028_);
  nand (_15030_, _13877_, _14789_);
  nand (_15031_, _13879_, _23584_);
  nand (_23585_, _15031_, _15030_);
  nand (_15032_, _14792_, _13877_);
  nand (_15033_, _13879_, _23586_);
  nand (_23587_, _15033_, _15032_);
  nand (_15034_, _14795_, _13877_);
  nand (_15035_, _13879_, _23588_);
  nand (_23589_, _15035_, _15034_);
  nand (_15036_, _14799_, _13877_);
  nand (_15037_, _13879_, _23590_);
  nand (_23591_, _15037_, _15036_);
  nand (_15038_, _14802_, _13877_);
  nand (_15039_, _13879_, _23592_);
  nand (_23593_, _15039_, _15038_);
  nand (_15040_, _14805_, _13877_);
  nand (_15041_, _13879_, _23594_);
  nand (_23595_, _15041_, _15040_);
  nand (_15042_, _14808_, _13877_);
  nand (_15043_, _13879_, _23596_);
  nand (_23597_, _15043_, _15042_);
  nand (_15044_, _13910_, _14789_);
  nand (_15045_, _13912_, _23598_);
  nand (_23599_, _15045_, _15044_);
  nand (_15046_, _14792_, _13910_);
  nand (_15047_, _13912_, _23600_);
  nand (_23601_, _15047_, _15046_);
  nand (_15048_, _14795_, _13910_);
  nand (_15050_, _13912_, _23602_);
  nand (_23603_, _15050_, _15048_);
  nand (_15051_, _14799_, _13910_);
  nand (_15052_, _13912_, _23604_);
  nand (_23605_, _15052_, _15051_);
  nand (_15053_, _14802_, _13910_);
  nand (_15054_, _13912_, _23606_);
  nand (_23607_, _15054_, _15053_);
  nand (_15055_, _14805_, _13910_);
  nand (_15056_, _13912_, _23608_);
  nand (_23609_, _15056_, _15055_);
  nand (_15057_, _14808_, _13910_);
  nand (_15058_, _13912_, _23610_);
  nand (_23611_, _15058_, _15057_);
  nand (_15059_, _13918_, _14789_);
  nand (_15060_, _13920_, _23612_);
  nand (_23613_, _15060_, _15059_);
  nand (_15061_, _14792_, _13918_);
  nand (_15062_, _13920_, _23614_);
  nand (_23615_, _15062_, _15061_);
  nand (_15063_, _14795_, _13918_);
  nand (_15064_, _13920_, _23616_);
  nand (_23617_, _15064_, _15063_);
  nand (_15065_, _14799_, _13918_);
  nand (_15066_, _13920_, _23618_);
  nand (_23619_, _15066_, _15065_);
  nand (_15067_, _14802_, _13918_);
  nand (_15068_, _13920_, _23620_);
  nand (_23621_, _15068_, _15067_);
  nand (_15069_, _14805_, _13918_);
  nand (_15070_, _13920_, _23623_);
  nand (_23624_, _15070_, _15069_);
  nand (_15071_, _14808_, _13918_);
  nand (_15072_, _13920_, _23625_);
  nand (_23626_, _15072_, _15071_);
  nand (_15073_, _14365_, _14789_);
  nand (_15074_, _14367_, _23627_);
  nand (_23628_, _15074_, _15073_);
  nand (_15075_, _14792_, _14365_);
  nand (_15076_, _14367_, _23629_);
  nand (_23630_, _15076_, _15075_);
  nand (_15078_, _14795_, _14365_);
  nand (_15079_, _14367_, _23631_);
  nand (_23632_, _15079_, _15078_);
  nand (_15080_, _14799_, _14365_);
  nand (_15081_, _14367_, _23633_);
  nand (_23634_, _15081_, _15080_);
  nand (_15082_, _14802_, _14365_);
  nand (_15083_, _14367_, _23635_);
  nand (_23636_, _15083_, _15082_);
  nand (_15084_, _14805_, _14365_);
  nand (_15085_, _14367_, _23637_);
  nand (_23638_, _15085_, _15084_);
  nand (_15086_, _14808_, _14365_);
  nand (_15087_, _14367_, _23639_);
  nand (_23640_, _15087_, _15086_);
  nand (_15088_, _14360_, _14789_);
  nand (_15089_, _14362_, _23641_);
  nand (_23642_, _15089_, _15088_);
  nand (_15090_, _14792_, _14360_);
  nand (_15091_, _14362_, _23643_);
  nand (_23644_, _15091_, _15090_);
  nand (_15092_, _14795_, _14360_);
  nand (_15093_, _14362_, _23645_);
  nand (_23646_, _15093_, _15092_);
  nand (_15094_, _14799_, _14360_);
  nand (_15095_, _14362_, _23647_);
  nand (_23648_, _15095_, _15094_);
  nand (_15096_, _14802_, _14360_);
  nand (_15097_, _14362_, _23649_);
  nand (_23650_, _15097_, _15096_);
  nand (_15098_, _14805_, _14360_);
  nand (_15099_, _14362_, _23651_);
  nand (_23652_, _15099_, _15098_);
  nand (_15100_, _14808_, _14360_);
  nand (_15101_, _14362_, _23653_);
  nand (_23654_, _15101_, _15100_);
  nand (_15102_, _14369_, _14789_);
  nand (_15103_, _14371_, _23655_);
  nand (_23656_, _15103_, _15102_);
  nand (_15105_, _14792_, _14369_);
  nand (_15106_, _14371_, _23657_);
  nand (_23658_, _15106_, _15105_);
  nand (_15107_, _14795_, _14369_);
  nand (_15108_, _14371_, _23659_);
  nand (_23660_, _15108_, _15107_);
  nand (_15109_, _14799_, _14369_);
  nand (_15110_, _14371_, _23661_);
  nand (_23662_, _15110_, _15109_);
  nand (_15111_, _14802_, _14369_);
  nand (_15112_, _14371_, _23664_);
  nand (_23665_, _15112_, _15111_);
  nand (_15113_, _14805_, _14369_);
  nand (_15114_, _14371_, _23666_);
  nand (_23667_, _15114_, _15113_);
  nand (_15115_, _14808_, _14369_);
  nand (_15116_, _14371_, _23668_);
  nand (_23669_, _15116_, _15115_);
  nand (_15117_, _14356_, _14789_);
  nand (_15118_, _14358_, _23670_);
  nand (_23671_, _15118_, _15117_);
  nand (_15119_, _14792_, _14356_);
  nand (_15120_, _14358_, _23672_);
  nand (_23673_, _15120_, _15119_);
  nand (_15121_, _14795_, _14356_);
  nand (_15122_, _14358_, _23674_);
  nand (_23675_, _15122_, _15121_);
  nand (_15123_, _14799_, _14356_);
  nand (_15124_, _14358_, _23676_);
  nand (_23677_, _15124_, _15123_);
  nand (_15125_, _14802_, _14356_);
  nand (_15126_, _14358_, _23678_);
  nand (_23679_, _15126_, _15125_);
  nand (_15127_, _14805_, _14356_);
  nand (_15128_, _14358_, _23680_);
  nand (_23681_, _15128_, _15127_);
  nand (_15129_, _14808_, _14356_);
  nand (_15130_, _14358_, _23682_);
  nand (_23683_, _15130_, _15129_);
  nand (_15131_, _13914_, _14789_);
  nand (_15133_, _13916_, _23692_);
  nand (_23693_, _15133_, _15131_);
  nand (_15134_, _14792_, _13914_);
  nand (_15135_, _13916_, _23694_);
  nand (_23695_, _15135_, _15134_);
  nand (_15136_, _14795_, _13914_);
  nand (_15137_, _13916_, _23696_);
  nand (_23697_, _15137_, _15136_);
  nand (_15138_, _14799_, _13914_);
  nand (_15139_, _13916_, _23701_);
  nand (_23702_, _15139_, _15138_);
  nand (_15141_, _14802_, _13914_);
  nand (_15142_, _13916_, _23703_);
  nand (_23704_, _15142_, _15141_);
  nand (_15143_, _14805_, _13914_);
  nand (_15144_, _13916_, _23705_);
  nand (_23706_, _15144_, _15143_);
  nand (_15145_, _14808_, _13914_);
  nand (_15146_, _13916_, _23707_);
  nand (_23708_, _15146_, _15145_);
  nand (_15147_, _14785_, _14789_);
  nand (_15148_, _14787_, _23709_);
  nand (_23710_, _15148_, _15147_);
  nand (_15149_, _14792_, _14785_);
  nand (_15150_, _14787_, _23711_);
  nand (_23712_, _15150_, _15149_);
  nand (_15151_, _14795_, _14785_);
  nand (_15152_, _14787_, _23713_);
  nand (_23714_, _15152_, _15151_);
  nand (_15153_, _14799_, _14785_);
  nand (_15154_, _14787_, _23715_);
  nand (_23716_, _15154_, _15153_);
  nand (_15155_, _14802_, _14785_);
  nand (_15156_, _14787_, _23717_);
  nand (_23718_, _15156_, _15155_);
  nand (_15157_, _14805_, _14785_);
  nand (_15158_, _14787_, _23719_);
  nand (_23720_, _15158_, _15157_);
  nand (_15159_, _14808_, _14785_);
  nand (_15160_, _14787_, _23721_);
  nand (_23722_, _15160_, _15159_);
  nand (_15162_, _14781_, _14789_);
  nand (_15163_, _14783_, _23723_);
  nand (_23724_, _15163_, _15162_);
  nand (_15164_, _14792_, _14781_);
  nand (_15165_, _14783_, _23725_);
  nand (_23726_, _15165_, _15164_);
  nand (_15166_, _14795_, _14781_);
  nand (_15167_, _14783_, _23727_);
  nand (_23728_, _15167_, _15166_);
  nand (_15168_, _14799_, _14781_);
  nand (_15169_, _14783_, _23729_);
  nand (_23730_, _15169_, _15168_);
  nand (_15170_, _14802_, _14781_);
  nand (_15171_, _14783_, _23731_);
  nand (_23732_, _15171_, _15170_);
  nand (_15172_, _14805_, _14781_);
  nand (_15173_, _14783_, _23733_);
  nand (_23734_, _15173_, _15172_);
  nand (_15174_, _14808_, _14781_);
  nand (_15175_, _14783_, _23735_);
  nand (_23736_, _15175_, _15174_);
  nand (_15176_, _14777_, _14789_);
  nand (_15177_, _14779_, _23737_);
  nand (_23738_, _15177_, _15176_);
  nand (_15178_, _14792_, _14777_);
  nand (_15179_, _14779_, _23739_);
  nand (_23740_, _15179_, _15178_);
  nand (_15180_, _14795_, _14777_);
  nand (_15181_, _14779_, _23742_);
  nand (_23743_, _15181_, _15180_);
  nand (_15182_, _14799_, _14777_);
  nand (_15183_, _14779_, _23744_);
  nand (_23745_, _15183_, _15182_);
  nand (_15184_, _14802_, _14777_);
  nand (_15185_, _14779_, _23746_);
  nand (_23747_, _15185_, _15184_);
  nand (_15186_, _14805_, _14777_);
  nand (_15187_, _14779_, _23748_);
  nand (_23749_, _15187_, _15186_);
  nand (_15189_, _14808_, _14777_);
  nand (_15190_, _14779_, _23750_);
  nand (_23751_, _15190_, _15189_);
  nand (_15191_, _14773_, _14789_);
  nand (_15192_, _14775_, _23752_);
  nand (_23753_, _15192_, _15191_);
  nand (_15193_, _14792_, _14773_);
  nand (_15194_, _14775_, _23754_);
  nand (_23755_, _15194_, _15193_);
  nand (_15195_, _14795_, _14773_);
  nand (_15196_, _14775_, _23756_);
  nand (_23757_, _15196_, _15195_);
  nand (_15197_, _14799_, _14773_);
  nand (_15198_, _14775_, _23758_);
  nand (_23759_, _15198_, _15197_);
  nand (_15199_, _14802_, _14773_);
  nand (_15200_, _14775_, _23760_);
  nand (_23761_, _15200_, _15199_);
  nand (_15201_, _14805_, _14773_);
  nand (_15202_, _14775_, _23762_);
  nand (_23763_, _15202_, _15201_);
  nand (_15203_, _14808_, _14773_);
  nand (_15204_, _14775_, _23764_);
  nand (_23765_, _15204_, _15203_);
  nand (_15205_, _14769_, _14789_);
  nand (_15206_, _14771_, _23766_);
  nand (_23767_, _15206_, _15205_);
  nand (_15207_, _14792_, _14769_);
  nand (_15208_, _14771_, _23768_);
  nand (_23769_, _15208_, _15207_);
  nand (_15209_, _14795_, _14769_);
  nand (_15210_, _14771_, _23770_);
  nand (_23771_, _15210_, _15209_);
  nand (_15211_, _14799_, _14769_);
  nand (_15212_, _14771_, _23772_);
  nand (_23773_, _15212_, _15211_);
  nand (_15213_, _14802_, _14769_);
  nand (_15214_, _14771_, _23774_);
  nand (_23775_, _15214_, _15213_);
  nand (_15215_, _14805_, _14769_);
  nand (_15217_, _14771_, _23776_);
  nand (_23777_, _15217_, _15215_);
  nand (_15218_, _14808_, _14769_);
  nand (_15219_, _14771_, _23778_);
  nand (_23779_, _15219_, _15218_);
  nand (_15220_, _14764_, _14789_);
  nand (_15221_, _14767_, _23780_);
  nand (_23781_, _15221_, _15220_);
  nand (_15222_, _14792_, _14764_);
  nand (_15223_, _14767_, _23783_);
  nand (_23784_, _15223_, _15222_);
  nand (_15224_, _14795_, _14764_);
  nand (_15225_, _14767_, _23785_);
  nand (_23786_, _15225_, _15224_);
  nand (_15226_, _14799_, _14764_);
  nand (_15227_, _14767_, _23787_);
  nand (_23788_, _15227_, _15226_);
  nand (_15228_, _14802_, _14764_);
  nand (_15229_, _14767_, _23789_);
  nand (_23790_, _15229_, _15228_);
  nand (_15230_, _14805_, _14764_);
  nand (_15231_, _14767_, _23791_);
  nand (_23792_, _15231_, _15230_);
  nand (_15232_, _14808_, _14764_);
  nand (_15233_, _14767_, _23793_);
  nand (_23794_, _15233_, _15232_);
  nand (_15234_, _14760_, _14789_);
  nand (_15235_, _14762_, _23795_);
  nand (_23796_, _15235_, _15234_);
  nand (_15236_, _14792_, _14760_);
  nand (_15237_, _14762_, _23797_);
  nand (_23798_, _15237_, _15236_);
  nand (_15238_, _14795_, _14760_);
  nand (_15239_, _14762_, _23799_);
  nand (_23800_, _15239_, _15238_);
  nand (_15240_, _14799_, _14760_);
  nand (_15241_, _14762_, _23801_);
  nand (_23802_, _15241_, _15240_);
  nand (_15242_, _14802_, _14760_);
  nand (_15243_, _14762_, _23803_);
  nand (_23804_, _15243_, _15242_);
  nand (_15245_, _14805_, _14760_);
  nand (_15246_, _14762_, _23805_);
  nand (_23806_, _15246_, _15245_);
  nand (_15247_, _14808_, _14760_);
  nand (_15248_, _14762_, _23807_);
  nand (_23808_, _15248_, _15247_);
  nand (_15249_, _14756_, _14789_);
  nand (_15250_, _14758_, _23809_);
  nand (_23810_, _15250_, _15249_);
  nand (_15251_, _14792_, _14756_);
  nand (_15252_, _14758_, _23811_);
  nand (_23812_, _15252_, _15251_);
  nand (_15253_, _14795_, _14756_);
  nand (_15254_, _14758_, _23813_);
  nand (_23814_, _15254_, _15253_);
  nand (_15255_, _14799_, _14756_);
  nand (_15256_, _14758_, _23815_);
  nand (_23816_, _15256_, _15255_);
  nand (_15257_, _14802_, _14756_);
  nand (_15258_, _14758_, _23817_);
  nand (_23818_, _15258_, _15257_);
  nand (_15259_, _14805_, _14756_);
  nand (_15260_, _14758_, _23819_);
  nand (_23820_, _15260_, _15259_);
  nand (_15261_, _14808_, _14756_);
  nand (_15262_, _14758_, _23821_);
  nand (_23822_, _15262_, _15261_);
  nand (_15263_, _14752_, _14789_);
  nand (_15264_, _14754_, _23824_);
  nand (_23825_, _15264_, _15263_);
  nand (_15265_, _14792_, _14752_);
  nand (_15266_, _14754_, _23826_);
  nand (_23827_, _15266_, _15265_);
  nand (_15267_, _14795_, _14752_);
  nand (_15268_, _14754_, _23828_);
  nand (_23829_, _15268_, _15267_);
  nand (_15269_, _14799_, _14752_);
  nand (_15270_, _14754_, _23830_);
  nand (_23831_, _15270_, _15269_);
  nand (_15272_, _14802_, _14752_);
  nand (_15273_, _14754_, _23832_);
  nand (_23833_, _15273_, _15272_);
  nand (_15274_, _14805_, _14752_);
  nand (_15275_, _14754_, _23834_);
  nand (_23835_, _15275_, _15274_);
  nand (_15276_, _14808_, _14752_);
  nand (_15277_, _14754_, _23836_);
  nand (_23837_, _15277_, _15276_);
  nand (_15278_, _14748_, _14789_);
  nand (_15279_, _14750_, _23838_);
  nand (_23839_, _15279_, _15278_);
  nand (_15280_, _14792_, _14748_);
  nand (_15281_, _14750_, _23840_);
  nand (_23841_, _15281_, _15280_);
  nand (_15282_, _14795_, _14748_);
  nand (_15283_, _14750_, _23842_);
  nand (_23843_, _15283_, _15282_);
  nand (_15284_, _14799_, _14748_);
  nand (_15285_, _14750_, _23844_);
  nand (_23845_, _15285_, _15284_);
  nand (_15286_, _14802_, _14748_);
  nand (_15287_, _14750_, _23846_);
  nand (_23847_, _15287_, _15286_);
  nand (_15288_, _14805_, _14748_);
  nand (_15289_, _14750_, _23848_);
  nand (_23849_, _15289_, _15288_);
  nand (_15290_, _14808_, _14748_);
  nand (_15291_, _14750_, _23850_);
  nand (_23851_, _15291_, _15290_);
  nand (_15292_, _14744_, _14789_);
  nand (_15293_, _14746_, _23852_);
  nand (_23853_, _15293_, _15292_);
  nand (_15294_, _14792_, _14744_);
  nand (_15295_, _14746_, _23854_);
  nand (_23855_, _15295_, _15294_);
  nand (_15296_, _14795_, _14744_);
  nand (_15297_, _14746_, _23856_);
  nand (_23857_, _15297_, _15296_);
  nand (_15298_, _14799_, _14744_);
  nand (_15299_, _14746_, _23858_);
  nand (_23859_, _15299_, _15298_);
  nand (_15300_, _14802_, _14744_);
  nand (_15301_, _14746_, _23860_);
  nand (_23861_, _15301_, _15300_);
  nand (_15302_, _14805_, _14744_);
  nand (_15303_, _14746_, _23862_);
  nand (_23863_, _15303_, _15302_);
  nand (_15304_, _14808_, _14744_);
  nand (_15305_, _14746_, _23865_);
  nand (_23866_, _15305_, _15304_);
  nand (_15306_, _14740_, _14789_);
  nand (_15307_, _14742_, _23867_);
  nand (_23868_, _15307_, _15306_);
  nand (_15308_, _14792_, _14740_);
  nand (_15309_, _14742_, _23869_);
  nand (_23870_, _15309_, _15308_);
  nand (_15310_, _14795_, _14740_);
  nand (_15311_, _14742_, _23871_);
  nand (_23872_, _15311_, _15310_);
  nand (_15312_, _14799_, _14740_);
  nand (_15313_, _14742_, _23873_);
  nand (_23874_, _15313_, _15312_);
  nand (_15314_, _14802_, _14740_);
  nand (_15315_, _14742_, _23875_);
  nand (_23876_, _15315_, _15314_);
  nand (_15316_, _14805_, _14740_);
  nand (_15317_, _14742_, _23877_);
  nand (_23878_, _15317_, _15316_);
  nand (_15318_, _14808_, _14740_);
  nand (_15319_, _14742_, _23879_);
  nand (_23880_, _15319_, _15318_);
  nand (_15320_, _14736_, _14789_);
  nand (_15321_, _14738_, _23881_);
  nand (_23882_, _15321_, _15320_);
  nand (_15322_, _14792_, _14736_);
  nand (_15323_, _14738_, _23883_);
  nand (_23884_, _15323_, _15322_);
  nand (_15324_, _14795_, _14736_);
  nand (_15325_, _14738_, _23885_);
  nand (_23886_, _15325_, _15324_);
  nand (_15326_, _14799_, _14736_);
  nand (_15327_, _14738_, _23887_);
  nand (_23888_, _15327_, _15326_);
  nand (_15328_, _14802_, _14736_);
  nand (_15329_, _14738_, _23889_);
  nand (_23890_, _15329_, _15328_);
  nand (_15330_, _14805_, _14736_);
  nand (_15331_, _14738_, _23891_);
  nand (_23892_, _15331_, _15330_);
  nand (_15332_, _14808_, _14736_);
  nand (_15333_, _14738_, _23893_);
  nand (_23894_, _15333_, _15332_);
  nand (_15334_, _14731_, _14789_);
  nand (_15335_, _14734_, _23895_);
  nand (_23896_, _15335_, _15334_);
  nand (_15336_, _14792_, _14731_);
  nand (_15337_, _14734_, _23897_);
  nand (_23898_, _15337_, _15336_);
  nand (_15338_, _14795_, _14731_);
  nand (_15339_, _14734_, _23899_);
  nand (_23900_, _15339_, _15338_);
  nand (_15340_, _14799_, _14731_);
  nand (_15341_, _14734_, _23901_);
  nand (_23902_, _15341_, _15340_);
  nand (_15342_, _14802_, _14731_);
  nand (_15343_, _14734_, _23903_);
  nand (_23904_, _15343_, _15342_);
  nand (_15344_, _14805_, _14731_);
  nand (_15345_, _14734_, _23906_);
  nand (_23907_, _15345_, _15344_);
  nand (_15346_, _14808_, _14731_);
  nand (_15347_, _14734_, _23908_);
  nand (_23909_, _15347_, _15346_);
  nand (_15348_, _14727_, _14789_);
  nand (_15349_, _14729_, _23910_);
  nand (_23911_, _15349_, _15348_);
  nand (_15350_, _14792_, _14727_);
  nand (_15351_, _14729_, _23912_);
  nand (_23913_, _15351_, _15350_);
  nand (_15352_, _14795_, _14727_);
  nand (_15353_, _14729_, _23914_);
  nand (_23915_, _15353_, _15352_);
  nand (_15354_, _14799_, _14727_);
  nand (_15355_, _14729_, _23916_);
  nand (_23917_, _15355_, _15354_);
  nand (_15356_, _14802_, _14727_);
  nand (_15357_, _14729_, _23918_);
  nand (_23919_, _15357_, _15356_);
  nand (_15358_, _14805_, _14727_);
  nand (_15359_, _14729_, _23920_);
  nand (_23921_, _15359_, _15358_);
  nand (_15360_, _14808_, _14727_);
  nand (_15361_, _14729_, _23922_);
  nand (_23923_, _15361_, _15360_);
  nand (_15362_, _14723_, _14789_);
  nand (_15363_, _14725_, _23924_);
  nand (_23925_, _15363_, _15362_);
  nand (_15364_, _14792_, _14723_);
  nand (_15365_, _14725_, _23926_);
  nand (_23927_, _15365_, _15364_);
  nand (_15366_, _14795_, _14723_);
  nand (_15367_, _14725_, _23928_);
  nand (_23929_, _15367_, _15366_);
  nand (_15368_, _14799_, _14723_);
  nand (_15369_, _14725_, _23930_);
  nand (_23931_, _15369_, _15368_);
  nand (_15370_, _14802_, _14723_);
  nand (_15371_, _14725_, _23932_);
  nand (_23933_, _15371_, _15370_);
  nand (_15372_, _14805_, _14723_);
  nand (_15373_, _14725_, _23934_);
  nand (_23935_, _15373_, _15372_);
  nand (_15374_, _14808_, _14723_);
  nand (_15375_, _14725_, _23936_);
  nand (_23937_, _15375_, _15374_);
  nand (_15376_, _14718_, _23938_);
  nand (_15377_, _14717_, _14789_);
  nand (_23939_, _15377_, _15376_);
  nand (_15378_, _14718_, _23940_);
  nand (_15379_, _14792_, _14717_);
  nand (_23941_, _15379_, _15378_);
  nand (_15380_, _14718_, _23942_);
  nand (_15381_, _14795_, _14717_);
  nand (_23943_, _15381_, _15380_);
  nand (_15382_, _14718_, _23944_);
  nand (_15383_, _14799_, _14717_);
  nand (_23945_, _15383_, _15382_);
  nand (_15384_, _14718_, _23947_);
  nand (_15385_, _14802_, _14717_);
  nand (_23948_, _15385_, _15384_);
  nand (_15386_, _14718_, _23949_);
  nand (_15387_, _14805_, _14717_);
  nand (_23950_, _15387_, _15386_);
  nand (_15388_, _14718_, _23951_);
  nand (_15389_, _14808_, _14717_);
  nand (_23952_, _15389_, _15388_);
  nand (_15390_, _14714_, _23953_);
  nand (_15391_, _14713_, _14789_);
  nand (_23954_, _15391_, _15390_);
  nand (_15392_, _14714_, _23955_);
  nand (_15393_, _14792_, _14713_);
  nand (_23956_, _15393_, _15392_);
  nand (_15394_, _14714_, _23957_);
  nand (_15395_, _14795_, _14713_);
  nand (_23958_, _15395_, _15394_);
  nand (_15396_, _14714_, _23959_);
  nand (_15397_, _14799_, _14713_);
  nand (_23960_, _15397_, _15396_);
  nand (_15398_, _14714_, _23961_);
  nand (_15399_, _14802_, _14713_);
  nand (_23962_, _15399_, _15398_);
  nand (_15400_, _14714_, _23963_);
  nand (_15401_, _14805_, _14713_);
  nand (_23964_, _15401_, _15400_);
  nand (_15402_, _14714_, _23965_);
  nand (_15403_, _14808_, _14713_);
  nand (_23966_, _15403_, _15402_);
  nand (_15404_, _14710_, _23967_);
  nand (_15405_, _14709_, _14789_);
  nand (_23968_, _15405_, _15404_);
  nand (_15406_, _14710_, _23969_);
  nand (_15407_, _14792_, _14709_);
  nand (_23970_, _15407_, _15406_);
  nand (_15408_, _14710_, _23971_);
  nand (_15409_, _14795_, _14709_);
  nand (_23972_, _15409_, _15408_);
  nand (_15410_, _14710_, _23973_);
  nand (_15411_, _14799_, _14709_);
  nand (_23974_, _15411_, _15410_);
  nand (_15413_, _14710_, _23975_);
  nand (_15414_, _14802_, _14709_);
  nand (_23976_, _15414_, _15413_);
  nand (_15415_, _14710_, _23977_);
  nand (_15416_, _14805_, _14709_);
  nand (_23978_, _15416_, _15415_);
  nand (_15417_, _14710_, _23979_);
  nand (_15418_, _14808_, _14709_);
  nand (_23980_, _15418_, _15417_);
  nand (_15419_, _14706_, _23981_);
  nand (_15420_, _14705_, _14789_);
  nand (_23982_, _15420_, _15419_);
  nand (_15421_, _14706_, _23983_);
  nand (_15422_, _14792_, _14705_);
  nand (_23984_, _15422_, _15421_);
  nand (_15423_, _14706_, _23985_);
  nand (_15424_, _14795_, _14705_);
  nand (_23986_, _15424_, _15423_);
  nand (_15425_, _14706_, _23988_);
  nand (_15426_, _14799_, _14705_);
  nand (_23989_, _15426_, _15425_);
  nand (_15427_, _14706_, _23990_);
  nand (_15428_, _14802_, _14705_);
  nand (_23991_, _15428_, _15427_);
  nand (_15429_, _14706_, _23992_);
  nand (_15430_, _14805_, _14705_);
  nand (_23993_, _15430_, _15429_);
  nand (_15431_, _14706_, _23994_);
  nand (_15432_, _14808_, _14705_);
  nand (_23995_, _15432_, _15431_);
  nand (_15433_, _14702_, _23996_);
  nand (_15434_, _14701_, _14789_);
  nand (_23997_, _15434_, _15433_);
  nand (_15435_, _14702_, _23998_);
  nand (_15436_, _14792_, _14701_);
  nand (_23999_, _15436_, _15435_);
  nand (_15437_, _14702_, _24000_);
  nand (_15438_, _14795_, _14701_);
  nand (_24001_, _15438_, _15437_);
  nand (_15439_, _14702_, _24002_);
  nand (_15440_, _14799_, _14701_);
  nand (_24003_, _15440_, _15439_);
  nand (_15441_, _14702_, _24004_);
  nand (_15442_, _14802_, _14701_);
  nand (_24005_, _15442_, _15441_);
  nand (_15443_, _14702_, _24006_);
  nand (_15444_, _14805_, _14701_);
  nand (_24007_, _15444_, _15443_);
  nand (_15445_, _14702_, _24008_);
  nand (_15446_, _14808_, _14701_);
  nand (_24009_, _15446_, _15445_);
  nand (_15447_, _14697_, _24010_);
  nand (_15448_, _14696_, _14789_);
  nand (_24011_, _15448_, _15447_);
  nand (_15449_, _14697_, _24012_);
  nand (_15450_, _14792_, _14696_);
  nand (_24013_, _15450_, _15449_);
  nand (_15451_, _14697_, _24014_);
  nand (_15452_, _14795_, _14696_);
  nand (_24015_, _15452_, _15451_);
  nand (_15453_, _14697_, _24016_);
  nand (_15454_, _14799_, _14696_);
  nand (_24017_, _15454_, _15453_);
  nand (_15455_, _14697_, _24018_);
  nand (_15456_, _14802_, _14696_);
  nand (_24019_, _15456_, _15455_);
  nand (_15457_, _14697_, _24020_);
  nand (_15458_, _14805_, _14696_);
  nand (_24021_, _15458_, _15457_);
  nand (_15459_, _14697_, _24022_);
  nand (_15460_, _14808_, _14696_);
  nand (_24023_, _15460_, _15459_);
  nand (_15461_, _14693_, _24024_);
  nand (_15462_, _14692_, _14789_);
  nand (_24025_, _15462_, _15461_);
  nand (_15463_, _14693_, _24026_);
  nand (_15464_, _14792_, _14692_);
  nand (_24027_, _15464_, _15463_);
  nand (_15465_, _14693_, _24029_);
  nand (_15466_, _14795_, _14692_);
  nand (_24030_, _15466_, _15465_);
  nand (_15467_, _14693_, _24031_);
  nand (_15468_, _14799_, _14692_);
  nand (_24032_, _15468_, _15467_);
  nand (_15469_, _14693_, _24033_);
  nand (_15470_, _14802_, _14692_);
  nand (_24034_, _15470_, _15469_);
  nand (_15471_, _14693_, _24035_);
  nand (_15472_, _14805_, _14692_);
  nand (_24036_, _15472_, _15471_);
  nand (_15474_, _14693_, _24037_);
  nand (_15475_, _14808_, _14692_);
  nand (_24038_, _15475_, _15474_);
  nand (_15476_, _14689_, _24039_);
  nand (_15477_, _14688_, _14789_);
  nand (_24040_, _15477_, _15476_);
  nand (_15478_, _14689_, _24041_);
  nand (_15479_, _14792_, _14688_);
  nand (_24042_, _15479_, _15478_);
  nand (_15480_, _14689_, _24043_);
  nand (_15481_, _14795_, _14688_);
  nand (_24044_, _15481_, _15480_);
  nand (_15482_, _14689_, _24045_);
  nand (_15483_, _14799_, _14688_);
  nand (_24046_, _15483_, _15482_);
  nand (_15484_, _14689_, _24047_);
  nand (_15485_, _14802_, _14688_);
  nand (_24048_, _15485_, _15484_);
  nand (_15486_, _14689_, _24049_);
  nand (_15487_, _14805_, _14688_);
  nand (_24050_, _15487_, _15486_);
  nand (_15489_, _14689_, _24051_);
  nand (_15490_, _14808_, _14688_);
  nand (_24052_, _15490_, _15489_);
  nand (_15491_, _14685_, _24053_);
  nand (_15492_, _14684_, _14789_);
  nand (_24054_, _15492_, _15491_);
  nand (_15493_, _14685_, _24055_);
  nand (_15494_, _14792_, _14684_);
  nand (_24056_, _15494_, _15493_);
  nand (_15495_, _14685_, _24057_);
  nand (_15496_, _14795_, _14684_);
  nand (_24058_, _15496_, _15495_);
  nand (_15497_, _14685_, _24059_);
  nand (_15498_, _14799_, _14684_);
  nand (_24060_, _15498_, _15497_);
  nand (_15499_, _14685_, _24061_);
  nand (_15500_, _14802_, _14684_);
  nand (_24062_, _15500_, _15499_);
  nand (_15501_, _14685_, _24063_);
  nand (_15502_, _14805_, _14684_);
  nand (_24064_, _15502_, _15501_);
  nand (_15503_, _14685_, _24065_);
  nand (_15504_, _14808_, _14684_);
  nand (_24066_, _15504_, _15503_);
  nand (_15505_, _14681_, _24067_);
  nand (_15506_, _14680_, _14789_);
  nand (_24068_, _15506_, _15505_);
  nand (_15507_, _14681_, _24070_);
  nand (_15508_, _14792_, _14680_);
  nand (_24071_, _15508_, _15507_);
  nand (_15509_, _14681_, _24072_);
  nand (_15510_, _14795_, _14680_);
  nand (_24073_, _15510_, _15509_);
  nand (_15511_, _14681_, _24074_);
  nand (_15512_, _14799_, _14680_);
  nand (_24075_, _15512_, _15511_);
  nand (_15513_, _14681_, _24076_);
  nand (_15514_, _14802_, _14680_);
  nand (_24077_, _15514_, _15513_);
  nand (_15515_, _14681_, _24078_);
  nand (_15516_, _14805_, _14680_);
  nand (_24079_, _15516_, _15515_);
  nand (_15517_, _14681_, _24080_);
  nand (_15518_, _14808_, _14680_);
  nand (_24081_, _15518_, _15517_);
  nand (_15519_, _14677_, _24082_);
  nand (_15520_, _14676_, _14789_);
  nand (_24083_, _15520_, _15519_);
  nand (_15521_, _14677_, _24084_);
  nand (_15522_, _14792_, _14676_);
  nand (_24085_, _15522_, _15521_);
  nand (_15523_, _14677_, _24086_);
  nand (_15524_, _14795_, _14676_);
  nand (_24087_, _15524_, _15523_);
  nand (_15525_, _14677_, _24088_);
  nand (_15526_, _14799_, _14676_);
  nand (_24089_, _15526_, _15525_);
  nand (_15527_, _14677_, _24090_);
  nand (_15528_, _14802_, _14676_);
  nand (_24091_, _15528_, _15527_);
  nand (_15529_, _14677_, _24092_);
  nand (_15530_, _14805_, _14676_);
  nand (_24093_, _15530_, _15529_);
  nand (_15531_, _14677_, _24094_);
  nand (_15532_, _14808_, _14676_);
  nand (_24095_, _15532_, _15531_);
  nand (_15533_, _14673_, _24096_);
  nand (_15534_, _14672_, _14789_);
  nand (_24097_, _15534_, _15533_);
  nand (_15536_, _14673_, _24098_);
  nand (_15537_, _14792_, _14672_);
  nand (_24099_, _15537_, _15536_);
  nand (_15538_, _14673_, _24100_);
  nand (_15539_, _14795_, _14672_);
  nand (_24101_, _15539_, _15538_);
  nand (_15540_, _14673_, _24102_);
  nand (_15541_, _14799_, _14672_);
  nand (_24103_, _15541_, _15540_);
  nand (_15542_, _14673_, _24104_);
  nand (_15544_, _14802_, _14672_);
  nand (_24105_, _15544_, _15542_);
  nand (_15545_, _14673_, _24106_);
  nand (_15546_, _14805_, _14672_);
  nand (_24107_, _15546_, _15545_);
  nand (_15547_, _14673_, _24108_);
  nand (_15548_, _14808_, _14672_);
  nand (_24109_, _15548_, _15547_);
  nand (_15549_, _14669_, _24112_);
  nand (_15550_, _14668_, _14789_);
  nand (_24113_, _15550_, _15549_);
  nand (_15551_, _14669_, _24114_);
  nand (_15552_, _14792_, _14668_);
  nand (_24115_, _15552_, _15551_);
  nand (_15553_, _14669_, _24116_);
  nand (_15554_, _14795_, _14668_);
  nand (_24117_, _15554_, _15553_);
  nand (_15555_, _14669_, _24118_);
  nand (_15556_, _14799_, _14668_);
  nand (_24119_, _15556_, _15555_);
  nand (_15557_, _14669_, _24120_);
  nand (_15558_, _14802_, _14668_);
  nand (_24121_, _15558_, _15557_);
  nand (_15559_, _14669_, _24122_);
  nand (_15560_, _14805_, _14668_);
  nand (_24123_, _15560_, _15559_);
  nand (_15561_, _14669_, _24124_);
  nand (_15562_, _14808_, _14668_);
  nand (_24125_, _15562_, _15561_);
  nand (_15563_, _14664_, _24126_);
  nand (_15564_, _14663_, _14789_);
  nand (_24127_, _15564_, _15563_);
  nand (_15565_, _14664_, _24128_);
  nand (_15566_, _14792_, _14663_);
  nand (_24129_, _15566_, _15565_);
  nand (_15567_, _14664_, _24130_);
  nand (_15568_, _14795_, _14663_);
  nand (_24131_, _15568_, _15567_);
  nand (_15569_, _14664_, _24132_);
  nand (_15570_, _14799_, _14663_);
  nand (_24133_, _15570_, _15569_);
  nand (_15571_, _14664_, _24134_);
  nand (_15572_, _14802_, _14663_);
  nand (_24135_, _15572_, _15571_);
  nand (_15573_, _14664_, _24136_);
  nand (_15574_, _14805_, _14663_);
  nand (_24137_, _15574_, _15573_);
  nand (_15575_, _14664_, _24138_);
  nand (_15576_, _14808_, _14663_);
  nand (_24139_, _15576_, _15575_);
  nand (_15577_, _14660_, _24140_);
  nand (_15578_, _14659_, _14789_);
  nand (_24141_, _15578_, _15577_);
  nand (_15579_, _14660_, _24142_);
  nand (_15580_, _14792_, _14659_);
  nand (_24143_, _15580_, _15579_);
  nand (_15581_, _14660_, _24144_);
  nand (_15582_, _14795_, _14659_);
  nand (_24145_, _15582_, _15581_);
  nand (_15583_, _14660_, _24146_);
  nand (_15584_, _14799_, _14659_);
  nand (_24147_, _15584_, _15583_);
  nand (_15585_, _14660_, _24148_);
  nand (_15586_, _14802_, _14659_);
  nand (_24149_, _15586_, _15585_);
  nand (_15587_, _14660_, _24150_);
  nand (_15588_, _14805_, _14659_);
  nand (_24151_, _15588_, _15587_);
  nand (_15589_, _14660_, _24153_);
  nand (_15590_, _14808_, _14659_);
  nand (_24154_, _15590_, _15589_);
  nand (_15592_, _14656_, _24155_);
  nand (_15593_, _14655_, _14789_);
  nand (_24156_, _15593_, _15592_);
  nand (_15594_, _14656_, _24157_);
  nand (_15595_, _14792_, _14655_);
  nand (_24158_, _15595_, _15594_);
  nand (_15596_, _14656_, _24159_);
  nand (_15597_, _14795_, _14655_);
  nand (_24160_, _15597_, _15596_);
  nand (_15599_, _14656_, _24161_);
  nand (_15600_, _14799_, _14655_);
  nand (_24162_, _15600_, _15599_);
  nand (_15601_, _14656_, _24163_);
  nand (_15602_, _14802_, _14655_);
  nand (_24164_, _15602_, _15601_);
  nand (_15603_, _14656_, _24165_);
  nand (_15604_, _14805_, _14655_);
  nand (_24166_, _15604_, _15603_);
  nand (_15605_, _14656_, _24167_);
  nand (_15606_, _14808_, _14655_);
  nand (_24168_, _15606_, _15605_);
  nand (_15607_, _14649_, _14789_);
  nand (_15608_, _14651_, _24169_);
  nand (_24170_, _15608_, _15607_);
  nand (_15609_, _14792_, _14649_);
  nand (_15610_, _14651_, _24171_);
  nand (_24172_, _15610_, _15609_);
  nand (_15611_, _14795_, _14649_);
  nand (_15612_, _14651_, _24173_);
  nand (_24174_, _15612_, _15611_);
  nand (_15613_, _14799_, _14649_);
  nand (_15614_, _14651_, _24175_);
  nand (_24176_, _15614_, _15613_);
  nand (_15615_, _14802_, _14649_);
  nand (_15616_, _14651_, _24177_);
  nand (_24178_, _15616_, _15615_);
  nand (_15617_, _14805_, _14649_);
  nand (_15618_, _14651_, _24179_);
  nand (_24180_, _15618_, _15617_);
  nand (_15619_, _14808_, _14649_);
  nand (_15620_, _14651_, _24181_);
  nand (_24182_, _15620_, _15619_);
  nand (_15621_, _14645_, _14789_);
  nand (_15622_, _14647_, _24183_);
  nand (_24184_, _15622_, _15621_);
  nand (_15623_, _14792_, _14645_);
  nand (_15624_, _14647_, _24185_);
  nand (_24186_, _15624_, _15623_);
  nand (_15625_, _14795_, _14645_);
  nand (_15626_, _14647_, _24187_);
  nand (_24188_, _15626_, _15625_);
  nand (_15627_, _14799_, _14645_);
  nand (_15628_, _14647_, _24189_);
  nand (_24190_, _15628_, _15627_);
  nand (_15629_, _14802_, _14645_);
  nand (_15630_, _14647_, _24191_);
  nand (_24192_, _15630_, _15629_);
  nand (_15631_, _14805_, _14645_);
  nand (_15632_, _14647_, _24194_);
  nand (_24195_, _15632_, _15631_);
  nand (_15634_, _14808_, _14645_);
  nand (_15635_, _14647_, _24196_);
  nand (_24197_, _15635_, _15634_);
  nand (_15636_, _14641_, _14789_);
  nand (_15637_, _14643_, _24198_);
  nand (_24199_, _15637_, _15636_);
  nand (_15638_, _14792_, _14641_);
  nand (_15639_, _14643_, _24200_);
  nand (_24201_, _15639_, _15638_);
  nand (_15641_, _14795_, _14641_);
  nand (_15642_, _14643_, _24202_);
  nand (_24203_, _15642_, _15641_);
  nand (_15643_, _14799_, _14641_);
  nand (_15644_, _14643_, _24204_);
  nand (_24205_, _15644_, _15643_);
  nand (_15645_, _14802_, _14641_);
  nand (_15646_, _14643_, _24206_);
  nand (_24207_, _15646_, _15645_);
  nand (_15647_, _14805_, _14641_);
  nand (_15648_, _14643_, _24208_);
  nand (_24209_, _15648_, _15647_);
  nand (_15649_, _14808_, _14641_);
  nand (_15650_, _14643_, _24210_);
  nand (_24211_, _15650_, _15649_);
  nand (_15651_, _14637_, _14789_);
  nand (_15652_, _14639_, _24212_);
  nand (_24213_, _15652_, _15651_);
  nand (_15653_, _14792_, _14637_);
  nand (_15654_, _14639_, _24214_);
  nand (_24215_, _15654_, _15653_);
  nand (_15655_, _14795_, _14637_);
  nand (_15656_, _14639_, _24216_);
  nand (_24217_, _15656_, _15655_);
  nand (_15657_, _14799_, _14637_);
  nand (_15658_, _14639_, _24218_);
  nand (_24219_, _15658_, _15657_);
  nand (_15659_, _14802_, _14637_);
  nand (_15660_, _14639_, _24220_);
  nand (_24221_, _15660_, _15659_);
  nand (_15661_, _14805_, _14637_);
  nand (_15662_, _14639_, _24222_);
  nand (_24223_, _15662_, _15661_);
  nand (_15663_, _14808_, _14637_);
  nand (_15664_, _14639_, _24224_);
  nand (_24225_, _15664_, _15663_);
  nand (_15665_, _14633_, _14789_);
  nand (_15666_, _14635_, _24226_);
  nand (_24227_, _15666_, _15665_);
  nand (_15667_, _14792_, _14633_);
  nand (_15668_, _14635_, _24228_);
  nand (_24229_, _15668_, _15667_);
  nand (_15669_, _14795_, _14633_);
  nand (_15670_, _14635_, _24230_);
  nand (_24231_, _15670_, _15669_);
  nand (_15671_, _14799_, _14633_);
  nand (_15672_, _14635_, _24232_);
  nand (_24233_, _15672_, _15671_);
  nand (_15673_, _14802_, _14633_);
  nand (_15674_, _14635_, _24235_);
  nand (_24236_, _15674_, _15673_);
  nand (_15675_, _14805_, _14633_);
  nand (_15676_, _14635_, _24237_);
  nand (_24238_, _15676_, _15675_);
  nand (_15677_, _14808_, _14633_);
  nand (_15678_, _14635_, _24239_);
  nand (_24240_, _15678_, _15677_);
  nand (_15679_, _14628_, _14789_);
  nand (_15680_, _14630_, _24241_);
  nand (_24242_, _15680_, _15679_);
  nand (_15681_, _14792_, _14628_);
  nand (_15682_, _14630_, _24243_);
  nand (_24244_, _15682_, _15681_);
  nand (_15683_, _14795_, _14628_);
  nand (_15684_, _14630_, _24245_);
  nand (_24246_, _15684_, _15683_);
  nand (_15685_, _14799_, _14628_);
  nand (_15686_, _14630_, _24247_);
  nand (_24248_, _15686_, _15685_);
  nand (_15687_, _14802_, _14628_);
  nand (_15690_, _14630_, _24249_);
  nand (_24250_, _15690_, _15687_);
  nand (_15691_, _14805_, _14628_);
  nand (_15692_, _14630_, _24251_);
  nand (_24252_, _15692_, _15691_);
  nand (_15693_, _14808_, _14628_);
  nand (_15694_, _14630_, _24253_);
  nand (_24254_, _15694_, _15693_);
  nand (_15695_, _14624_, _14789_);
  nand (_15696_, _14626_, _24255_);
  nand (_24256_, _15696_, _15695_);
  nand (_15698_, _14792_, _14624_);
  nand (_15699_, _14626_, _24257_);
  nand (_24258_, _15699_, _15698_);
  nand (_15700_, _14795_, _14624_);
  nand (_15701_, _14626_, _24259_);
  nand (_24260_, _15701_, _15700_);
  nand (_15702_, _14799_, _14624_);
  nand (_15703_, _14626_, _24261_);
  nand (_24262_, _15703_, _15702_);
  nand (_15704_, _14802_, _14624_);
  nand (_15705_, _14626_, _24263_);
  nand (_24264_, _15705_, _15704_);
  nand (_15706_, _14805_, _14624_);
  nand (_15707_, _14626_, _24265_);
  nand (_24266_, _15707_, _15706_);
  nand (_15708_, _14808_, _14624_);
  nand (_15709_, _14626_, _24267_);
  nand (_24268_, _15709_, _15708_);
  nand (_15710_, _14620_, _14789_);
  nand (_15711_, _14622_, _24269_);
  nand (_24270_, _15711_, _15710_);
  nand (_15712_, _14792_, _14620_);
  nand (_15713_, _14622_, _24271_);
  nand (_24272_, _15713_, _15712_);
  nand (_15714_, _14795_, _14620_);
  nand (_15715_, _14622_, _24273_);
  nand (_24274_, _15715_, _15714_);
  nand (_15716_, _14799_, _14620_);
  nand (_15717_, _14622_, _24276_);
  nand (_24277_, _15717_, _15716_);
  nand (_15718_, _14802_, _14620_);
  nand (_15719_, _14622_, _24278_);
  nand (_24279_, _15719_, _15718_);
  nand (_15720_, _14805_, _14620_);
  nand (_15721_, _14622_, _24280_);
  nand (_24281_, _15721_, _15720_);
  nand (_15722_, _14808_, _14620_);
  nand (_15723_, _14622_, _24282_);
  nand (_24283_, _15723_, _15722_);
  nand (_15725_, _14616_, _14789_);
  nand (_15726_, _14618_, _24284_);
  nand (_24285_, _15726_, _15725_);
  nand (_15727_, _14792_, _14616_);
  nand (_15728_, _14618_, _24286_);
  nand (_24287_, _15728_, _15727_);
  nand (_15729_, _14795_, _14616_);
  nand (_15730_, _14618_, _24288_);
  nand (_24289_, _15730_, _15729_);
  nand (_15731_, _14799_, _14616_);
  nand (_15733_, _14618_, _24290_);
  nand (_24291_, _15733_, _15731_);
  nand (_15734_, _14802_, _14616_);
  nand (_15735_, _14618_, _24292_);
  nand (_24293_, _15735_, _15734_);
  nand (_15736_, _14805_, _14616_);
  nand (_15737_, _14618_, _24294_);
  nand (_24295_, _15737_, _15736_);
  nand (_15738_, _14808_, _14616_);
  nand (_15739_, _14618_, _24296_);
  nand (_24297_, _15739_, _15738_);
  nand (_15740_, _14612_, _14789_);
  nand (_15741_, _14614_, _24298_);
  nand (_24299_, _15741_, _15740_);
  nand (_15742_, _14792_, _14612_);
  nand (_15743_, _14614_, _24300_);
  nand (_24301_, _15743_, _15742_);
  nand (_15744_, _14795_, _14612_);
  nand (_15745_, _14614_, _24302_);
  nand (_24303_, _15745_, _15744_);
  nand (_15746_, _14799_, _14612_);
  nand (_15747_, _14614_, _24304_);
  nand (_24305_, _15747_, _15746_);
  nand (_15748_, _14802_, _14612_);
  nand (_15749_, _14614_, _24306_);
  nand (_24307_, _15749_, _15748_);
  nand (_15750_, _14805_, _14612_);
  nand (_15751_, _14614_, _24308_);
  nand (_24309_, _15751_, _15750_);
  nand (_15752_, _14808_, _14612_);
  nand (_15753_, _14614_, _24310_);
  nand (_24311_, _15753_, _15752_);
  nand (_15754_, _14608_, _14789_);
  nand (_15755_, _14610_, _24312_);
  nand (_24313_, _15755_, _15754_);
  nand (_15756_, _14792_, _14608_);
  nand (_15757_, _14610_, _24314_);
  nand (_24315_, _15757_, _15756_);
  nand (_15758_, _14795_, _14608_);
  nand (_15759_, _14610_, _24317_);
  nand (_24318_, _15759_, _15758_);
  nand (_15761_, _14799_, _14608_);
  nand (_15762_, _14610_, _24319_);
  nand (_24320_, _15762_, _15761_);
  nand (_15763_, _14802_, _14608_);
  nand (_15764_, _14610_, _24321_);
  nand (_24322_, _15764_, _15763_);
  nand (_15765_, _14805_, _14608_);
  nand (_15766_, _14610_, _24323_);
  nand (_24324_, _15766_, _15765_);
  nand (_15768_, _14808_, _14608_);
  nand (_15769_, _14610_, _24325_);
  nand (_24326_, _15769_, _15768_);
  nand (_15770_, _14604_, _14789_);
  nand (_15771_, _14606_, _24327_);
  nand (_24328_, _15771_, _15770_);
  nand (_15772_, _14792_, _14604_);
  nand (_15773_, _14606_, _24329_);
  nand (_24330_, _15773_, _15772_);
  nand (_15774_, _14795_, _14604_);
  nand (_15775_, _14606_, _24331_);
  nand (_24332_, _15775_, _15774_);
  nand (_15776_, _14799_, _14604_);
  nand (_15777_, _14606_, _24333_);
  nand (_24334_, _15777_, _15776_);
  nand (_15778_, _14802_, _14604_);
  nand (_15779_, _14606_, _24335_);
  nand (_24336_, _15779_, _15778_);
  nand (_15780_, _14805_, _14604_);
  nand (_15781_, _14606_, _24337_);
  nand (_24338_, _15781_, _15780_);
  nand (_15782_, _14808_, _14604_);
  nand (_15783_, _14606_, _24339_);
  nand (_24340_, _15783_, _15782_);
  nand (_15784_, _14600_, _14789_);
  nand (_15785_, _14602_, _24341_);
  nand (_24342_, _15785_, _15784_);
  nand (_15786_, _14792_, _14600_);
  nand (_15787_, _14602_, _24343_);
  nand (_24344_, _15787_, _15786_);
  nand (_15788_, _14795_, _14600_);
  nand (_15789_, _14602_, _24345_);
  nand (_24346_, _15789_, _15788_);
  nand (_15790_, _14799_, _14600_);
  nand (_15791_, _14602_, _24347_);
  nand (_24348_, _15791_, _15790_);
  nand (_15792_, _14802_, _14600_);
  nand (_15793_, _14602_, _24349_);
  nand (_24350_, _15793_, _15792_);
  nand (_15794_, _14805_, _14600_);
  nand (_15796_, _14602_, _24351_);
  nand (_24352_, _15796_, _15794_);
  nand (_15797_, _14808_, _14600_);
  nand (_15798_, _14602_, _24353_);
  nand (_24354_, _15798_, _15797_);
  nand (_15799_, _14595_, _14789_);
  nand (_15800_, _14597_, _24355_);
  nand (_24356_, _15800_, _15799_);
  nand (_15801_, _14792_, _14595_);
  nand (_15802_, _14597_, _24358_);
  nand (_24359_, _15802_, _15801_);
  nand (_15804_, _14795_, _14595_);
  nand (_15805_, _14597_, _24360_);
  nand (_24361_, _15805_, _15804_);
  nand (_15806_, _14799_, _14595_);
  nand (_15807_, _14597_, _24362_);
  nand (_24363_, _15807_, _15806_);
  nand (_15808_, _14802_, _14595_);
  nand (_15809_, _14597_, _24364_);
  nand (_24365_, _15809_, _15808_);
  nand (_15810_, _14805_, _14595_);
  nand (_15811_, _14597_, _24366_);
  nand (_24367_, _15811_, _15810_);
  nand (_15812_, _14808_, _14595_);
  nand (_15813_, _14597_, _24368_);
  nand (_24369_, _15813_, _15812_);
  nand (_15814_, _14591_, _14789_);
  nand (_15815_, _14593_, _24370_);
  nand (_24371_, _15815_, _15814_);
  nand (_15816_, _14792_, _14591_);
  nand (_15817_, _14593_, _24372_);
  nand (_24373_, _15817_, _15816_);
  nand (_15818_, _14795_, _14591_);
  nand (_15819_, _14593_, _24374_);
  nand (_24375_, _15819_, _15818_);
  nand (_15820_, _14799_, _14591_);
  nand (_15821_, _14593_, _24376_);
  nand (_24377_, _15821_, _15820_);
  nand (_15822_, _14802_, _14591_);
  nand (_15823_, _14593_, _24378_);
  nand (_24379_, _15823_, _15822_);
  nand (_15824_, _14805_, _14591_);
  nand (_15825_, _14593_, _24380_);
  nand (_24381_, _15825_, _15824_);
  nand (_15826_, _14808_, _14591_);
  nand (_15827_, _14593_, _24382_);
  nand (_24383_, _15827_, _15826_);
  nand (_15828_, _14587_, _14789_);
  nand (_15829_, _14589_, _24384_);
  nand (_24385_, _15829_, _15828_);
  nand (_15830_, _14792_, _14587_);
  nand (_15831_, _14589_, _24386_);
  nand (_24387_, _15831_, _15830_);
  nand (_15832_, _14795_, _14587_);
  nand (_15833_, _14589_, _24388_);
  nand (_24389_, _15833_, _15832_);
  nand (_15834_, _14799_, _14587_);
  nand (_15835_, _14589_, _24390_);
  nand (_24391_, _15835_, _15834_);
  nand (_15836_, _14802_, _14587_);
  nand (_15837_, _14589_, _24392_);
  nand (_24393_, _15837_, _15836_);
  nand (_15838_, _14805_, _14587_);
  nand (_15839_, _14589_, _24394_);
  nand (_24395_, _15839_, _15838_);
  nand (_15840_, _14808_, _14587_);
  nand (_15841_, _14589_, _24396_);
  nand (_24397_, _15841_, _15840_);
  nand (_15842_, _14581_, _14789_);
  nand (_15843_, _14583_, _24399_);
  nand (_24400_, _15843_, _15842_);
  nand (_15844_, _14792_, _14581_);
  nand (_15845_, _14583_, _24401_);
  nand (_24402_, _15845_, _15844_);
  nand (_15846_, _14795_, _14581_);
  nand (_15847_, _14583_, _24403_);
  nand (_24404_, _15847_, _15846_);
  nand (_15848_, _14799_, _14581_);
  nand (_15849_, _14583_, _24405_);
  nand (_24406_, _15849_, _15848_);
  nand (_15851_, _14802_, _14581_);
  nand (_15852_, _14583_, _24407_);
  nand (_24408_, _15852_, _15851_);
  nand (_15853_, _14805_, _14581_);
  nand (_15854_, _14583_, _24409_);
  nand (_24410_, _15854_, _15853_);
  nand (_15855_, _14808_, _14581_);
  nand (_15856_, _14583_, _24411_);
  nand (_24412_, _15856_, _15855_);
  nand (_15857_, _14577_, _14789_);
  nand (_15859_, _14579_, _24413_);
  nand (_24414_, _15859_, _15857_);
  nand (_15860_, _14792_, _14577_);
  nand (_15861_, _14579_, _24415_);
  nand (_24416_, _15861_, _15860_);
  nand (_15862_, _14795_, _14577_);
  nand (_15863_, _14579_, _24417_);
  nand (_24418_, _15863_, _15862_);
  nand (_15864_, _14799_, _14577_);
  nand (_15865_, _14579_, _24419_);
  nand (_24420_, _15865_, _15864_);
  nand (_15866_, _14802_, _14577_);
  nand (_15867_, _14579_, _24421_);
  nand (_24422_, _15867_, _15866_);
  nand (_15868_, _14805_, _14577_);
  nand (_15869_, _14579_, _24423_);
  nand (_24424_, _15869_, _15868_);
  nand (_15870_, _14808_, _14577_);
  nand (_15871_, _14579_, _24425_);
  nand (_24426_, _15871_, _15870_);
  nand (_15872_, _14573_, _14789_);
  nand (_15873_, _14575_, _24427_);
  nand (_24428_, _15873_, _15872_);
  nand (_15874_, _14792_, _14573_);
  nand (_15875_, _14575_, _24429_);
  nand (_24430_, _15875_, _15874_);
  nand (_15876_, _14795_, _14573_);
  nand (_15877_, _14575_, _24431_);
  nand (_24432_, _15877_, _15876_);
  nand (_15878_, _14799_, _14573_);
  nand (_15879_, _14575_, _24433_);
  nand (_24434_, _15879_, _15878_);
  nand (_15880_, _14802_, _14573_);
  nand (_15881_, _14575_, _24435_);
  nand (_24436_, _15881_, _15880_);
  nand (_15882_, _14805_, _14573_);
  nand (_15883_, _14575_, _24437_);
  nand (_24438_, _15883_, _15882_);
  nand (_15884_, _14808_, _14573_);
  nand (_15885_, _14575_, _24440_);
  nand (_24441_, _15885_, _15884_);
  nand (_15887_, _14569_, _14789_);
  nand (_15888_, _14571_, _24442_);
  nand (_24443_, _15888_, _15887_);
  nand (_15889_, _14792_, _14569_);
  nand (_15890_, _14571_, _24444_);
  nand (_24445_, _15890_, _15889_);
  nand (_15891_, _14795_, _14569_);
  nand (_15892_, _14571_, _24446_);
  nand (_24447_, _15892_, _15891_);
  nand (_15894_, _14799_, _14569_);
  nand (_15895_, _14571_, _24448_);
  nand (_24449_, _15895_, _15894_);
  nand (_15896_, _14802_, _14569_);
  nand (_15897_, _14571_, _24450_);
  nand (_24451_, _15897_, _15896_);
  nand (_15898_, _14805_, _14569_);
  nand (_15899_, _14571_, _24452_);
  nand (_24453_, _15899_, _15898_);
  nand (_15900_, _14808_, _14569_);
  nand (_15901_, _14571_, _24454_);
  nand (_24455_, _15901_, _15900_);
  nand (_15902_, _14564_, _14789_);
  nand (_15903_, _14567_, _24456_);
  nand (_24457_, _15903_, _15902_);
  nand (_15904_, _14792_, _14564_);
  nand (_15905_, _14567_, _24458_);
  nand (_24459_, _15905_, _15904_);
  nand (_15906_, _14795_, _14564_);
  nand (_15907_, _14567_, _24460_);
  nand (_24461_, _15907_, _15906_);
  nand (_15908_, _14799_, _14564_);
  nand (_15909_, _14567_, _24462_);
  nand (_24463_, _15909_, _15908_);
  nand (_15910_, _14802_, _14564_);
  nand (_15911_, _14567_, _24464_);
  nand (_24465_, _15911_, _15910_);
  nand (_15912_, _14805_, _14564_);
  nand (_15913_, _14567_, _24466_);
  nand (_24467_, _15913_, _15912_);
  nand (_15914_, _14808_, _14564_);
  nand (_15915_, _14567_, _24468_);
  nand (_24469_, _15915_, _15914_);
  nand (_15916_, _14560_, _14789_);
  nand (_15917_, _14562_, _24470_);
  nand (_24471_, _15917_, _15916_);
  nand (_15918_, _14792_, _14560_);
  nand (_15919_, _14562_, _24472_);
  nand (_24473_, _15919_, _15918_);
  nand (_15920_, _14795_, _14560_);
  nand (_15922_, _14562_, _24474_);
  nand (_24475_, _15922_, _15920_);
  nand (_15923_, _14799_, _14560_);
  nand (_15924_, _14562_, _24476_);
  nand (_24477_, _15924_, _15923_);
  nand (_15925_, _14802_, _14560_);
  nand (_15926_, _14562_, _24478_);
  nand (_24479_, _15926_, _15925_);
  nand (_15927_, _14805_, _14560_);
  nand (_15928_, _14562_, _24481_);
  nand (_24482_, _15928_, _15927_);
  nand (_15930_, _14808_, _14560_);
  nand (_15931_, _14562_, _24483_);
  nand (_24484_, _15931_, _15930_);
  nand (_15932_, _14556_, _14789_);
  nand (_15933_, _14558_, _24485_);
  nand (_24486_, _15933_, _15932_);
  nand (_15934_, _14792_, _14556_);
  nand (_15935_, _14558_, _24487_);
  nand (_24488_, _15935_, _15934_);
  nand (_15936_, _14795_, _14556_);
  nand (_15937_, _14558_, _24489_);
  nand (_24490_, _15937_, _15936_);
  nand (_15938_, _14799_, _14556_);
  nand (_15939_, _14558_, _24491_);
  nand (_24492_, _15939_, _15938_);
  nand (_15940_, _14802_, _14556_);
  nand (_15941_, _14558_, _24493_);
  nand (_24494_, _15941_, _15940_);
  nand (_15942_, _14805_, _14556_);
  nand (_15943_, _14558_, _24495_);
  nand (_24496_, _15943_, _15942_);
  nand (_15944_, _14808_, _14556_);
  nand (_15945_, _14558_, _24497_);
  nand (_24498_, _15945_, _15944_);
  nand (_15946_, _14552_, _14789_);
  nand (_15947_, _14554_, _24499_);
  nand (_24500_, _15947_, _15946_);
  nand (_15948_, _14792_, _14552_);
  nand (_15949_, _14554_, _24501_);
  nand (_24502_, _15949_, _15948_);
  nand (_15950_, _14795_, _14552_);
  nand (_15951_, _14554_, _24503_);
  nand (_24504_, _15951_, _15950_);
  nand (_15952_, _14799_, _14552_);
  nand (_15953_, _14554_, _24505_);
  nand (_24506_, _15953_, _15952_);
  nand (_15954_, _14802_, _14552_);
  nand (_15955_, _14554_, _24507_);
  nand (_24508_, _15955_, _15954_);
  nand (_15957_, _14805_, _14552_);
  nand (_15958_, _14554_, _24509_);
  nand (_24510_, _15958_, _15957_);
  nand (_15959_, _14808_, _14552_);
  nand (_15960_, _14554_, _24511_);
  nand (_24512_, _15960_, _15959_);
  nand (_15961_, _14548_, _14789_);
  nand (_15962_, _14550_, _24513_);
  nand (_24514_, _15962_, _15961_);
  nand (_15963_, _14792_, _14548_);
  nand (_15965_, _14550_, _24515_);
  nand (_24516_, _15965_, _15963_);
  nand (_15966_, _14795_, _14548_);
  nand (_15967_, _14550_, _24517_);
  nand (_24518_, _15967_, _15966_);
  nand (_15968_, _14799_, _14548_);
  nand (_15969_, _14550_, _24519_);
  nand (_24520_, _15969_, _15968_);
  nand (_15970_, _14802_, _14548_);
  nand (_15971_, _14550_, _24523_);
  nand (_24524_, _15971_, _15970_);
  nand (_15973_, _14805_, _14548_);
  nand (_15974_, _14550_, _24525_);
  nand (_24526_, _15974_, _15973_);
  nand (_15975_, _14808_, _14548_);
  nand (_15976_, _14550_, _24527_);
  nand (_24528_, _15976_, _15975_);
  nand (_15977_, _14544_, _14789_);
  nand (_15978_, _14546_, _24529_);
  nand (_24530_, _15978_, _15977_);
  nand (_15979_, _14792_, _14544_);
  nand (_15980_, _14546_, _24531_);
  nand (_24532_, _15980_, _15979_);
  nand (_15981_, _14795_, _14544_);
  nand (_15982_, _14546_, _24533_);
  nand (_24534_, _15982_, _15981_);
  nand (_15983_, _14799_, _14544_);
  nand (_15984_, _14546_, _24535_);
  nand (_24536_, _15984_, _15983_);
  nand (_15985_, _14802_, _14544_);
  nand (_15986_, _14546_, _24537_);
  nand (_24538_, _15986_, _15985_);
  nand (_15987_, _14805_, _14544_);
  nand (_15988_, _14546_, _24539_);
  nand (_24540_, _15988_, _15987_);
  nand (_15989_, _14808_, _14544_);
  nand (_15990_, _14546_, _24541_);
  nand (_24542_, _15990_, _15989_);
  nand (_15991_, _14538_, _14789_);
  nand (_15992_, _14542_, _24543_);
  nand (_24544_, _15992_, _15991_);
  nand (_15993_, _14792_, _14538_);
  nand (_15994_, _14542_, _24545_);
  nand (_24546_, _15994_, _15993_);
  nand (_15995_, _14795_, _14538_);
  nand (_15996_, _14542_, _24547_);
  nand (_24548_, _15996_, _15995_);
  nand (_15997_, _14799_, _14538_);
  nand (_15998_, _14542_, _24549_);
  nand (_24550_, _15998_, _15997_);
  nand (_16000_, _14802_, _14538_);
  nand (_16001_, _14542_, _24551_);
  nand (_24552_, _16001_, _16000_);
  nand (_16002_, _14805_, _14538_);
  nand (_16003_, _14542_, _24553_);
  nand (_24554_, _16003_, _16002_);
  nand (_16004_, _14808_, _14538_);
  nand (_16005_, _14542_, _24555_);
  nand (_24556_, _16005_, _16004_);
  nand (_16006_, _14534_, _14789_);
  nand (_16008_, _14536_, _24557_);
  nand (_24558_, _16008_, _16006_);
  nand (_16009_, _14792_, _14534_);
  nand (_16010_, _14536_, _24559_);
  nand (_24560_, _16010_, _16009_);
  nand (_16011_, _14795_, _14534_);
  nand (_16012_, _14536_, _24561_);
  nand (_24562_, _16012_, _16011_);
  nand (_16013_, _14799_, _14534_);
  nand (_16014_, _14536_, _24564_);
  nand (_24565_, _16014_, _16013_);
  nand (_16015_, _14802_, _14534_);
  nand (_16016_, _14536_, _24566_);
  nand (_24567_, _16016_, _16015_);
  nand (_16017_, _14805_, _14534_);
  nand (_16018_, _14536_, _24568_);
  nand (_24569_, _16018_, _16017_);
  nand (_16019_, _14808_, _14534_);
  nand (_16020_, _14536_, _24570_);
  nand (_24571_, _16020_, _16019_);
  nand (_16021_, _14529_, _14789_);
  nand (_16022_, _14532_, _24572_);
  nand (_24573_, _16022_, _16021_);
  nand (_16023_, _14792_, _14529_);
  nand (_16024_, _14532_, _24574_);
  nand (_24575_, _16024_, _16023_);
  nand (_16025_, _14795_, _14529_);
  nand (_16026_, _14532_, _24576_);
  nand (_24577_, _16026_, _16025_);
  nand (_16027_, _14799_, _14529_);
  nand (_16028_, _14532_, _24578_);
  nand (_24579_, _16028_, _16027_);
  nand (_16029_, _14802_, _14529_);
  nand (_16030_, _14532_, _24580_);
  nand (_24581_, _16030_, _16029_);
  nand (_16031_, _14805_, _14529_);
  nand (_16032_, _14532_, _24582_);
  nand (_24583_, _16032_, _16031_);
  nand (_16033_, _14808_, _14529_);
  nand (_16034_, _14532_, _24584_);
  nand (_24585_, _16034_, _16033_);
  nand (_16036_, _14525_, _14789_);
  nand (_16037_, _14527_, _24586_);
  nand (_24587_, _16037_, _16036_);
  nand (_16038_, _14792_, _14525_);
  nand (_16039_, _14527_, _24588_);
  nand (_24589_, _16039_, _16038_);
  nand (_16040_, _14795_, _14525_);
  nand (_16041_, _14527_, _24590_);
  nand (_24591_, _16041_, _16040_);
  nand (_16043_, _14799_, _14525_);
  nand (_16044_, _14527_, _24592_);
  nand (_24593_, _16044_, _16043_);
  nand (_16045_, _14802_, _14525_);
  nand (_16046_, _14527_, _24594_);
  nand (_24595_, _16046_, _16045_);
  nand (_16047_, _14805_, _14525_);
  nand (_16048_, _14527_, _24596_);
  nand (_24597_, _16048_, _16047_);
  nand (_16049_, _14808_, _14525_);
  nand (_16050_, _14527_, _24598_);
  nand (_24599_, _16050_, _16049_);
  nand (_16051_, _14521_, _14789_);
  nand (_16052_, _14523_, _24600_);
  nand (_24601_, _16052_, _16051_);
  nand (_16053_, _14792_, _14521_);
  nand (_16054_, _14523_, _24602_);
  nand (_24603_, _16054_, _16053_);
  nand (_16055_, _14795_, _14521_);
  nand (_16056_, _14523_, _24605_);
  nand (_24606_, _16056_, _16055_);
  nand (_16057_, _14799_, _14521_);
  nand (_16058_, _14523_, _24607_);
  nand (_24608_, _16058_, _16057_);
  nand (_16059_, _14802_, _14521_);
  nand (_16060_, _14523_, _24609_);
  nand (_24610_, _16060_, _16059_);
  nand (_16061_, _14805_, _14521_);
  nand (_16062_, _14523_, _24611_);
  nand (_24612_, _16062_, _16061_);
  nand (_16063_, _14808_, _14521_);
  nand (_16064_, _14523_, _24613_);
  nand (_24614_, _16064_, _16063_);
  nand (_16065_, _14517_, _14789_);
  nand (_16066_, _14519_, _24615_);
  nand (_24616_, _16066_, _16065_);
  nand (_16067_, _14792_, _14517_);
  nand (_16068_, _14519_, _24617_);
  nand (_24618_, _16068_, _16067_);
  nand (_16069_, _14795_, _14517_);
  nand (_16071_, _14519_, _24619_);
  nand (_24620_, _16071_, _16069_);
  nand (_16072_, _14799_, _14517_);
  nand (_16073_, _14519_, _24621_);
  nand (_24622_, _16073_, _16072_);
  nand (_16074_, _14802_, _14517_);
  nand (_16075_, _14519_, _24623_);
  nand (_24624_, _16075_, _16074_);
  nand (_16076_, _14805_, _14517_);
  nand (_16077_, _14519_, _24625_);
  nand (_24626_, _16077_, _16076_);
  nand (_16079_, _14808_, _14517_);
  nand (_16080_, _14519_, _24627_);
  nand (_24628_, _16080_, _16079_);
  nand (_16081_, _14510_, _24629_);
  nand (_16082_, _14509_, _14789_);
  nand (_24630_, _16082_, _16081_);
  nand (_16083_, _14510_, _24631_);
  nand (_16084_, _14792_, _14509_);
  nand (_24632_, _16084_, _16083_);
  nand (_16085_, _14510_, _24633_);
  nand (_16086_, _14795_, _14509_);
  nand (_24634_, _16086_, _16085_);
  nand (_16087_, _14510_, _24635_);
  nand (_16088_, _14799_, _14509_);
  nand (_24636_, _16088_, _16087_);
  nand (_16089_, _14510_, _24637_);
  nand (_16090_, _14802_, _14509_);
  nand (_24638_, _16090_, _16089_);
  nand (_16091_, _14510_, _24639_);
  nand (_16092_, _14805_, _14509_);
  nand (_24640_, _16092_, _16091_);
  nand (_16093_, _14510_, _24641_);
  nand (_16094_, _14808_, _14509_);
  nand (_24642_, _16094_, _16093_);
  nand (_16095_, _14506_, _24643_);
  nand (_16096_, _14505_, _14789_);
  nand (_24644_, _16096_, _16095_);
  nand (_16097_, _14506_, _24646_);
  nand (_16098_, _14792_, _14505_);
  nand (_24647_, _16098_, _16097_);
  nand (_16099_, _14506_, _24648_);
  nand (_16100_, _14795_, _14505_);
  nand (_24649_, _16100_, _16099_);
  nand (_16101_, _14506_, _24650_);
  nand (_16102_, _14799_, _14505_);
  nand (_24651_, _16102_, _16101_);
  nand (_16103_, _14506_, _24652_);
  nand (_16104_, _14802_, _14505_);
  nand (_24653_, _16104_, _16103_);
  nand (_16106_, _14506_, _24654_);
  nand (_16107_, _14805_, _14505_);
  nand (_24655_, _16107_, _16106_);
  nand (_16108_, _14506_, _24656_);
  nand (_16109_, _14808_, _14505_);
  nand (_24657_, _16109_, _16108_);
  nand (_16110_, _14502_, _24658_);
  nand (_16111_, _14501_, _14789_);
  nand (_24659_, _16111_, _16110_);
  nand (_16112_, _14502_, _24660_);
  nand (_16114_, _14792_, _14501_);
  nand (_24661_, _16114_, _16112_);
  nand (_16115_, _14502_, _24662_);
  nand (_16116_, _14795_, _14501_);
  nand (_24663_, _16116_, _16115_);
  nand (_16117_, _14502_, _24664_);
  nand (_16118_, _14799_, _14501_);
  nand (_24665_, _16118_, _16117_);
  nand (_16119_, _14502_, _24666_);
  nand (_16120_, _14802_, _14501_);
  nand (_24667_, _16120_, _16119_);
  nand (_16121_, _14502_, _24668_);
  nand (_16122_, _14805_, _14501_);
  nand (_24669_, _16122_, _16121_);
  nand (_16123_, _14502_, _24670_);
  nand (_16124_, _14808_, _14501_);
  nand (_24671_, _16124_, _16123_);
  nand (_16125_, _14498_, _24672_);
  nand (_16126_, _14496_, _14789_);
  nand (_24673_, _16126_, _16125_);
  nand (_16127_, _14498_, _24674_);
  nand (_16128_, _14792_, _14496_);
  nand (_24675_, _16128_, _16127_);
  nand (_16129_, _14498_, _24676_);
  nand (_16130_, _14795_, _14496_);
  nand (_24677_, _16130_, _16129_);
  nand (_16131_, _14498_, _24678_);
  nand (_16132_, _14799_, _14496_);
  nand (_24679_, _16132_, _16131_);
  nand (_16133_, _14498_, _24680_);
  nand (_16134_, _14802_, _14496_);
  nand (_24681_, _16134_, _16133_);
  nand (_16135_, _14498_, _24682_);
  nand (_16136_, _14805_, _14496_);
  nand (_24683_, _16136_, _16135_);
  nand (_16137_, _14498_, _24684_);
  nand (_16138_, _14808_, _14496_);
  nand (_24685_, _16138_, _16137_);
  nand (_16139_, _14493_, _24687_);
  nand (_16140_, _14492_, _14789_);
  nand (_24688_, _16140_, _16139_);
  nand (_16141_, _14493_, _24689_);
  nand (_16142_, _14792_, _14492_);
  nand (_24690_, _16142_, _16141_);
  nand (_16143_, _14493_, _24691_);
  nand (_16144_, _14795_, _14492_);
  nand (_24692_, _16144_, _16143_);
  nand (_16145_, _14493_, _24693_);
  nand (_16146_, _14799_, _14492_);
  nand (_24694_, _16146_, _16145_);
  nand (_16147_, _14493_, _24695_);
  nand (_16148_, _14802_, _14492_);
  nand (_24696_, _16148_, _16147_);
  nand (_16149_, _14493_, _24697_);
  nand (_16150_, _14805_, _14492_);
  nand (_24698_, _16150_, _16149_);
  nand (_16151_, _14493_, _24699_);
  nand (_16152_, _14808_, _14492_);
  nand (_24700_, _16152_, _16151_);
  nand (_16153_, _14489_, _24701_);
  nand (_16154_, _14488_, _14789_);
  nand (_24702_, _16154_, _16153_);
  nand (_16155_, _14489_, _24703_);
  nand (_16156_, _14792_, _14488_);
  nand (_24704_, _16156_, _16155_);
  nand (_16157_, _14489_, _24705_);
  nand (_16158_, _14795_, _14488_);
  nand (_24706_, _16158_, _16157_);
  nand (_16159_, _14489_, _24707_);
  nand (_16160_, _14799_, _14488_);
  nand (_24708_, _16160_, _16159_);
  nand (_16162_, _14489_, _24709_);
  nand (_16163_, _14802_, _14488_);
  nand (_24710_, _16163_, _16162_);
  nand (_16164_, _14489_, _24711_);
  nand (_16165_, _14805_, _14488_);
  nand (_24712_, _16165_, _16164_);
  nand (_16166_, _14489_, _24713_);
  nand (_16167_, _14808_, _14488_);
  nand (_24714_, _16167_, _16166_);
  nand (_16169_, _14485_, _24715_);
  nand (_16170_, _14484_, _14789_);
  nand (_24716_, _16170_, _16169_);
  nand (_16171_, _14485_, _24717_);
  nand (_16172_, _14792_, _14484_);
  nand (_24718_, _16172_, _16171_);
  nand (_16173_, _14485_, _24719_);
  nand (_16174_, _14795_, _14484_);
  nand (_24720_, _16174_, _16173_);
  nand (_16175_, _14485_, _24721_);
  nand (_16176_, _14799_, _14484_);
  nand (_24722_, _16176_, _16175_);
  nand (_16177_, _14485_, _24723_);
  nand (_16178_, _14802_, _14484_);
  nand (_24724_, _16178_, _16177_);
  nand (_16179_, _14485_, _24725_);
  nand (_16180_, _14805_, _14484_);
  nand (_24726_, _16180_, _16179_);
  nand (_16181_, _14485_, _24728_);
  nand (_16182_, _14808_, _14484_);
  nand (_24729_, _16182_, _16181_);
  nand (_16183_, _14481_, _24730_);
  nand (_16184_, _14480_, _14789_);
  nand (_24731_, _16184_, _16183_);
  nand (_16185_, _14481_, _24732_);
  nand (_16186_, _14792_, _14480_);
  nand (_24733_, _16186_, _16185_);
  nand (_16187_, _14481_, _24734_);
  nand (_16188_, _14795_, _14480_);
  nand (_24735_, _16188_, _16187_);
  nand (_16190_, _14481_, _24736_);
  nand (_16191_, _14799_, _14480_);
  nand (_24737_, _16191_, _16190_);
  nand (_16192_, _14481_, _24738_);
  nand (_16193_, _14802_, _14480_);
  nand (_24739_, _16193_, _16192_);
  nand (_16194_, _14481_, _24740_);
  nand (_16195_, _14805_, _14480_);
  nand (_24741_, _16195_, _16194_);
  nand (_16196_, _14481_, _24742_);
  nand (_16198_, _14808_, _14480_);
  nand (_24743_, _16198_, _16196_);
  nand (_16199_, _14477_, _24744_);
  nand (_16200_, _14476_, _14789_);
  nand (_24745_, _16200_, _16199_);
  nand (_16201_, _14477_, _24746_);
  nand (_16202_, _14792_, _14476_);
  nand (_24747_, _16202_, _16201_);
  nand (_16203_, _14477_, _24748_);
  nand (_16204_, _14795_, _14476_);
  nand (_24749_, _16204_, _16203_);
  nand (_16205_, _14477_, _24750_);
  nand (_16206_, _14799_, _14476_);
  nand (_24751_, _16206_, _16205_);
  nand (_16207_, _14477_, _24752_);
  nand (_16208_, _14802_, _14476_);
  nand (_24753_, _16208_, _16207_);
  nand (_16209_, _14477_, _24754_);
  nand (_16210_, _14805_, _14476_);
  nand (_24755_, _16210_, _16209_);
  nand (_16211_, _14477_, _24756_);
  nand (_16212_, _14808_, _14476_);
  nand (_24757_, _16212_, _16211_);
  nand (_16213_, _14473_, _24758_);
  nand (_16214_, _14472_, _14789_);
  nand (_24759_, _16214_, _16213_);
  nand (_16215_, _14473_, _24760_);
  nand (_16216_, _14792_, _14472_);
  nand (_24761_, _16216_, _16215_);
  nand (_16217_, _14473_, _24762_);
  nand (_16219_, _14795_, _14472_);
  nand (_24763_, _16219_, _16217_);
  nand (_16220_, _14473_, _24764_);
  nand (_16221_, _14799_, _14472_);
  nand (_24765_, _16221_, _16220_);
  nand (_16222_, _14473_, _24766_);
  nand (_16223_, _14802_, _14472_);
  nand (_24767_, _16223_, _16222_);
  nand (_16224_, _14473_, _24769_);
  nand (_16225_, _14805_, _14472_);
  nand (_24770_, _16225_, _16224_);
  nand (_16227_, _14473_, _24771_);
  nand (_16228_, _14808_, _14472_);
  nand (_24772_, _16228_, _16227_);
  nand (_16229_, _14469_, _24773_);
  nand (_16230_, _14468_, _14789_);
  nand (_24774_, _16230_, _16229_);
  nand (_16231_, _14469_, _24775_);
  nand (_16232_, _14792_, _14468_);
  nand (_24776_, _16232_, _16231_);
  nand (_16233_, _14469_, _24777_);
  nand (_16234_, _14795_, _14468_);
  nand (_24778_, _16234_, _16233_);
  nand (_16235_, _14469_, _24779_);
  nand (_16236_, _14799_, _14468_);
  nand (_24780_, _16236_, _16235_);
  nand (_16237_, _14469_, _24781_);
  nand (_16238_, _14802_, _14468_);
  nand (_24782_, _16238_, _16237_);
  nand (_16239_, _14469_, _24783_);
  nand (_16240_, _14805_, _14468_);
  nand (_24784_, _16240_, _16239_);
  nand (_16241_, _14469_, _24785_);
  nand (_16242_, _14808_, _14468_);
  nand (_24786_, _16242_, _16241_);
  nand (_16243_, _14465_, _24787_);
  nand (_16244_, _14463_, _14789_);
  nand (_24788_, _16244_, _16243_);
  nand (_16245_, _14465_, _24789_);
  nand (_16246_, _14792_, _14463_);
  nand (_24790_, _16246_, _16245_);
  nand (_16248_, _14465_, _24791_);
  nand (_16249_, _14795_, _14463_);
  nand (_24792_, _16249_, _16248_);
  nand (_16250_, _14465_, _24793_);
  nand (_16251_, _14799_, _14463_);
  nand (_24794_, _16251_, _16250_);
  nand (_16252_, _14465_, _24795_);
  nand (_16253_, _14802_, _14463_);
  nand (_24796_, _16253_, _16252_);
  nand (_16256_, _14465_, _24797_);
  nand (_16257_, _14805_, _14463_);
  nand (_24798_, _16257_, _16256_);
  nand (_16258_, _14465_, _24799_);
  nand (_16259_, _14808_, _14463_);
  nand (_24800_, _16259_, _16258_);
  nand (_16260_, _14460_, _24801_);
  nand (_16261_, _14459_, _14789_);
  nand (_24802_, _16261_, _16260_);
  nand (_16262_, _14460_, _24803_);
  nand (_16263_, _14792_, _14459_);
  nand (_24804_, _16263_, _16262_);
  nand (_16264_, _14460_, _24805_);
  nand (_16265_, _14795_, _14459_);
  nand (_24806_, _16265_, _16264_);
  nand (_16266_, _14460_, _24807_);
  nand (_16267_, _14799_, _14459_);
  nand (_24808_, _16267_, _16266_);
  nand (_16268_, _14460_, _24810_);
  nand (_16269_, _14802_, _14459_);
  nand (_24811_, _16269_, _16268_);
  nand (_16270_, _14460_, _24812_);
  nand (_16271_, _14805_, _14459_);
  nand (_24813_, _16271_, _16270_);
  nand (_16272_, _14460_, _24814_);
  nand (_16273_, _14808_, _14459_);
  nand (_24815_, _16273_, _16272_);
  nand (_16274_, _14456_, _24816_);
  nand (_16275_, _14455_, _14789_);
  nand (_24817_, _16275_, _16274_);
  nand (_16277_, _14456_, _24818_);
  nand (_16278_, _14792_, _14455_);
  nand (_24819_, _16278_, _16277_);
  nand (_16279_, _14456_, _24820_);
  nand (_16280_, _14795_, _14455_);
  nand (_24821_, _16280_, _16279_);
  nand (_16281_, _14456_, _24822_);
  nand (_16282_, _14799_, _14455_);
  nand (_24823_, _16282_, _16281_);
  nand (_16283_, _14456_, _24824_);
  nand (_16285_, _14802_, _14455_);
  nand (_24825_, _16285_, _16283_);
  nand (_16286_, _14456_, _24826_);
  nand (_16287_, _14805_, _14455_);
  nand (_24827_, _16287_, _16286_);
  nand (_16288_, _14456_, _24828_);
  nand (_16289_, _14808_, _14455_);
  nand (_24829_, _16289_, _16288_);
  nand (_16290_, _14452_, _24830_);
  nand (_16291_, _14451_, _14789_);
  nand (_24831_, _16291_, _16290_);
  nand (_16292_, _14452_, _24832_);
  nand (_16293_, _14792_, _14451_);
  nand (_24833_, _16293_, _16292_);
  nand (_16294_, _14452_, _24834_);
  nand (_16295_, _14795_, _14451_);
  nand (_24835_, _16295_, _16294_);
  nand (_16296_, _14452_, _24836_);
  nand (_16297_, _14799_, _14451_);
  nand (_24837_, _16297_, _16296_);
  nand (_16298_, _14452_, _24838_);
  nand (_16299_, _14802_, _14451_);
  nand (_24839_, _16299_, _16298_);
  nand (_16300_, _14452_, _24840_);
  nand (_16301_, _14805_, _14451_);
  nand (_24841_, _16301_, _16300_);
  nand (_16302_, _14452_, _24842_);
  nand (_16303_, _14808_, _14451_);
  nand (_24843_, _16303_, _16302_);
  nand (_16304_, _14448_, _24844_);
  nand (_16306_, _14447_, _14789_);
  nand (_24845_, _16306_, _16304_);
  nand (_16307_, _14448_, _24846_);
  nand (_16308_, _14792_, _14447_);
  nand (_24847_, _16308_, _16307_);
  nand (_16309_, _14448_, _24848_);
  nand (_16310_, _14795_, _14447_);
  nand (_24849_, _16310_, _16309_);
  nand (_16311_, _14448_, _24851_);
  nand (_16312_, _14799_, _14447_);
  nand (_24852_, _16312_, _16311_);
  nand (_16314_, _14448_, _24853_);
  nand (_16315_, _14802_, _14447_);
  nand (_24854_, _16315_, _16314_);
  nand (_16316_, _14448_, _24855_);
  nand (_16317_, _14805_, _14447_);
  nand (_24856_, _16317_, _16316_);
  nand (_16318_, _14448_, _24857_);
  nand (_16319_, _14808_, _14447_);
  nand (_24858_, _16319_, _16318_);
  nand (_16320_, _14442_, _24859_);
  nand (_16321_, _14441_, _14789_);
  nand (_24860_, _16321_, _16320_);
  nand (_16322_, _14442_, _24861_);
  nand (_16323_, _14792_, _14441_);
  nand (_24862_, _16323_, _16322_);
  nand (_16324_, _14442_, _24863_);
  nand (_16325_, _14795_, _14441_);
  nand (_24864_, _16325_, _16324_);
  nand (_16326_, _14442_, _24865_);
  nand (_16327_, _14799_, _14441_);
  nand (_24866_, _16327_, _16326_);
  nand (_16328_, _14442_, _24867_);
  nand (_16329_, _14802_, _14441_);
  nand (_24868_, _16329_, _16328_);
  nand (_16330_, _14442_, _24869_);
  nand (_16331_, _14805_, _14441_);
  nand (_24870_, _16331_, _16330_);
  nand (_16332_, _14442_, _24871_);
  nand (_16333_, _14808_, _14441_);
  nand (_24872_, _16333_, _16332_);
  nand (_16335_, _14438_, _24873_);
  nand (_16336_, _14437_, _14789_);
  nand (_24874_, _16336_, _16335_);
  nand (_16337_, _14438_, _24875_);
  nand (_16338_, _14792_, _14437_);
  nand (_24876_, _16338_, _16337_);
  nand (_16339_, _14438_, _24877_);
  nand (_16340_, _14795_, _14437_);
  nand (_24878_, _16340_, _16339_);
  nand (_16342_, _14438_, _24879_);
  nand (_16343_, _14799_, _14437_);
  nand (_24880_, _16343_, _16342_);
  nand (_16344_, _14438_, _24881_);
  nand (_16345_, _14802_, _14437_);
  nand (_24882_, _16345_, _16344_);
  nand (_16346_, _14438_, _24883_);
  nand (_16347_, _14805_, _14437_);
  nand (_24884_, _16347_, _16346_);
  nand (_16348_, _14438_, _24885_);
  nand (_16349_, _14808_, _14437_);
  nand (_24886_, _16349_, _16348_);
  nand (_16350_, _14434_, _24887_);
  nand (_16351_, _14433_, _14789_);
  nand (_24888_, _16351_, _16350_);
  nand (_16352_, _14434_, _24889_);
  nand (_16353_, _14792_, _14433_);
  nand (_24890_, _16353_, _16352_);
  nand (_16354_, _14434_, _24892_);
  nand (_16355_, _14795_, _14433_);
  nand (_24893_, _16355_, _16354_);
  nand (_16356_, _14434_, _24894_);
  nand (_16357_, _14799_, _14433_);
  nand (_24895_, _16357_, _16356_);
  nand (_16358_, _14434_, _24896_);
  nand (_16359_, _14802_, _14433_);
  nand (_24897_, _16359_, _16358_);
  nand (_16360_, _14434_, _24898_);
  nand (_16361_, _14805_, _14433_);
  nand (_24899_, _16361_, _16360_);
  nand (_16363_, _14434_, _24900_);
  nand (_16364_, _14808_, _14433_);
  nand (_24901_, _16364_, _16363_);
  nand (_16365_, _14429_, _24902_);
  nand (_16366_, _14428_, _14789_);
  nand (_24903_, _16366_, _16365_);
  nand (_16367_, _14429_, _24904_);
  nand (_16368_, _14792_, _14428_);
  nand (_24905_, _16368_, _16367_);
  nand (_16369_, _14429_, _24906_);
  nand (_16371_, _14795_, _14428_);
  nand (_24907_, _16371_, _16369_);
  nand (_16372_, _14429_, _24908_);
  nand (_16373_, _14799_, _14428_);
  nand (_24909_, _16373_, _16372_);
  nand (_16374_, _14429_, _24910_);
  nand (_16375_, _14802_, _14428_);
  nand (_24911_, _16375_, _16374_);
  nand (_16376_, _14429_, _24912_);
  nand (_16377_, _14805_, _14428_);
  nand (_24913_, _16377_, _16376_);
  nand (_16378_, _14429_, _24914_);
  nand (_16379_, _14808_, _14428_);
  nand (_24915_, _16379_, _16378_);
  nand (_16380_, _14425_, _24916_);
  nand (_16381_, _14424_, _14789_);
  nand (_24917_, _16381_, _16380_);
  nand (_16382_, _14425_, _24918_);
  nand (_16383_, _14792_, _14424_);
  nand (_24919_, _16383_, _16382_);
  nand (_16384_, _14425_, _24920_);
  nand (_16385_, _14795_, _14424_);
  nand (_24921_, _16385_, _16384_);
  nand (_16386_, _14425_, _24922_);
  nand (_16387_, _14799_, _14424_);
  nand (_24923_, _16387_, _16386_);
  nand (_16388_, _14425_, _24924_);
  nand (_16389_, _14802_, _14424_);
  nand (_24925_, _16389_, _16388_);
  nand (_16390_, _14425_, _24926_);
  nand (_16392_, _14805_, _14424_);
  nand (_24927_, _16392_, _16390_);
  nand (_16393_, _14425_, _24928_);
  nand (_16394_, _14808_, _14424_);
  nand (_24929_, _16394_, _16393_);
  nand (_16395_, _14421_, _24930_);
  nand (_16396_, _14420_, _14789_);
  nand (_24931_, _16396_, _16395_);
  nand (_16397_, _14421_, _24934_);
  nand (_16398_, _14792_, _14420_);
  nand (_24935_, _16398_, _16397_);
  nand (_16400_, _14421_, _24936_);
  nand (_16401_, _14795_, _14420_);
  nand (_24937_, _16401_, _16400_);
  nand (_16402_, _14421_, _24938_);
  nand (_16403_, _14799_, _14420_);
  nand (_24939_, _16403_, _16402_);
  nand (_16404_, _14421_, _24940_);
  nand (_16405_, _14802_, _14420_);
  nand (_24941_, _16405_, _16404_);
  nand (_16406_, _14421_, _24942_);
  nand (_16407_, _14805_, _14420_);
  nand (_24943_, _16407_, _16406_);
  nand (_16408_, _14421_, _24944_);
  nand (_16409_, _14808_, _14420_);
  nand (_24945_, _16409_, _16408_);
  nand (_16410_, _14417_, _24946_);
  nand (_16411_, _14416_, _14789_);
  nand (_24947_, _16411_, _16410_);
  nand (_16412_, _14417_, _24948_);
  nand (_16413_, _14792_, _14416_);
  nand (_24949_, _16413_, _16412_);
  nand (_16414_, _14417_, _24950_);
  nand (_16415_, _14795_, _14416_);
  nand (_24951_, _16415_, _16414_);
  nand (_16416_, _14417_, _24952_);
  nand (_16417_, _14799_, _14416_);
  nand (_24953_, _16417_, _16416_);
  nand (_16418_, _14417_, _24954_);
  nand (_16419_, _14802_, _14416_);
  nand (_24955_, _16419_, _16418_);
  nand (_16421_, _14417_, _24956_);
  nand (_16422_, _14805_, _14416_);
  nand (_24957_, _16422_, _16421_);
  nand (_16423_, _14417_, _24958_);
  nand (_16424_, _14808_, _14416_);
  nand (_24959_, _16424_, _16423_);
  nand (_16425_, _14413_, _24960_);
  nand (_16426_, _14412_, _14789_);
  nand (_24961_, _16426_, _16425_);
  nand (_16428_, _14413_, _24962_);
  nand (_16429_, _14792_, _14412_);
  nand (_24963_, _16429_, _16428_);
  nand (_16430_, _14413_, _24964_);
  nand (_16431_, _14795_, _14412_);
  nand (_24965_, _16431_, _16430_);
  nand (_16432_, _14413_, _24966_);
  nand (_16433_, _14799_, _14412_);
  nand (_24967_, _16433_, _16432_);
  nand (_16434_, _14413_, _24968_);
  nand (_16435_, _14802_, _14412_);
  nand (_24969_, _16435_, _16434_);
  nand (_16436_, _14413_, _24970_);
  nand (_16437_, _14805_, _14412_);
  nand (_24971_, _16437_, _16436_);
  nand (_16438_, _14413_, _24972_);
  nand (_16439_, _14808_, _14412_);
  nand (_24973_, _16439_, _16438_);
  nand (_16440_, _14409_, _24975_);
  nand (_16441_, _14408_, _14789_);
  nand (_24976_, _16441_, _16440_);
  nand (_16442_, _14409_, _24977_);
  nand (_16443_, _14792_, _14408_);
  nand (_24978_, _16443_, _16442_);
  nand (_16444_, _14409_, _24979_);
  nand (_16445_, _14795_, _14408_);
  nand (_24980_, _16445_, _16444_);
  nand (_16446_, _14409_, _24981_);
  nand (_16447_, _14799_, _14408_);
  nand (_24982_, _16447_, _16446_);
  nand (_16449_, _14409_, _24983_);
  nand (_16450_, _14802_, _14408_);
  nand (_24984_, _16450_, _16449_);
  nand (_16451_, _14409_, _24985_);
  nand (_16452_, _14805_, _14408_);
  nand (_24986_, _16452_, _16451_);
  nand (_16453_, _14409_, _24987_);
  nand (_16454_, _14808_, _14408_);
  nand (_24988_, _16454_, _16453_);
  nand (_16455_, _14405_, _24989_);
  nand (_16457_, _14404_, _14789_);
  nand (_24990_, _16457_, _16455_);
  nand (_16458_, _14405_, _24991_);
  nand (_16459_, _14792_, _14404_);
  nand (_24992_, _16459_, _16458_);
  nand (_16460_, _14405_, _24993_);
  nand (_16461_, _14795_, _14404_);
  nand (_24994_, _16461_, _16460_);
  nand (_16462_, _14405_, _24995_);
  nand (_16463_, _14799_, _14404_);
  nand (_24996_, _16463_, _16462_);
  nand (_16464_, _14405_, _24997_);
  nand (_16465_, _14802_, _14404_);
  nand (_24998_, _16465_, _16464_);
  nand (_16466_, _14405_, _24999_);
  nand (_16467_, _14805_, _14404_);
  nand (_25000_, _16467_, _16466_);
  nand (_16468_, _14405_, _25001_);
  nand (_16469_, _14808_, _14404_);
  nand (_25002_, _16469_, _16468_);
  nand (_16470_, _14401_, _25003_);
  nand (_16471_, _14400_, _14789_);
  nand (_25004_, _16471_, _16470_);
  nand (_16472_, _14401_, _25005_);
  nand (_16473_, _14792_, _14400_);
  nand (_25006_, _16473_, _16472_);
  nand (_16474_, _14401_, _25007_);
  nand (_16475_, _14795_, _14400_);
  nand (_25008_, _16475_, _16474_);
  nand (_16476_, _14401_, _25009_);
  nand (_16478_, _14799_, _14400_);
  nand (_25010_, _16478_, _16476_);
  nand (_16479_, _14401_, _25011_);
  nand (_16480_, _14802_, _14400_);
  nand (_25012_, _16480_, _16479_);
  nand (_16481_, _14401_, _25013_);
  nand (_16482_, _14805_, _14400_);
  nand (_25014_, _16482_, _16481_);
  nand (_16483_, _14401_, _25016_);
  nand (_16484_, _14808_, _14400_);
  nand (_25017_, _16484_, _16483_);
  nand (_16486_, _14396_, _25018_);
  nand (_16487_, _14395_, _14789_);
  nand (_25019_, _16487_, _16486_);
  nand (_16488_, _14396_, _25020_);
  nand (_16489_, _14792_, _14395_);
  nand (_25021_, _16489_, _16488_);
  nand (_16490_, _14396_, _25022_);
  nand (_16491_, _14795_, _14395_);
  nand (_25023_, _16491_, _16490_);
  nand (_16492_, _14396_, _25024_);
  nand (_16493_, _14799_, _14395_);
  nand (_25025_, _16493_, _16492_);
  nand (_16494_, _14396_, _25026_);
  nand (_16495_, _14802_, _14395_);
  nand (_25027_, _16495_, _16494_);
  nand (_16496_, _14396_, _25028_);
  nand (_16497_, _14805_, _14395_);
  nand (_25029_, _16497_, _16496_);
  nand (_16498_, _14396_, _25030_);
  nand (_16499_, _14808_, _14395_);
  nand (_25031_, _16499_, _16498_);
  nand (_16500_, _14392_, _25032_);
  nand (_16501_, _14391_, _14789_);
  nand (_25033_, _16501_, _16500_);
  nand (_16502_, _14392_, _25034_);
  nand (_16503_, _14792_, _14391_);
  nand (_25035_, _16503_, _16502_);
  nand (_16504_, _14392_, _25036_);
  nand (_16505_, _14795_, _14391_);
  nand (_25037_, _16505_, _16504_);
  nand (_16507_, _14392_, _25038_);
  nand (_16508_, _14799_, _14391_);
  nand (_25039_, _16508_, _16507_);
  nand (_16509_, _14392_, _25040_);
  nand (_16510_, _14802_, _14391_);
  nand (_25041_, _16510_, _16509_);
  nand (_16511_, _14392_, _25042_);
  nand (_16512_, _14805_, _14391_);
  nand (_25043_, _16512_, _16511_);
  nand (_16514_, _14392_, _25044_);
  nand (_16515_, _14808_, _14391_);
  nand (_25045_, _16515_, _16514_);
  nand (_16516_, _14388_, _25046_);
  nand (_16517_, _14387_, _14789_);
  nand (_25047_, _16517_, _16516_);
  nand (_16518_, _14388_, _25048_);
  nand (_16519_, _14792_, _14387_);
  nand (_25049_, _16519_, _16518_);
  nand (_16520_, _14388_, _25050_);
  nand (_16521_, _14795_, _14387_);
  nand (_25051_, _16521_, _16520_);
  nand (_16522_, _14388_, _25052_);
  nand (_16523_, _14799_, _14387_);
  nand (_25053_, _16523_, _16522_);
  nand (_16524_, _14388_, _25054_);
  nand (_16525_, _14802_, _14387_);
  nand (_25055_, _16525_, _16524_);
  nand (_16526_, _14388_, _25057_);
  nand (_16527_, _14805_, _14387_);
  nand (_25058_, _16527_, _16526_);
  nand (_16528_, _14388_, _25059_);
  nand (_16529_, _14808_, _14387_);
  nand (_25060_, _16529_, _16528_);
  nand (_16530_, _14384_, _25061_);
  nand (_16531_, _14383_, _14789_);
  nand (_25062_, _16531_, _16530_);
  nand (_16532_, _14384_, _25063_);
  nand (_16533_, _14792_, _14383_);
  nand (_25064_, _16533_, _16532_);
  nand (_16535_, _14384_, _25065_);
  nand (_16536_, _14795_, _14383_);
  nand (_25066_, _16536_, _16535_);
  nand (_16537_, _14384_, _25067_);
  nand (_16538_, _14799_, _14383_);
  nand (_25068_, _16538_, _16537_);
  nand (_16539_, _14384_, _25069_);
  nand (_16540_, _14802_, _14383_);
  nand (_25070_, _16540_, _16539_);
  nand (_16541_, _14384_, _25071_);
  nand (_16544_, _14805_, _14383_);
  nand (_25072_, _16544_, _16541_);
  nand (_16545_, _14384_, _25073_);
  nand (_16546_, _14808_, _14383_);
  nand (_25074_, _16546_, _16545_);
  nand (_16547_, _14380_, _25075_);
  nand (_16548_, _14379_, _14789_);
  nand (_25076_, _16548_, _16547_);
  nand (_16549_, _14380_, _25077_);
  nand (_16550_, _14792_, _14379_);
  nand (_25078_, _16550_, _16549_);
  nand (_16551_, _14380_, _25079_);
  nand (_16552_, _14795_, _14379_);
  nand (_25080_, _16552_, _16551_);
  nand (_16553_, _14380_, _25081_);
  nand (_16554_, _14799_, _14379_);
  nand (_25082_, _16554_, _16553_);
  nand (_16555_, _14380_, _25083_);
  nand (_16556_, _14802_, _14379_);
  nand (_25084_, _16556_, _16555_);
  nand (_16557_, _14380_, _25085_);
  nand (_16558_, _14805_, _14379_);
  nand (_25086_, _16558_, _16557_);
  nand (_16559_, _14380_, _25087_);
  nand (_16560_, _14808_, _14379_);
  nand (_25088_, _16560_, _16559_);
  nand (_16561_, _14373_, _14789_);
  nand (_16562_, _14375_, _25089_);
  nand (_25090_, _16562_, _16561_);
  nand (_16563_, _14792_, _14373_);
  nand (_16565_, _14375_, _25091_);
  nand (_25092_, _16565_, _16563_);
  nand (_16566_, _14795_, _14373_);
  nand (_16567_, _14375_, _25093_);
  nand (_25094_, _16567_, _16566_);
  nand (_16568_, _14799_, _14373_);
  nand (_16569_, _14375_, _25095_);
  nand (_25096_, _16569_, _16568_);
  nand (_16570_, _14802_, _14373_);
  nand (_16571_, _14375_, _25098_);
  nand (_25099_, _16571_, _16570_);
  nand (_16573_, _14805_, _14373_);
  nand (_16574_, _14375_, _25100_);
  nand (_25101_, _16574_, _16573_);
  nand (_16575_, _14808_, _14373_);
  nand (_16576_, _14375_, _25102_);
  nand (_25103_, _16576_, _16575_);
  nand (_16577_, _14352_, _14789_);
  nand (_16578_, _14354_, _25104_);
  nand (_25105_, _16578_, _16577_);
  nand (_16579_, _14792_, _14352_);
  nand (_16580_, _14354_, _25106_);
  nand (_25107_, _16580_, _16579_);
  nand (_16581_, _14795_, _14352_);
  nand (_16582_, _14354_, _25108_);
  nand (_25109_, _16582_, _16581_);
  nand (_16583_, _14799_, _14352_);
  nand (_16584_, _14354_, _25110_);
  nand (_25111_, _16584_, _16583_);
  nand (_16585_, _14802_, _14352_);
  nand (_16586_, _14354_, _25112_);
  nand (_25113_, _16586_, _16585_);
  nand (_16587_, _14805_, _14352_);
  nand (_16588_, _14354_, _25114_);
  nand (_25115_, _16588_, _16587_);
  nand (_16589_, _14808_, _14352_);
  nand (_16590_, _14354_, _25116_);
  nand (_25117_, _16590_, _16589_);
  nand (_16591_, _14348_, _14789_);
  nand (_16592_, _14350_, _25118_);
  nand (_25119_, _16592_, _16591_);
  nand (_16594_, _14792_, _14348_);
  nand (_16595_, _14350_, _25120_);
  nand (_25121_, _16595_, _16594_);
  nand (_16596_, _14795_, _14348_);
  nand (_16597_, _14350_, _25122_);
  nand (_25123_, _16597_, _16596_);
  nand (_16598_, _14799_, _14348_);
  nand (_16599_, _14350_, _25124_);
  nand (_25125_, _16599_, _16598_);
  nand (_16601_, _14802_, _14348_);
  nand (_16602_, _14350_, _25126_);
  nand (_25127_, _16602_, _16601_);
  nand (_16603_, _14805_, _14348_);
  nand (_16604_, _14350_, _25128_);
  nand (_25129_, _16604_, _16603_);
  nand (_16605_, _14808_, _14348_);
  nand (_16606_, _14350_, _25130_);
  nand (_25131_, _16606_, _16605_);
  nand (_16607_, _14344_, _14789_);
  nand (_16608_, _14346_, _25132_);
  nand (_25133_, _16608_, _16607_);
  nand (_16609_, _14792_, _14344_);
  nand (_16610_, _14346_, _25134_);
  nand (_25135_, _16610_, _16609_);
  nand (_16611_, _14795_, _14344_);
  nand (_16612_, _14346_, _25136_);
  nand (_25137_, _16612_, _16611_);
  nand (_16613_, _14799_, _14344_);
  nand (_16614_, _14346_, _25139_);
  nand (_25140_, _16614_, _16613_);
  nand (_16615_, _14802_, _14344_);
  nand (_16616_, _14346_, _25141_);
  nand (_25142_, _16616_, _16615_);
  nand (_16617_, _14805_, _14344_);
  nand (_16618_, _14346_, _25143_);
  nand (_25144_, _16618_, _16617_);
  nand (_16619_, _14808_, _14344_);
  nand (_16620_, _14346_, _25145_);
  nand (_25146_, _16620_, _16619_);
  nand (_16621_, _14340_, _14789_);
  nand (_16622_, _14342_, _25147_);
  nand (_25148_, _16622_, _16621_);
  nand (_16623_, _14792_, _14340_);
  nand (_16624_, _14342_, _25149_);
  nand (_25150_, _16624_, _16623_);
  nand (_16625_, _14795_, _14340_);
  nand (_16626_, _14342_, _25151_);
  nand (_25152_, _16626_, _16625_);
  nand (_16627_, _14799_, _14340_);
  nand (_16628_, _14342_, _25153_);
  nand (_25154_, _16628_, _16627_);
  nand (_16629_, _14802_, _14340_);
  nand (_16630_, _14342_, _25155_);
  nand (_25156_, _16630_, _16629_);
  nand (_16631_, _14805_, _14340_);
  nand (_16632_, _14342_, _25157_);
  nand (_25158_, _16632_, _16631_);
  nand (_16633_, _14808_, _14340_);
  nand (_16634_, _14342_, _25159_);
  nand (_25160_, _16634_, _16633_);
  nand (_16635_, _14336_, _14789_);
  nand (_16636_, _14338_, _25161_);
  nand (_25162_, _16636_, _16635_);
  nand (_16637_, _14792_, _14336_);
  nand (_16638_, _14338_, _25163_);
  nand (_25164_, _16638_, _16637_);
  nand (_16639_, _14795_, _14336_);
  nand (_16640_, _14338_, _25165_);
  nand (_25166_, _16640_, _16639_);
  nand (_16641_, _14799_, _14336_);
  nand (_16642_, _14338_, _25167_);
  nand (_25168_, _16642_, _16641_);
  nand (_16643_, _14802_, _14336_);
  nand (_16644_, _14338_, _25169_);
  nand (_25170_, _16644_, _16643_);
  nand (_16645_, _14805_, _14336_);
  nand (_16646_, _14338_, _25171_);
  nand (_25172_, _16646_, _16645_);
  nand (_16647_, _14808_, _14336_);
  nand (_16649_, _14338_, _25173_);
  nand (_25174_, _16649_, _16647_);
  nand (_16650_, _14332_, _14789_);
  nand (_16651_, _14334_, _25175_);
  nand (_25176_, _16651_, _16650_);
  nand (_16652_, _14792_, _14332_);
  nand (_16653_, _14334_, _25177_);
  nand (_25178_, _16653_, _16652_);
  nand (_16654_, _14795_, _14332_);
  nand (_16655_, _14334_, _25180_);
  nand (_25181_, _16655_, _16654_);
  nand (_16657_, _14799_, _14332_);
  nand (_16658_, _14334_, _25182_);
  nand (_25183_, _16658_, _16657_);
  nand (_16659_, _14802_, _14332_);
  nand (_16660_, _14334_, _25184_);
  nand (_25185_, _16660_, _16659_);
  nand (_16661_, _14805_, _14332_);
  nand (_16662_, _14334_, _25186_);
  nand (_25187_, _16662_, _16661_);
  nand (_16663_, _14808_, _14332_);
  nand (_16664_, _14334_, _25188_);
  nand (_25189_, _16664_, _16663_);
  nand (_16665_, _14327_, _14789_);
  nand (_16666_, _14329_, _25190_);
  nand (_25191_, _16666_, _16665_);
  nand (_16667_, _14792_, _14327_);
  nand (_16668_, _14329_, _25192_);
  nand (_25193_, _16668_, _16667_);
  nand (_16669_, _14795_, _14327_);
  nand (_16670_, _14329_, _25194_);
  nand (_25195_, _16670_, _16669_);
  nand (_16671_, _14799_, _14327_);
  nand (_16672_, _14329_, _25196_);
  nand (_25197_, _16672_, _16671_);
  nand (_16673_, _14802_, _14327_);
  nand (_16674_, _14329_, _25198_);
  nand (_25199_, _16674_, _16673_);
  nand (_16675_, _14805_, _14327_);
  nand (_16676_, _14329_, _25200_);
  nand (_25201_, _16676_, _16675_);
  nand (_16678_, _14808_, _14327_);
  nand (_16679_, _14329_, _25202_);
  nand (_25203_, _16679_, _16678_);
  nand (_16680_, _14323_, _14789_);
  nand (_16681_, _14325_, _25204_);
  nand (_25205_, _16681_, _16680_);
  nand (_16682_, _14792_, _14323_);
  nand (_16683_, _14325_, _25206_);
  nand (_25207_, _16683_, _16682_);
  nand (_16685_, _14795_, _14323_);
  nand (_16686_, _14325_, _25208_);
  nand (_25209_, _16686_, _16685_);
  nand (_16687_, _14799_, _14323_);
  nand (_16688_, _14325_, _25210_);
  nand (_25211_, _16688_, _16687_);
  nand (_16689_, _14802_, _14323_);
  nand (_16690_, _14325_, _25212_);
  nand (_25213_, _16690_, _16689_);
  nand (_16691_, _14805_, _14323_);
  nand (_16692_, _14325_, _25214_);
  nand (_25215_, _16692_, _16691_);
  nand (_16693_, _14808_, _14323_);
  nand (_16694_, _14325_, _25216_);
  nand (_25217_, _16694_, _16693_);
  nand (_16695_, _14319_, _14789_);
  nand (_16696_, _14321_, _25218_);
  nand (_25219_, _16696_, _16695_);
  nand (_16697_, _14792_, _14319_);
  nand (_16698_, _14321_, _25221_);
  nand (_25222_, _16698_, _16697_);
  nand (_16699_, _14795_, _14319_);
  nand (_16700_, _14321_, _25223_);
  nand (_25224_, _16700_, _16699_);
  nand (_16701_, _14799_, _14319_);
  nand (_16702_, _14321_, _25225_);
  nand (_25226_, _16702_, _16701_);
  nand (_16703_, _14802_, _14319_);
  nand (_16704_, _14321_, _25227_);
  nand (_25228_, _16704_, _16703_);
  nand (_16706_, _14805_, _14319_);
  nand (_16707_, _14321_, _25229_);
  nand (_25230_, _16707_, _16706_);
  nand (_16708_, _14808_, _14319_);
  nand (_16709_, _14321_, _25231_);
  nand (_25232_, _16709_, _16708_);
  nand (_16710_, _14315_, _14789_);
  nand (_16711_, _14317_, _25233_);
  nand (_25234_, _16711_, _16710_);
  nand (_16712_, _14792_, _14315_);
  nand (_16714_, _14317_, _25235_);
  nand (_25236_, _16714_, _16712_);
  nand (_16715_, _14795_, _14315_);
  nand (_16716_, _14317_, _25237_);
  nand (_25238_, _16716_, _16715_);
  nand (_16717_, _14799_, _14315_);
  nand (_16718_, _14317_, _25239_);
  nand (_25240_, _16718_, _16717_);
  nand (_16719_, _14802_, _14315_);
  nand (_16720_, _14317_, _25241_);
  nand (_25242_, _16720_, _16719_);
  nand (_16721_, _14805_, _14315_);
  nand (_16722_, _14317_, _25243_);
  nand (_25244_, _16722_, _16721_);
  nand (_16723_, _14808_, _14315_);
  nand (_16724_, _14317_, _25245_);
  nand (_25246_, _16724_, _16723_);
  nand (_16725_, _14311_, _14789_);
  nand (_16726_, _14313_, _25247_);
  nand (_25248_, _16726_, _16725_);
  nand (_16727_, _14792_, _14311_);
  nand (_16728_, _14313_, _25249_);
  nand (_25250_, _16728_, _16727_);
  nand (_16729_, _14795_, _14311_);
  nand (_16730_, _14313_, _25251_);
  nand (_25252_, _16730_, _16729_);
  nand (_16731_, _14799_, _14311_);
  nand (_16732_, _14313_, _25253_);
  nand (_25254_, _16732_, _16731_);
  nand (_16733_, _14802_, _14311_);
  nand (_16735_, _14313_, _25255_);
  nand (_25256_, _16735_, _16733_);
  nand (_16736_, _14805_, _14311_);
  nand (_16737_, _14313_, _25257_);
  nand (_25258_, _16737_, _16736_);
  nand (_16738_, _14808_, _14311_);
  nand (_16739_, _14313_, _25259_);
  nand (_25260_, _16739_, _16738_);
  nand (_16740_, _14305_, _14789_);
  nand (_16741_, _14307_, _25262_);
  nand (_25263_, _16741_, _16740_);
  nand (_16743_, _14792_, _14305_);
  nand (_16744_, _14307_, _25264_);
  nand (_25265_, _16744_, _16743_);
  nand (_16745_, _14795_, _14305_);
  nand (_16746_, _14307_, _25266_);
  nand (_25267_, _16746_, _16745_);
  nand (_16747_, _14799_, _14305_);
  nand (_16748_, _14307_, _25268_);
  nand (_25269_, _16748_, _16747_);
  nand (_16749_, _14802_, _14305_);
  nand (_16750_, _14307_, _25270_);
  nand (_25271_, _16750_, _16749_);
  nand (_16751_, _14805_, _14305_);
  nand (_16752_, _14307_, _25272_);
  nand (_25273_, _16752_, _16751_);
  nand (_16753_, _14808_, _14305_);
  nand (_16754_, _14307_, _25274_);
  nand (_25275_, _16754_, _16753_);
  nand (_16755_, _14301_, _14789_);
  nand (_16756_, _14303_, _25276_);
  nand (_25277_, _16756_, _16755_);
  nand (_16757_, _14792_, _14301_);
  nand (_16758_, _14303_, _25278_);
  nand (_25279_, _16758_, _16757_);
  nand (_16759_, _14795_, _14301_);
  nand (_16760_, _14303_, _25280_);
  nand (_25281_, _16760_, _16759_);
  nand (_16761_, _14799_, _14301_);
  nand (_16762_, _14303_, _25282_);
  nand (_25283_, _16762_, _16761_);
  nand (_16764_, _14802_, _14301_);
  nand (_16765_, _14303_, _25284_);
  nand (_25285_, _16765_, _16764_);
  nand (_16766_, _14805_, _14301_);
  nand (_16767_, _14303_, _25286_);
  nand (_25287_, _16767_, _16766_);
  nand (_16768_, _14808_, _14301_);
  nand (_16769_, _14303_, _25288_);
  nand (_25289_, _16769_, _16768_);
  nand (_16771_, _14296_, _14789_);
  nand (_16772_, _14299_, _25290_);
  nand (_25291_, _16772_, _16771_);
  nand (_16773_, _14792_, _14296_);
  nand (_16774_, _14299_, _25292_);
  nand (_25293_, _16774_, _16773_);
  nand (_16775_, _14795_, _14296_);
  nand (_16776_, _14299_, _25294_);
  nand (_25295_, _16776_, _16775_);
  nand (_16777_, _14799_, _14296_);
  nand (_16778_, _14299_, _25296_);
  nand (_25297_, _16778_, _16777_);
  nand (_16779_, _14802_, _14296_);
  nand (_16780_, _14299_, _25298_);
  nand (_25299_, _16780_, _16779_);
  nand (_16781_, _14805_, _14296_);
  nand (_16782_, _14299_, _25300_);
  nand (_25301_, _16782_, _16781_);
  nand (_16783_, _14808_, _14296_);
  nand (_16784_, _14299_, _25303_);
  nand (_25304_, _16784_, _16783_);
  nand (_16785_, _14292_, _14789_);
  nand (_16786_, _14294_, _25305_);
  nand (_25306_, _16786_, _16785_);
  nand (_16787_, _14792_, _14292_);
  nand (_16788_, _14294_, _25307_);
  nand (_25308_, _16788_, _16787_);
  nand (_16789_, _14795_, _14292_);
  nand (_16790_, _14294_, _25309_);
  nand (_25310_, _16790_, _16789_);
  nand (_16792_, _14799_, _14292_);
  nand (_16793_, _14294_, _25311_);
  nand (_25312_, _16793_, _16792_);
  nand (_16794_, _14802_, _14292_);
  nand (_16795_, _14294_, _25313_);
  nand (_25314_, _16795_, _16794_);
  nand (_16796_, _14805_, _14292_);
  nand (_16797_, _14294_, _25315_);
  nand (_25316_, _16797_, _16796_);
  nand (_16798_, _14808_, _14292_);
  nand (_16800_, _14294_, _25317_);
  nand (_25318_, _16800_, _16798_);
  nand (_16801_, _14288_, _14789_);
  nand (_16802_, _14290_, _25319_);
  nand (_25320_, _16802_, _16801_);
  nand (_16803_, _14792_, _14288_);
  nand (_16804_, _14290_, _25321_);
  nand (_25322_, _16804_, _16803_);
  nand (_16805_, _14795_, _14288_);
  nand (_16806_, _14290_, _25323_);
  nand (_25324_, _16806_, _16805_);
  nand (_16807_, _14799_, _14288_);
  nand (_16808_, _14290_, _25325_);
  nand (_25326_, _16808_, _16807_);
  nand (_16809_, _14802_, _14288_);
  nand (_16810_, _14290_, _25327_);
  nand (_25328_, _16810_, _16809_);
  nand (_16811_, _14805_, _14288_);
  nand (_16812_, _14290_, _25329_);
  nand (_25330_, _16812_, _16811_);
  nand (_16813_, _14808_, _14288_);
  nand (_16814_, _14290_, _25331_);
  nand (_25332_, _16814_, _16813_);
  nand (_16815_, _14284_, _14789_);
  nand (_16816_, _14286_, _25333_);
  nand (_25334_, _16816_, _16815_);
  nand (_16817_, _14792_, _14284_);
  nand (_16818_, _14286_, _25335_);
  nand (_25336_, _16818_, _16817_);
  nand (_16819_, _14795_, _14284_);
  nand (_16821_, _14286_, _25337_);
  nand (_25338_, _16821_, _16819_);
  nand (_16822_, _14799_, _14284_);
  nand (_16823_, _14286_, _25339_);
  nand (_25340_, _16823_, _16822_);
  nand (_16824_, _14802_, _14284_);
  nand (_16825_, _14286_, _25341_);
  nand (_25342_, _16825_, _16824_);
  nand (_16826_, _14805_, _14284_);
  nand (_16827_, _14286_, _25345_);
  nand (_25346_, _16827_, _16826_);
  nand (_16830_, _14808_, _14284_);
  nand (_16831_, _14286_, _25347_);
  nand (_25348_, _16831_, _16830_);
  nand (_16832_, _14280_, _14789_);
  nand (_16833_, _14282_, _25349_);
  nand (_25350_, _16833_, _16832_);
  nand (_16834_, _14792_, _14280_);
  nand (_16835_, _14282_, _25351_);
  nand (_25352_, _16835_, _16834_);
  nand (_16836_, _14795_, _14280_);
  nand (_16837_, _14282_, _25353_);
  nand (_25354_, _16837_, _16836_);
  nand (_16838_, _14799_, _14280_);
  nand (_16839_, _14282_, _25355_);
  nand (_25356_, _16839_, _16838_);
  nand (_16840_, _14802_, _14280_);
  nand (_16841_, _14282_, _25357_);
  nand (_25358_, _16841_, _16840_);
  nand (_16842_, _14805_, _14280_);
  nand (_16843_, _14282_, _25359_);
  nand (_25360_, _16843_, _16842_);
  nand (_16844_, _14808_, _14280_);
  nand (_16845_, _14282_, _25361_);
  nand (_25362_, _16845_, _16844_);
  nand (_16846_, _14276_, _14789_);
  nand (_16847_, _14278_, _25363_);
  nand (_25364_, _16847_, _16846_);
  nand (_16848_, _14792_, _14276_);
  nand (_16849_, _14278_, _25365_);
  nand (_25366_, _16849_, _16848_);
  nand (_16851_, _14795_, _14276_);
  nand (_16852_, _14278_, _25367_);
  nand (_25368_, _16852_, _16851_);
  nand (_16853_, _14799_, _14276_);
  nand (_16854_, _14278_, _25369_);
  nand (_25370_, _16854_, _16853_);
  nand (_16855_, _14802_, _14276_);
  nand (_16856_, _14278_, _25371_);
  nand (_25372_, _16856_, _16855_);
  nand (_16858_, _14805_, _14276_);
  nand (_16859_, _14278_, _25373_);
  nand (_25374_, _16859_, _16858_);
  nand (_16860_, _14808_, _14276_);
  nand (_16861_, _14278_, _25375_);
  nand (_25376_, _16861_, _16860_);
  nand (_16862_, _14272_, _14789_);
  nand (_16863_, _14274_, _25377_);
  nand (_25378_, _16863_, _16862_);
  nand (_16864_, _14792_, _14272_);
  nand (_16865_, _14274_, _25379_);
  nand (_25380_, _16865_, _16864_);
  nand (_16866_, _14795_, _14272_);
  nand (_16867_, _14274_, _25381_);
  nand (_25382_, _16867_, _16866_);
  nand (_16868_, _14799_, _14272_);
  nand (_16869_, _14274_, _25383_);
  nand (_25384_, _16869_, _16868_);
  nand (_16870_, _14802_, _14272_);
  nand (_16871_, _14274_, _25386_);
  nand (_25387_, _16871_, _16870_);
  nand (_16872_, _14805_, _14272_);
  nand (_16873_, _14274_, _25388_);
  nand (_25389_, _16873_, _16872_);
  nand (_16874_, _14808_, _14272_);
  nand (_16875_, _14274_, _25390_);
  nand (_25391_, _16875_, _16874_);
  nand (_16876_, _14268_, _14789_);
  nand (_16877_, _14270_, _25392_);
  nand (_25393_, _16877_, _16876_);
  nand (_16879_, _14792_, _14268_);
  nand (_16880_, _14270_, _25394_);
  nand (_25395_, _16880_, _16879_);
  nand (_16881_, _14795_, _14268_);
  nand (_16882_, _14270_, _25396_);
  nand (_25397_, _16882_, _16881_);
  nand (_16883_, _14799_, _14268_);
  nand (_16884_, _14270_, _25398_);
  nand (_25399_, _16884_, _16883_);
  nand (_16885_, _14802_, _14268_);
  nand (_16887_, _14270_, _25400_);
  nand (_25401_, _16887_, _16885_);
  nand (_16888_, _14805_, _14268_);
  nand (_16889_, _14270_, _25402_);
  nand (_25403_, _16889_, _16888_);
  nand (_16890_, _14808_, _14268_);
  nand (_16891_, _14270_, _25404_);
  nand (_25405_, _16891_, _16890_);
  nand (_16892_, _14263_, _14789_);
  nand (_16893_, _14266_, _25406_);
  nand (_25407_, _16893_, _16892_);
  nand (_16894_, _14792_, _14263_);
  nand (_16895_, _14266_, _25408_);
  nand (_25409_, _16895_, _16894_);
  nand (_16896_, _14795_, _14263_);
  nand (_16897_, _14266_, _25410_);
  nand (_25411_, _16897_, _16896_);
  nand (_16898_, _14799_, _14263_);
  nand (_16899_, _14266_, _25412_);
  nand (_25413_, _16899_, _16898_);
  nand (_16900_, _14802_, _14263_);
  nand (_16901_, _14266_, _25414_);
  nand (_25415_, _16901_, _16900_);
  nand (_16902_, _14805_, _14263_);
  nand (_16903_, _14266_, _25416_);
  nand (_25417_, _16903_, _16902_);
  nand (_16904_, _14808_, _14263_);
  nand (_16905_, _14266_, _25418_);
  nand (_25419_, _16905_, _16904_);
  nand (_16906_, _14259_, _14789_);
  nand (_16908_, _14261_, _25420_);
  nand (_25421_, _16908_, _16906_);
  nand (_16909_, _14792_, _14259_);
  nand (_16910_, _14261_, _25422_);
  nand (_25423_, _16910_, _16909_);
  nand (_16911_, _14795_, _14259_);
  nand (_16912_, _14261_, _25424_);
  nand (_25425_, _16912_, _16911_);
  nand (_16913_, _14799_, _14259_);
  nand (_16914_, _14261_, _25427_);
  nand (_25428_, _16914_, _16913_);
  nand (_16916_, _14802_, _14259_);
  nand (_16917_, _14261_, _25429_);
  nand (_25430_, _16917_, _16916_);
  nand (_16918_, _14805_, _14259_);
  nand (_16919_, _14261_, _25431_);
  nand (_25432_, _16919_, _16918_);
  nand (_16920_, _14808_, _14259_);
  nand (_16921_, _14261_, _25433_);
  nand (_25434_, _16921_, _16920_);
  nand (_16922_, _14255_, _14789_);
  nand (_16923_, _14257_, _25435_);
  nand (_25436_, _16923_, _16922_);
  nand (_16924_, _14792_, _14255_);
  nand (_16925_, _14257_, _25437_);
  nand (_25438_, _16925_, _16924_);
  nand (_16926_, _14795_, _14255_);
  nand (_16927_, _14257_, _25439_);
  nand (_25440_, _16927_, _16926_);
  nand (_16928_, _14799_, _14255_);
  nand (_16929_, _14257_, _25441_);
  nand (_25442_, _16929_, _16928_);
  nand (_16930_, _14802_, _14255_);
  nand (_16931_, _14257_, _25443_);
  nand (_25444_, _16931_, _16930_);
  nand (_16932_, _14805_, _14255_);
  nand (_16933_, _14257_, _25445_);
  nand (_25446_, _16933_, _16932_);
  nand (_16934_, _14808_, _14255_);
  nand (_16935_, _14257_, _25447_);
  nand (_25448_, _16935_, _16934_);
  nand (_16937_, _14251_, _14789_);
  nand (_16938_, _14253_, _25449_);
  nand (_25450_, _16938_, _16937_);
  nand (_16939_, _14792_, _14251_);
  nand (_16940_, _14253_, _25451_);
  nand (_25452_, _16940_, _16939_);
  nand (_16941_, _14795_, _14251_);
  nand (_16942_, _14253_, _25453_);
  nand (_25454_, _16942_, _16941_);
  nand (_16944_, _14799_, _14251_);
  nand (_16945_, _14253_, _25455_);
  nand (_25456_, _16945_, _16944_);
  nand (_16946_, _14802_, _14251_);
  nand (_16947_, _14253_, _25457_);
  nand (_25458_, _16947_, _16946_);
  nand (_16948_, _14805_, _14251_);
  nand (_16949_, _14253_, _25459_);
  nand (_25460_, _16949_, _16948_);
  nand (_16950_, _14808_, _14251_);
  nand (_16951_, _14253_, _25461_);
  nand (_25462_, _16951_, _16950_);
  nand (_16952_, _14247_, _14789_);
  nand (_16953_, _14249_, _25463_);
  nand (_25464_, _16953_, _16952_);
  nand (_16954_, _14792_, _14247_);
  nand (_16955_, _14249_, _25465_);
  nand (_25466_, _16955_, _16954_);
  nand (_16956_, _14795_, _14247_);
  nand (_16957_, _14249_, _25468_);
  nand (_25469_, _16957_, _16956_);
  nand (_16958_, _14799_, _14247_);
  nand (_16959_, _14249_, _25470_);
  nand (_25471_, _16959_, _16958_);
  nand (_16960_, _14802_, _14247_);
  nand (_16961_, _14249_, _25472_);
  nand (_25473_, _16961_, _16960_);
  nand (_16962_, _14805_, _14247_);
  nand (_16963_, _14249_, _25474_);
  nand (_25475_, _16963_, _16962_);
  nand (_16965_, _14808_, _14247_);
  nand (_16966_, _14249_, _25476_);
  nand (_25477_, _16966_, _16965_);
  nand (_16967_, _14243_, _14789_);
  nand (_16968_, _14245_, _25478_);
  nand (_25479_, _16968_, _16967_);
  nand (_16969_, _14792_, _14243_);
  nand (_16970_, _14245_, _25480_);
  nand (_25481_, _16970_, _16969_);
  nand (_16971_, _14795_, _14243_);
  nand (_16973_, _14245_, _25482_);
  nand (_25483_, _16973_, _16971_);
  nand (_16974_, _14799_, _14243_);
  nand (_16975_, _14245_, _25484_);
  nand (_25485_, _16975_, _16974_);
  nand (_16976_, _14802_, _14243_);
  nand (_16977_, _14245_, _25486_);
  nand (_25487_, _16977_, _16976_);
  nand (_16978_, _14805_, _14243_);
  nand (_16979_, _14245_, _25488_);
  nand (_25489_, _16979_, _16978_);
  nand (_16980_, _14808_, _14243_);
  nand (_16981_, _14245_, _25490_);
  nand (_25491_, _16981_, _16980_);
  nand (_16982_, _14235_, _14789_);
  nand (_16983_, _14237_, _25492_);
  nand (_25493_, _16983_, _16982_);
  nand (_16984_, _14792_, _14235_);
  nand (_16985_, _14237_, _25494_);
  nand (_25495_, _16985_, _16984_);
  nand (_16986_, _14795_, _14235_);
  nand (_16987_, _14237_, _25496_);
  nand (_25497_, _16987_, _16986_);
  nand (_16988_, _14799_, _14235_);
  nand (_16989_, _14237_, _25498_);
  nand (_25499_, _16989_, _16988_);
  nand (_16990_, _14802_, _14235_);
  nand (_16991_, _14237_, _25500_);
  nand (_25501_, _16991_, _16990_);
  nand (_16992_, _14805_, _14235_);
  nand (_16994_, _14237_, _25502_);
  nand (_25503_, _16994_, _16992_);
  nand (_16995_, _14808_, _14235_);
  nand (_16996_, _14237_, _25504_);
  nand (_25505_, _16996_, _16995_);
  nand (_16997_, _14230_, _14789_);
  nand (_16998_, _14233_, _25506_);
  nand (_25507_, _16998_, _16997_);
  nand (_16999_, _14792_, _14230_);
  nand (_17000_, _14233_, _25509_);
  nand (_25510_, _17000_, _16999_);
  nand (_17002_, _14795_, _14230_);
  nand (_17003_, _14233_, _25511_);
  nand (_25512_, _17003_, _17002_);
  nand (_17004_, _14799_, _14230_);
  nand (_17005_, _14233_, _25513_);
  nand (_25514_, _17005_, _17004_);
  nand (_17006_, _14802_, _14230_);
  nand (_17007_, _14233_, _25515_);
  nand (_25516_, _17007_, _17006_);
  nand (_17008_, _14805_, _14230_);
  nand (_17009_, _14233_, _25517_);
  nand (_25518_, _17009_, _17008_);
  nand (_17010_, _14808_, _14230_);
  nand (_17011_, _14233_, _25519_);
  nand (_25520_, _17011_, _17010_);
  nand (_17012_, _14226_, _14789_);
  nand (_17013_, _14228_, _25521_);
  nand (_25522_, _17013_, _17012_);
  nand (_17014_, _14792_, _14226_);
  nand (_17015_, _14228_, _25523_);
  nand (_25524_, _17015_, _17014_);
  nand (_17016_, _14795_, _14226_);
  nand (_17017_, _14228_, _25525_);
  nand (_25526_, _17017_, _17016_);
  nand (_17018_, _14799_, _14226_);
  nand (_17019_, _14228_, _25527_);
  nand (_25528_, _17019_, _17018_);
  nand (_17020_, _14802_, _14226_);
  nand (_17021_, _14228_, _25529_);
  nand (_25530_, _17021_, _17020_);
  nand (_17023_, _14805_, _14226_);
  nand (_17024_, _14228_, _25531_);
  nand (_25532_, _17024_, _17023_);
  nand (_17025_, _14808_, _14226_);
  nand (_17026_, _14228_, _25533_);
  nand (_25534_, _17026_, _17025_);
  nand (_17027_, _14222_, _14789_);
  nand (_17028_, _14224_, _25535_);
  nand (_25536_, _17028_, _17027_);
  nand (_17030_, _14792_, _14222_);
  nand (_17031_, _14224_, _25537_);
  nand (_25538_, _17031_, _17030_);
  nand (_17032_, _14795_, _14222_);
  nand (_17033_, _14224_, _25539_);
  nand (_25540_, _17033_, _17032_);
  nand (_17034_, _14799_, _14222_);
  nand (_17035_, _14224_, _25541_);
  nand (_25542_, _17035_, _17034_);
  nand (_17036_, _14802_, _14222_);
  nand (_17037_, _14224_, _25543_);
  nand (_25544_, _17037_, _17036_);
  nand (_17038_, _14805_, _14222_);
  nand (_17039_, _14224_, _25545_);
  nand (_25546_, _17039_, _17038_);
  nand (_17040_, _14808_, _14222_);
  nand (_17041_, _14224_, _25547_);
  nand (_25548_, _17041_, _17040_);
  nand (_17042_, _14218_, _14789_);
  nand (_17043_, _14220_, _25550_);
  nand (_25551_, _17043_, _17042_);
  nand (_17044_, _14792_, _14218_);
  nand (_17045_, _14220_, _25552_);
  nand (_25553_, _17045_, _17044_);
  nand (_17046_, _14795_, _14218_);
  nand (_17047_, _14220_, _25554_);
  nand (_25555_, _17047_, _17046_);
  nand (_17048_, _14799_, _14218_);
  nand (_17049_, _14220_, _25556_);
  nand (_25557_, _17049_, _17048_);
  nand (_17051_, _14802_, _14218_);
  nand (_17052_, _14220_, _25558_);
  nand (_25559_, _17052_, _17051_);
  nand (_17053_, _14805_, _14218_);
  nand (_17054_, _14220_, _25560_);
  nand (_25561_, _17054_, _17053_);
  nand (_17055_, _14808_, _14218_);
  nand (_17056_, _14220_, _25562_);
  nand (_25563_, _17056_, _17055_);
  nand (_17057_, _14214_, _14789_);
  nand (_17059_, _14216_, _25564_);
  nand (_25565_, _17059_, _17057_);
  nand (_17060_, _14792_, _14214_);
  nand (_17061_, _14216_, _25566_);
  nand (_25567_, _17061_, _17060_);
  nand (_17062_, _14795_, _14214_);
  nand (_17063_, _14216_, _25568_);
  nand (_25569_, _17063_, _17062_);
  nand (_17064_, _14799_, _14214_);
  nand (_17065_, _14216_, _25570_);
  nand (_25571_, _17065_, _17064_);
  nand (_17066_, _14802_, _14214_);
  nand (_17067_, _14216_, _25572_);
  nand (_25573_, _17067_, _17066_);
  nand (_17068_, _14805_, _14214_);
  nand (_17069_, _14216_, _25574_);
  nand (_25575_, _17069_, _17068_);
  nand (_17070_, _14808_, _14214_);
  nand (_17071_, _14216_, _25576_);
  nand (_25577_, _17071_, _17070_);
  nand (_17072_, _14210_, _14789_);
  nand (_17073_, _14212_, _25578_);
  nand (_25579_, _17073_, _17072_);
  nand (_17074_, _14792_, _14210_);
  nand (_17075_, _14212_, _25580_);
  nand (_25581_, _17075_, _17074_);
  nand (_17076_, _14795_, _14210_);
  nand (_17077_, _14212_, _25582_);
  nand (_25583_, _17077_, _17076_);
  nand (_17078_, _14799_, _14210_);
  nand (_17080_, _14212_, _25584_);
  nand (_25585_, _17080_, _17078_);
  nand (_17081_, _14802_, _14210_);
  nand (_17082_, _14212_, _25586_);
  nand (_25587_, _17082_, _17081_);
  nand (_17083_, _14805_, _14210_);
  nand (_17084_, _14212_, _25589_);
  nand (_25591_, _17084_, _17083_);
  nand (_17085_, _14808_, _14210_);
  nand (_17086_, _14212_, _25594_);
  nand (_25596_, _17086_, _17085_);
  nand (_17088_, _14205_, _14789_);
  nand (_17089_, _14208_, _25598_);
  nand (_25600_, _17089_, _17088_);
  nand (_17090_, _14792_, _14205_);
  nand (_17091_, _14208_, _25602_);
  nand (_25604_, _17091_, _17090_);
  nand (_17092_, _14795_, _14205_);
  nand (_17093_, _14208_, _25606_);
  nand (_25608_, _17093_, _17092_);
  nand (_17094_, _14799_, _14205_);
  nand (_17095_, _14208_, _25610_);
  nand (_25612_, _17095_, _17094_);
  nand (_17096_, _14802_, _14205_);
  nand (_17097_, _14208_, _25614_);
  nand (_25616_, _17097_, _17096_);
  nand (_17098_, _14805_, _14205_);
  nand (_17099_, _14208_, _25618_);
  nand (_25620_, _17099_, _17098_);
  nand (_17100_, _14808_, _14205_);
  nand (_17101_, _14208_, _25622_);
  nand (_25624_, _17101_, _17100_);
  nand (_17102_, _14201_, _14789_);
  nand (_17103_, _14203_, _25626_);
  nand (_25628_, _17103_, _17102_);
  nand (_17104_, _14792_, _14201_);
  nand (_17105_, _14203_, _25630_);
  nand (_25632_, _17105_, _17104_);
  nand (_17106_, _14795_, _14201_);
  nand (_17107_, _14203_, _25634_);
  nand (_25636_, _17107_, _17106_);
  nand (_17108_, _14799_, _14201_);
  nand (_17109_, _14203_, _25638_);
  nand (_25640_, _17109_, _17108_);
  nand (_17110_, _14802_, _14201_);
  nand (_17111_, _14203_, _25642_);
  nand (_25644_, _17111_, _17110_);
  nand (_17112_, _14805_, _14201_);
  nand (_17113_, _14203_, _25646_);
  nand (_25648_, _17113_, _17112_);
  nand (_17115_, _14808_, _14201_);
  nand (_17116_, _14203_, _25650_);
  nand (_25652_, _17116_, _17115_);
  nand (_17117_, _14196_, _14789_);
  nand (_17118_, _14199_, _25654_);
  nand (_25656_, _17118_, _17117_);
  nand (_17119_, _14792_, _14196_);
  nand (_17120_, _14199_, _25658_);
  nand (_25660_, _17120_, _17119_);
  nand (_17121_, _14795_, _14196_);
  nand (_17123_, _14199_, _25662_);
  nand (_25664_, _17123_, _17121_);
  nand (_17124_, _14799_, _14196_);
  nand (_17125_, _14199_, _25666_);
  nand (_25668_, _17125_, _17124_);
  nand (_17126_, _14802_, _14196_);
  nand (_17127_, _14199_, _25670_);
  nand (_25672_, _17127_, _17126_);
  nand (_17128_, _14805_, _14196_);
  nand (_17129_, _14199_, _25675_);
  nand (_25677_, _17129_, _17128_);
  nand (_17131_, _14808_, _14196_);
  nand (_17132_, _14199_, _25679_);
  nand (_25681_, _17132_, _17131_);
  nand (_17133_, _14192_, _14789_);
  nand (_17134_, _14194_, _25683_);
  nand (_25685_, _17134_, _17133_);
  nand (_17135_, _14792_, _14192_);
  nand (_17136_, _14194_, _25687_);
  nand (_25689_, _17136_, _17135_);
  nand (_17137_, _14795_, _14192_);
  nand (_17138_, _14194_, _25691_);
  nand (_25693_, _17138_, _17137_);
  nand (_17139_, _14799_, _14192_);
  nand (_17140_, _14194_, _25695_);
  nand (_25697_, _17140_, _17139_);
  nand (_17141_, _14802_, _14192_);
  nand (_17142_, _14194_, _25699_);
  nand (_25701_, _17142_, _17141_);
  nand (_17143_, _14805_, _14192_);
  nand (_17144_, _14194_, _25703_);
  nand (_25705_, _17144_, _17143_);
  nand (_17145_, _14808_, _14192_);
  nand (_17146_, _14194_, _25707_);
  nand (_25709_, _17146_, _17145_);
  nand (_17147_, _14188_, _14789_);
  nand (_17148_, _14190_, _25711_);
  nand (_25713_, _17148_, _17147_);
  nand (_17149_, _14792_, _14188_);
  nand (_17150_, _14190_, _25715_);
  nand (_25717_, _17150_, _17149_);
  nand (_17152_, _14795_, _14188_);
  nand (_17153_, _14190_, _25719_);
  nand (_25721_, _17153_, _17152_);
  nand (_17154_, _14799_, _14188_);
  nand (_17155_, _14190_, _25723_);
  nand (_25725_, _17155_, _17154_);
  nand (_17156_, _14802_, _14188_);
  nand (_17157_, _14190_, _25727_);
  nand (_25729_, _17157_, _17156_);
  nand (_17159_, _14805_, _14188_);
  nand (_17160_, _14190_, _25731_);
  nand (_25733_, _17160_, _17159_);
  nand (_17161_, _14808_, _14188_);
  nand (_17162_, _14190_, _25735_);
  nand (_25737_, _17162_, _17161_);
  nand (_17163_, _14184_, _14789_);
  nand (_17164_, _14186_, _25739_);
  nand (_25741_, _17164_, _17163_);
  nand (_17165_, _14792_, _14184_);
  nand (_17166_, _14186_, _25743_);
  nand (_25745_, _17166_, _17165_);
  nand (_17167_, _14795_, _14184_);
  nand (_17168_, _14186_, _25747_);
  nand (_25749_, _17168_, _17167_);
  nand (_17169_, _14799_, _14184_);
  nand (_17170_, _14186_, _25751_);
  nand (_25753_, _17170_, _17169_);
  nand (_17171_, _14802_, _14184_);
  nand (_17172_, _14186_, _25756_);
  nand (_25758_, _17172_, _17171_);
  nand (_17173_, _14805_, _14184_);
  nand (_17174_, _14186_, _25760_);
  nand (_25762_, _17174_, _17173_);
  nand (_17175_, _14808_, _14184_);
  nand (_17176_, _14186_, _25764_);
  nand (_25766_, _17176_, _17175_);
  nand (_17177_, _14180_, _14789_);
  nand (_17178_, _14182_, _25768_);
  nand (_25770_, _17178_, _17177_);
  nand (_17180_, _14792_, _14180_);
  nand (_17181_, _14182_, _25772_);
  nand (_25774_, _17181_, _17180_);
  nand (_17182_, _14795_, _14180_);
  nand (_17183_, _14182_, _25776_);
  nand (_25778_, _17183_, _17182_);
  nand (_17184_, _14799_, _14180_);
  nand (_17185_, _14182_, _25780_);
  nand (_25782_, _17185_, _17184_);
  nand (_17186_, _14802_, _14180_);
  nand (_17188_, _14182_, _25784_);
  nand (_25786_, _17188_, _17186_);
  nand (_17189_, _14805_, _14180_);
  nand (_17190_, _14182_, _25788_);
  nand (_25790_, _17190_, _17189_);
  nand (_17191_, _14808_, _14180_);
  nand (_17192_, _14182_, _25792_);
  nand (_25794_, _17192_, _17191_);
  nand (_17193_, _14176_, _14789_);
  nand (_17194_, _14178_, _25796_);
  nand (_25798_, _17194_, _17193_);
  nand (_17195_, _14792_, _14176_);
  nand (_17196_, _14178_, _25800_);
  nand (_25802_, _17196_, _17195_);
  nand (_17197_, _14795_, _14176_);
  nand (_17198_, _14178_, _25804_);
  nand (_25806_, _17198_, _17197_);
  nand (_17199_, _14799_, _14176_);
  nand (_17200_, _14178_, _25808_);
  nand (_25810_, _17200_, _17199_);
  nand (_17201_, _14802_, _14176_);
  nand (_17202_, _14178_, _25812_);
  nand (_25814_, _17202_, _17201_);
  nand (_17203_, _14805_, _14176_);
  nand (_17204_, _14178_, _25816_);
  nand (_25818_, _17204_, _17203_);
  nand (_17205_, _14808_, _14176_);
  nand (_17206_, _14178_, _25820_);
  nand (_25822_, _17206_, _17205_);
  nand (_17207_, _14172_, _14789_);
  nand (_17209_, _14174_, _25824_);
  nand (_25826_, _17209_, _17207_);
  nand (_17210_, _14792_, _14172_);
  nand (_17211_, _14174_, _25828_);
  nand (_25830_, _17211_, _17210_);
  nand (_17212_, _14795_, _14172_);
  nand (_17213_, _14174_, _25832_);
  nand (_25834_, _17213_, _17212_);
  nand (_17214_, _14799_, _14172_);
  nand (_17215_, _14174_, _25837_);
  nand (_25839_, _17215_, _17214_);
  nand (_17217_, _14802_, _14172_);
  nand (_17218_, _14174_, _25841_);
  nand (_25843_, _17218_, _17217_);
  nand (_17219_, _14805_, _14172_);
  nand (_17220_, _14174_, _25845_);
  nand (_25847_, _17220_, _17219_);
  nand (_17221_, _14808_, _14172_);
  nand (_17222_, _14174_, _25849_);
  nand (_25851_, _17222_, _17221_);
  nand (_17223_, _14166_, _14789_);
  nand (_17224_, _14168_, _25853_);
  nand (_25855_, _17224_, _17223_);
  nand (_17225_, _14792_, _14166_);
  nand (_17226_, _14168_, _25857_);
  nand (_25859_, _17226_, _17225_);
  nand (_17227_, _14795_, _14166_);
  nand (_17228_, _14168_, _25861_);
  nand (_25863_, _17228_, _17227_);
  nand (_17229_, _14799_, _14166_);
  nand (_17230_, _14168_, _25865_);
  nand (_25867_, _17230_, _17229_);
  nand (_17231_, _14802_, _14166_);
  nand (_17232_, _14168_, _25869_);
  nand (_25871_, _17232_, _17231_);
  nand (_17233_, _14805_, _14166_);
  nand (_17234_, _14168_, _25873_);
  nand (_25875_, _17234_, _17233_);
  nand (_17235_, _14808_, _14166_);
  nand (_17236_, _14168_, _25877_);
  nand (_25879_, _17236_, _17235_);
  nand (_17238_, _14161_, _14789_);
  nand (_17239_, _14163_, _25881_);
  nand (_25883_, _17239_, _17238_);
  nand (_17240_, _14792_, _14161_);
  nand (_17241_, _14163_, _25885_);
  nand (_25887_, _17241_, _17240_);
  nand (_17242_, _14795_, _14161_);
  nand (_17243_, _14163_, _25889_);
  nand (_25891_, _17243_, _17242_);
  nand (_17245_, _14799_, _14161_);
  nand (_17246_, _14163_, _25893_);
  nand (_25895_, _17246_, _17245_);
  nand (_17247_, _14802_, _14161_);
  nand (_17248_, _14163_, _25897_);
  nand (_25899_, _17248_, _17247_);
  nand (_17249_, _14805_, _14161_);
  nand (_17250_, _14163_, _25901_);
  nand (_25903_, _17250_, _17249_);
  nand (_17251_, _14808_, _14161_);
  nand (_17252_, _14163_, _25905_);
  nand (_25907_, _17252_, _17251_);
  nand (_17253_, _14157_, _14789_);
  nand (_17254_, _14159_, _25909_);
  nand (_25911_, _17254_, _17253_);
  nand (_17255_, _14792_, _14157_);
  nand (_17256_, _14159_, _25913_);
  nand (_25915_, _17256_, _17255_);
  nand (_17257_, _14795_, _14157_);
  nand (_17258_, _14159_, _25919_);
  nand (_25921_, _17258_, _17257_);
  nand (_17259_, _14799_, _14157_);
  nand (_17260_, _14159_, _25923_);
  nand (_25925_, _17260_, _17259_);
  nand (_17261_, _14802_, _14157_);
  nand (_17262_, _14159_, _25927_);
  nand (_25929_, _17262_, _17261_);
  nand (_17263_, _14805_, _14157_);
  nand (_17264_, _14159_, _25931_);
  nand (_25933_, _17264_, _17263_);
  nand (_17266_, _14808_, _14157_);
  nand (_17267_, _14159_, _25935_);
  nand (_25937_, _17267_, _17266_);
  nand (_17268_, _14153_, _14789_);
  nand (_17269_, _14155_, _25939_);
  nand (_25941_, _17269_, _17268_);
  nand (_17270_, _14792_, _14153_);
  nand (_17271_, _14155_, _25943_);
  nand (_25945_, _17271_, _17270_);
  nand (_17272_, _14795_, _14153_);
  nand (_17274_, _14155_, _25947_);
  nand (_25949_, _17274_, _17272_);
  nand (_17275_, _14799_, _14153_);
  nand (_17276_, _14155_, _25951_);
  nand (_25953_, _17276_, _17275_);
  nand (_17277_, _14802_, _14153_);
  nand (_17278_, _14155_, _25955_);
  nand (_25957_, _17278_, _17277_);
  nand (_17279_, _14805_, _14153_);
  nand (_17280_, _14155_, _25959_);
  nand (_25961_, _17280_, _17279_);
  nand (_17281_, _14808_, _14153_);
  nand (_17282_, _14155_, _25963_);
  nand (_25965_, _17282_, _17281_);
  nand (_17283_, _14149_, _14789_);
  nand (_17284_, _14151_, _25967_);
  nand (_25969_, _17284_, _17283_);
  nand (_17285_, _14792_, _14149_);
  nand (_17286_, _14151_, _25971_);
  nand (_25973_, _17286_, _17285_);
  nand (_17287_, _14795_, _14149_);
  nand (_17288_, _14151_, _25975_);
  nand (_25977_, _17288_, _17287_);
  nand (_17289_, _14799_, _14149_);
  nand (_17290_, _14151_, _25979_);
  nand (_25981_, _17290_, _17289_);
  nand (_17291_, _14802_, _14149_);
  nand (_17292_, _14151_, _25983_);
  nand (_25985_, _17292_, _17291_);
  nand (_17293_, _14805_, _14149_);
  nand (_17295_, _14151_, _25987_);
  nand (_25989_, _17295_, _17293_);
  nand (_17296_, _14808_, _14149_);
  nand (_17297_, _14151_, _25991_);
  nand (_25993_, _17297_, _17296_);
  nand (_17298_, _14145_, _14789_);
  nand (_17299_, _14147_, _25995_);
  nand (_25997_, _17299_, _17298_);
  nand (_17300_, _14792_, _14145_);
  nand (_17301_, _14147_, _26000_);
  nand (_26002_, _17301_, _17300_);
  nand (_17303_, _14795_, _14145_);
  nand (_17304_, _14147_, _26004_);
  nand (_26006_, _17304_, _17303_);
  nand (_17305_, _14799_, _14145_);
  nand (_17306_, _14147_, _26008_);
  nand (_26010_, _17306_, _17305_);
  nand (_17307_, _14802_, _14145_);
  nand (_17308_, _14147_, _26012_);
  nand (_26014_, _17308_, _17307_);
  nand (_17309_, _14805_, _14145_);
  nand (_17310_, _14147_, _26016_);
  nand (_26018_, _17310_, _17309_);
  nand (_17311_, _14808_, _14145_);
  nand (_17312_, _14147_, _26020_);
  nand (_26022_, _17312_, _17311_);
  nand (_17313_, _14141_, _14789_);
  nand (_17314_, _14143_, _26024_);
  nand (_26026_, _17314_, _17313_);
  nand (_17315_, _14792_, _14141_);
  nand (_17316_, _14143_, _26028_);
  nand (_26030_, _17316_, _17315_);
  nand (_17317_, _14795_, _14141_);
  nand (_17318_, _14143_, _26032_);
  nand (_26034_, _17318_, _17317_);
  nand (_17319_, _14799_, _14141_);
  nand (_17320_, _14143_, _26036_);
  nand (_26038_, _17320_, _17319_);
  nand (_17321_, _14802_, _14141_);
  nand (_17322_, _14143_, _26040_);
  nand (_26042_, _17322_, _17321_);
  nand (_17324_, _14805_, _14141_);
  nand (_17325_, _14143_, _26044_);
  nand (_26046_, _17325_, _17324_);
  nand (_17326_, _14808_, _14141_);
  nand (_17327_, _14143_, _26048_);
  nand (_26050_, _17327_, _17326_);
  nand (_17328_, _14137_, _14789_);
  nand (_17329_, _14139_, _26052_);
  nand (_26054_, _17329_, _17328_);
  nand (_17331_, _14792_, _14137_);
  nand (_17332_, _14139_, _26056_);
  nand (_26058_, _17332_, _17331_);
  nand (_17333_, _14795_, _14137_);
  nand (_17334_, _14139_, _26060_);
  nand (_26062_, _17334_, _17333_);
  nand (_17335_, _14799_, _14137_);
  nand (_17336_, _14139_, _26064_);
  nand (_26066_, _17336_, _17335_);
  nand (_17337_, _14802_, _14137_);
  nand (_17338_, _14139_, _26068_);
  nand (_26070_, _17338_, _17337_);
  nand (_17339_, _14805_, _14137_);
  nand (_17340_, _14139_, _26072_);
  nand (_26074_, _17340_, _17339_);
  nand (_17341_, _14808_, _14137_);
  nand (_17342_, _14139_, _26076_);
  nand (_26078_, _17342_, _17341_);
  nand (_17343_, _14133_, _14789_);
  nand (_17344_, _14135_, _26081_);
  nand (_26083_, _17344_, _17343_);
  nand (_17345_, _14792_, _14133_);
  nand (_17346_, _14135_, _26085_);
  nand (_26087_, _17346_, _17345_);
  nand (_17347_, _14795_, _14133_);
  nand (_17348_, _14135_, _26089_);
  nand (_26091_, _17348_, _17347_);
  nand (_17349_, _14799_, _14133_);
  nand (_17350_, _14135_, _26093_);
  nand (_26095_, _17350_, _17349_);
  nand (_17352_, _14802_, _14133_);
  nand (_17353_, _14135_, _26097_);
  nand (_26099_, _17353_, _17352_);
  nand (_17354_, _14805_, _14133_);
  nand (_17355_, _14135_, _26101_);
  nand (_26103_, _17355_, _17354_);
  nand (_17356_, _14808_, _14133_);
  nand (_17357_, _14135_, _26105_);
  nand (_26107_, _17357_, _17356_);
  nand (_17358_, _14128_, _14789_);
  nand (_17360_, _14130_, _26109_);
  nand (_26111_, _17360_, _17358_);
  nand (_17361_, _14792_, _14128_);
  nand (_17362_, _14130_, _26113_);
  nand (_26115_, _17362_, _17361_);
  nand (_17363_, _14795_, _14128_);
  nand (_17364_, _14130_, _26117_);
  nand (_26119_, _17364_, _17363_);
  nand (_17365_, _14799_, _14128_);
  nand (_17366_, _14130_, _26121_);
  nand (_26123_, _17366_, _17365_);
  nand (_17367_, _14802_, _14128_);
  nand (_17368_, _14130_, _26125_);
  nand (_26127_, _17368_, _17367_);
  nand (_17369_, _14805_, _14128_);
  nand (_17370_, _14130_, _26129_);
  nand (_26131_, _17370_, _17369_);
  nand (_17371_, _14808_, _14128_);
  nand (_17372_, _14130_, _26133_);
  nand (_26135_, _17372_, _17371_);
  nand (_17373_, _14124_, _14789_);
  nand (_17374_, _14126_, _26137_);
  nand (_26139_, _17374_, _17373_);
  nand (_17375_, _14792_, _14124_);
  nand (_17376_, _14126_, _26141_);
  nand (_26143_, _17376_, _17375_);
  nand (_17377_, _14795_, _14124_);
  nand (_17378_, _14126_, _26145_);
  nand (_26147_, _17378_, _17377_);
  nand (_17379_, _14799_, _14124_);
  nand (_17381_, _14126_, _26149_);
  nand (_26151_, _17381_, _17379_);
  nand (_17382_, _14802_, _14124_);
  nand (_17383_, _14126_, _26153_);
  nand (_26155_, _17383_, _17382_);
  nand (_17384_, _14805_, _14124_);
  nand (_17385_, _14126_, _26157_);
  nand (_26159_, _17385_, _17384_);
  nand (_17386_, _14808_, _14124_);
  nand (_17387_, _14126_, _26162_);
  nand (_26164_, _17387_, _17386_);
  nand (_17389_, _14120_, _14789_);
  nand (_17390_, _14122_, _26166_);
  nand (_26168_, _17390_, _17389_);
  nand (_17391_, _14792_, _14120_);
  nand (_17392_, _14122_, _26170_);
  nand (_26172_, _17392_, _17391_);
  nand (_17393_, _14795_, _14120_);
  nand (_17394_, _14122_, _26174_);
  nand (_26176_, _17394_, _17393_);
  nand (_17395_, _14799_, _14120_);
  nand (_17396_, _14122_, _26178_);
  nand (_26180_, _17396_, _17395_);
  nand (_17397_, _14802_, _14120_);
  nand (_17398_, _14122_, _26182_);
  nand (_26184_, _17398_, _17397_);
  nand (_17399_, _14805_, _14120_);
  nand (_17400_, _14122_, _26186_);
  nand (_26188_, _17400_, _17399_);
  nand (_17401_, _14808_, _14120_);
  nand (_17404_, _14122_, _26190_);
  nand (_26192_, _17404_, _17401_);
  nand (_17405_, _14116_, _14789_);
  nand (_17406_, _14118_, _26194_);
  nand (_26196_, _17406_, _17405_);
  nand (_17407_, _14792_, _14116_);
  nand (_17408_, _14118_, _26198_);
  nand (_26200_, _17408_, _17407_);
  nand (_17409_, _14795_, _14116_);
  nand (_17410_, _14118_, _26202_);
  nand (_26204_, _17410_, _17409_);
  nand (_17412_, _14799_, _14116_);
  nand (_17413_, _14118_, _26206_);
  nand (_26208_, _17413_, _17412_);
  nand (_17414_, _14802_, _14116_);
  nand (_17415_, _14118_, _26210_);
  nand (_26212_, _17415_, _17414_);
  nand (_17416_, _14805_, _14116_);
  nand (_17417_, _14118_, _26214_);
  nand (_26216_, _17417_, _17416_);
  nand (_17419_, _14808_, _14116_);
  nand (_17420_, _14118_, _26218_);
  nand (_26220_, _17420_, _17419_);
  nand (_17421_, _14112_, _14789_);
  nand (_17422_, _14114_, _26222_);
  nand (_26224_, _17422_, _17421_);
  nand (_17423_, _14792_, _14112_);
  nand (_17424_, _14114_, _26226_);
  nand (_26228_, _17424_, _17423_);
  nand (_17425_, _14795_, _14112_);
  nand (_17426_, _14114_, _26230_);
  nand (_26232_, _17426_, _17425_);
  nand (_17427_, _14799_, _14112_);
  nand (_17428_, _14114_, _26234_);
  nand (_26236_, _17428_, _17427_);
  nand (_17429_, _14802_, _14112_);
  nand (_17430_, _14114_, _26238_);
  nand (_26240_, _17430_, _17429_);
  nand (_17431_, _14805_, _14112_);
  nand (_17432_, _14114_, _26243_);
  nand (_26245_, _17432_, _17431_);
  nand (_17433_, _14808_, _14112_);
  nand (_17434_, _14114_, _26247_);
  nand (_26249_, _17434_, _17433_);
  nand (_17435_, _14108_, _14789_);
  nand (_17436_, _14110_, _26251_);
  nand (_26253_, _17436_, _17435_);
  nand (_17437_, _14792_, _14108_);
  nand (_17438_, _14110_, _26255_);
  nand (_26257_, _17438_, _17437_);
  nand (_17440_, _14795_, _14108_);
  nand (_17441_, _14110_, _26259_);
  nand (_26261_, _17441_, _17440_);
  nand (_17442_, _14799_, _14108_);
  nand (_17443_, _14110_, _26263_);
  nand (_26265_, _17443_, _17442_);
  nand (_17444_, _14802_, _14108_);
  nand (_17445_, _14110_, _26267_);
  nand (_26269_, _17445_, _17444_);
  nand (_17446_, _14805_, _14108_);
  nand (_17448_, _14110_, _26271_);
  nand (_26273_, _17448_, _17446_);
  nand (_17449_, _14808_, _14108_);
  nand (_17450_, _14110_, _26275_);
  nand (_26277_, _17450_, _17449_);
  nand (_17451_, _14104_, _14789_);
  nand (_17452_, _14106_, _26279_);
  nand (_26281_, _17452_, _17451_);
  nand (_17453_, _14792_, _14104_);
  nand (_17454_, _14106_, _26283_);
  nand (_26285_, _17454_, _17453_);
  nand (_17455_, _14795_, _14104_);
  nand (_17456_, _14106_, _26287_);
  nand (_26289_, _17456_, _17455_);
  nand (_17457_, _14799_, _14104_);
  nand (_17458_, _14106_, _26291_);
  nand (_26293_, _17458_, _17457_);
  nand (_17459_, _14802_, _14104_);
  nand (_17460_, _14106_, _26295_);
  nand (_26297_, _17460_, _17459_);
  nand (_17461_, _14805_, _14104_);
  nand (_17462_, _14106_, _26299_);
  nand (_26301_, _17462_, _17461_);
  nand (_17463_, _14808_, _14104_);
  nand (_17464_, _14106_, _26303_);
  nand (_26305_, _17464_, _17463_);
  nand (_17465_, _14098_, _14789_);
  nand (_17466_, _14100_, _26307_);
  nand (_26309_, _17466_, _17465_);
  nand (_17467_, _14792_, _14098_);
  nand (_17469_, _14100_, _26311_);
  nand (_26313_, _17469_, _17467_);
  nand (_17470_, _14795_, _14098_);
  nand (_17471_, _14100_, _26315_);
  nand (_26317_, _17471_, _17470_);
  nand (_17472_, _14799_, _14098_);
  nand (_17473_, _14100_, _26319_);
  nand (_26321_, _17473_, _17472_);
  nand (_17474_, _14802_, _14098_);
  nand (_17475_, _14100_, _26324_);
  nand (_26326_, _17475_, _17474_);
  nand (_17477_, _14805_, _14098_);
  nand (_17478_, _14100_, _26328_);
  nand (_26330_, _17478_, _17477_);
  nand (_17479_, _14808_, _14098_);
  nand (_17480_, _14100_, _26332_);
  nand (_26334_, _17480_, _17479_);
  nand (_17481_, _14093_, _14789_);
  nand (_17482_, _14095_, _26336_);
  nand (_26338_, _17482_, _17481_);
  nand (_17483_, _14792_, _14093_);
  nand (_17484_, _14095_, _26340_);
  nand (_26342_, _17484_, _17483_);
  nand (_17485_, _14795_, _14093_);
  nand (_17486_, _14095_, _26344_);
  nand (_26346_, _17486_, _17485_);
  nand (_17487_, _14799_, _14093_);
  nand (_17488_, _14095_, _26348_);
  nand (_26350_, _17488_, _17487_);
  nand (_17489_, _14802_, _14093_);
  nand (_17490_, _14095_, _26352_);
  nand (_26354_, _17490_, _17489_);
  nand (_17491_, _14805_, _14093_);
  nand (_17492_, _14095_, _26356_);
  nand (_26358_, _17492_, _17491_);
  nand (_17493_, _14808_, _14093_);
  nand (_17494_, _14095_, _26360_);
  nand (_26362_, _17494_, _17493_);
  nand (_17495_, _14089_, _14789_);
  nand (_17496_, _14091_, _26364_);
  nand (_26366_, _17496_, _17495_);
  nand (_17498_, _14792_, _14089_);
  nand (_17499_, _14091_, _26368_);
  nand (_26370_, _17499_, _17498_);
  nand (_17500_, _14795_, _14089_);
  nand (_17501_, _14091_, _26372_);
  nand (_26374_, _17501_, _17500_);
  nand (_17502_, _14799_, _14089_);
  nand (_17503_, _14091_, _26376_);
  nand (_26378_, _17503_, _17502_);
  nand (_17505_, _14802_, _14089_);
  nand (_17506_, _14091_, _26380_);
  nand (_26382_, _17506_, _17505_);
  nand (_17507_, _14805_, _14089_);
  nand (_17508_, _14091_, _26384_);
  nand (_26386_, _17508_, _17507_);
  nand (_17509_, _14808_, _14089_);
  nand (_17510_, _14091_, _26388_);
  nand (_26390_, _17510_, _17509_);
  nand (_17511_, _14085_, _14789_);
  nand (_17512_, _14087_, _26392_);
  nand (_26394_, _17512_, _17511_);
  nand (_17513_, _14792_, _14085_);
  nand (_17514_, _14087_, _26396_);
  nand (_26398_, _17514_, _17513_);
  nand (_17515_, _14795_, _14085_);
  nand (_17516_, _14087_, _26400_);
  nand (_26402_, _17516_, _17515_);
  nand (_17517_, _14799_, _14085_);
  nand (_17518_, _14087_, _26405_);
  nand (_26407_, _17518_, _17517_);
  nand (_17519_, _14802_, _14085_);
  nand (_17520_, _14087_, _26409_);
  nand (_26411_, _17520_, _17519_);
  nand (_17521_, _14805_, _14085_);
  nand (_17522_, _14087_, _26413_);
  nand (_26415_, _17522_, _17521_);
  nand (_17523_, _14808_, _14085_);
  nand (_17524_, _14087_, _26417_);
  nand (_26419_, _17524_, _17523_);
  nand (_17526_, _14081_, _14789_);
  nand (_17527_, _14083_, _26421_);
  nand (_26423_, _17527_, _17526_);
  nand (_17528_, _14792_, _14081_);
  nand (_17529_, _14083_, _26425_);
  nand (_26427_, _17529_, _17528_);
  nand (_17530_, _14795_, _14081_);
  nand (_17531_, _14083_, _26429_);
  nand (_26431_, _17531_, _17530_);
  nand (_17532_, _14799_, _14081_);
  nand (_17534_, _14083_, _26433_);
  nand (_26435_, _17534_, _17532_);
  nand (_17535_, _14802_, _14081_);
  nand (_17536_, _14083_, _26437_);
  nand (_26439_, _17536_, _17535_);
  nand (_17537_, _14805_, _14081_);
  nand (_17538_, _14083_, _26441_);
  nand (_26443_, _17538_, _17537_);
  nand (_17539_, _14808_, _14081_);
  nand (_17540_, _14083_, _26445_);
  nand (_26447_, _17540_, _17539_);
  nand (_17541_, _14077_, _14789_);
  nand (_17542_, _14079_, _26449_);
  nand (_26451_, _17542_, _17541_);
  nand (_17543_, _14792_, _14077_);
  nand (_17544_, _14079_, _26453_);
  nand (_26455_, _17544_, _17543_);
  nand (_17545_, _14795_, _14077_);
  nand (_17546_, _14079_, _26457_);
  nand (_26459_, _17546_, _17545_);
  nand (_17547_, _14799_, _14077_);
  nand (_17548_, _14079_, _26461_);
  nand (_26463_, _17548_, _17547_);
  nand (_17549_, _14802_, _14077_);
  nand (_17550_, _14079_, _26465_);
  nand (_26467_, _17550_, _17549_);
  nand (_17551_, _14805_, _14077_);
  nand (_17552_, _14079_, _26469_);
  nand (_26471_, _17552_, _17551_);
  nand (_17553_, _14808_, _14077_);
  nand (_17555_, _14079_, _26473_);
  nand (_26475_, _17555_, _17553_);
  nand (_17556_, _14073_, _14789_);
  nand (_17557_, _14075_, _26477_);
  nand (_26479_, _17557_, _17556_);
  nand (_17558_, _14792_, _14073_);
  nand (_17559_, _14075_, _26481_);
  nand (_26483_, _17559_, _17558_);
  nand (_17560_, _14795_, _14073_);
  nand (_17561_, _14075_, _26486_);
  nand (_26488_, _17561_, _17560_);
  nand (_17563_, _14799_, _14073_);
  nand (_17564_, _14075_, _26490_);
  nand (_26492_, _17564_, _17563_);
  nand (_17565_, _14802_, _14073_);
  nand (_17566_, _14075_, _26494_);
  nand (_26496_, _17566_, _17565_);
  nand (_17567_, _14805_, _14073_);
  nand (_17568_, _14075_, _26498_);
  nand (_26500_, _17568_, _17567_);
  nand (_17569_, _14808_, _14073_);
  nand (_17570_, _14075_, _26502_);
  nand (_26504_, _17570_, _17569_);
  nand (_17571_, _14069_, _14789_);
  nand (_17572_, _14071_, _26506_);
  nand (_26508_, _17572_, _17571_);
  nand (_17573_, _14792_, _14069_);
  nand (_17574_, _14071_, _26510_);
  nand (_26512_, _17574_, _17573_);
  nand (_17575_, _14795_, _14069_);
  nand (_17576_, _14071_, _26514_);
  nand (_26516_, _17576_, _17575_);
  nand (_17577_, _14799_, _14069_);
  nand (_17578_, _14071_, _26518_);
  nand (_26520_, _17578_, _17577_);
  nand (_17579_, _14802_, _14069_);
  nand (_17580_, _14071_, _26522_);
  nand (_26524_, _17580_, _17579_);
  nand (_17581_, _14805_, _14069_);
  nand (_17582_, _14071_, _26526_);
  nand (_26528_, _17582_, _17581_);
  nand (_17583_, _14808_, _14069_);
  nand (_17584_, _14071_, _26530_);
  nand (_26532_, _17584_, _17583_);
  nand (_17585_, _14065_, _14789_);
  nand (_17586_, _14067_, _26534_);
  nand (_26536_, _17586_, _17585_);
  nand (_17587_, _14792_, _14065_);
  nand (_17588_, _14067_, _26538_);
  nand (_26540_, _17588_, _17587_);
  nand (_17589_, _14795_, _14065_);
  nand (_17590_, _14067_, _26542_);
  nand (_26544_, _17590_, _17589_);
  nand (_17591_, _14799_, _14065_);
  nand (_17592_, _14067_, _26546_);
  nand (_26548_, _17592_, _17591_);
  nand (_17593_, _14802_, _14065_);
  nand (_17594_, _14067_, _26550_);
  nand (_26552_, _17594_, _17593_);
  nand (_17595_, _14805_, _14065_);
  nand (_17596_, _14067_, _26554_);
  nand (_26556_, _17596_, _17595_);
  nand (_17597_, _14808_, _14065_);
  nand (_17598_, _14067_, _26558_);
  nand (_26560_, _17598_, _17597_);
  nand (_17599_, _14060_, _14789_);
  nand (_17600_, _14062_, _26562_);
  nand (_26564_, _17600_, _17599_);
  nand (_17601_, _14792_, _14060_);
  nand (_17602_, _14062_, _26567_);
  nand (_26569_, _17602_, _17601_);
  nand (_17603_, _14795_, _14060_);
  nand (_17604_, _14062_, _26571_);
  nand (_26573_, _17604_, _17603_);
  nand (_17605_, _14799_, _14060_);
  nand (_17606_, _14062_, _26575_);
  nand (_26577_, _17606_, _17605_);
  nand (_17607_, _14802_, _14060_);
  nand (_17608_, _14062_, _26579_);
  nand (_26581_, _17608_, _17607_);
  nand (_17610_, _14805_, _14060_);
  nand (_17611_, _14062_, _26583_);
  nand (_26585_, _17611_, _17610_);
  nand (_17612_, _14808_, _14060_);
  nand (_17613_, _14062_, _26587_);
  nand (_26589_, _17613_, _17612_);
  nand (_17614_, _14056_, _14789_);
  nand (_17615_, _14058_, _26591_);
  nand (_26593_, _17615_, _17614_);
  nand (_17616_, _14792_, _14056_);
  nand (_17618_, _14058_, _26595_);
  nand (_26597_, _17618_, _17616_);
  nand (_17619_, _14795_, _14056_);
  nand (_17620_, _14058_, _26599_);
  nand (_26601_, _17620_, _17619_);
  nand (_17621_, _14799_, _14056_);
  nand (_17622_, _14058_, _26603_);
  nand (_26605_, _17622_, _17621_);
  nand (_17623_, _14802_, _14056_);
  nand (_17624_, _14058_, _26607_);
  nand (_26609_, _17624_, _17623_);
  nand (_17625_, _14805_, _14056_);
  nand (_17626_, _14058_, _26611_);
  nand (_26613_, _17626_, _17625_);
  nand (_17627_, _14808_, _14056_);
  nand (_17628_, _14058_, _26615_);
  nand (_26617_, _17628_, _17627_);
  nand (_17629_, _14052_, _14789_);
  nand (_17630_, _14054_, _26619_);
  nand (_26621_, _17630_, _17629_);
  nand (_17631_, _14792_, _14052_);
  nand (_17632_, _14054_, _26623_);
  nand (_26625_, _17632_, _17631_);
  nand (_17633_, _14795_, _14052_);
  nand (_17634_, _14054_, _26627_);
  nand (_26629_, _17634_, _17633_);
  nand (_17635_, _14799_, _14052_);
  nand (_17636_, _14054_, _26631_);
  nand (_26633_, _17636_, _17635_);
  nand (_17637_, _14802_, _14052_);
  nand (_17639_, _14054_, _26635_);
  nand (_26637_, _17639_, _17637_);
  nand (_17640_, _14805_, _14052_);
  nand (_17641_, _14054_, _26639_);
  nand (_26641_, _17641_, _17640_);
  nand (_17642_, _14808_, _14052_);
  nand (_17643_, _14054_, _26643_);
  nand (_26645_, _17643_, _17642_);
  nand (_17644_, _14048_, _14789_);
  nand (_17645_, _14050_, _26648_);
  nand (_26650_, _17645_, _17644_);
  nand (_17647_, _14792_, _14048_);
  nand (_17648_, _14050_, _26652_);
  nand (_26654_, _17648_, _17647_);
  nand (_17649_, _14795_, _14048_);
  nand (_17650_, _14050_, _26656_);
  nand (_26658_, _17650_, _17649_);
  nand (_17651_, _14799_, _14048_);
  nand (_17652_, _14050_, _26660_);
  nand (_26662_, _17652_, _17651_);
  nand (_17653_, _14802_, _14048_);
  nand (_17654_, _14050_, _26664_);
  nand (_26666_, _17654_, _17653_);
  nand (_17655_, _14805_, _14048_);
  nand (_17656_, _14050_, _26668_);
  nand (_26670_, _17656_, _17655_);
  nand (_17657_, _14808_, _14048_);
  nand (_17658_, _14050_, _26672_);
  nand (_26674_, _17658_, _17657_);
  nand (_17659_, _14044_, _14789_);
  nand (_17660_, _14046_, _26676_);
  nand (_26678_, _17660_, _17659_);
  nand (_17661_, _14792_, _14044_);
  nand (_17662_, _14046_, _26680_);
  nand (_26682_, _17662_, _17661_);
  nand (_17663_, _14795_, _14044_);
  nand (_17664_, _14046_, _26684_);
  nand (_26686_, _17664_, _17663_);
  nand (_17665_, _14799_, _14044_);
  nand (_17666_, _14046_, _26688_);
  nand (_26690_, _17666_, _17665_);
  nand (_17668_, _14802_, _14044_);
  nand (_17669_, _14046_, _26692_);
  nand (_26694_, _17669_, _17668_);
  nand (_17670_, _14805_, _14044_);
  nand (_17671_, _14046_, _26696_);
  nand (_26698_, _17671_, _17670_);
  nand (_17672_, _14808_, _14044_);
  nand (_17673_, _14046_, _26700_);
  nand (_26702_, _17673_, _17672_);
  nand (_17675_, _14040_, _14789_);
  nand (_17676_, _14042_, _26704_);
  nand (_26706_, _17676_, _17675_);
  nand (_17677_, _14792_, _14040_);
  nand (_17678_, _14042_, _26708_);
  nand (_26710_, _17678_, _17677_);
  nand (_17679_, _14795_, _14040_);
  nand (_17680_, _14042_, _26712_);
  nand (_26714_, _17680_, _17679_);
  nand (_17681_, _14799_, _14040_);
  nand (_17682_, _14042_, _26716_);
  nand (_26718_, _17682_, _17681_);
  nand (_17683_, _14802_, _14040_);
  nand (_17684_, _14042_, _26720_);
  nand (_26722_, _17684_, _17683_);
  nand (_17685_, _14805_, _14040_);
  nand (_17686_, _14042_, _26724_);
  nand (_26726_, _17686_, _17685_);
  nand (_17687_, _14808_, _14040_);
  nand (_17688_, _14042_, _26730_);
  nand (_26732_, _17688_, _17687_);
  nand (_17690_, _14036_, _14789_);
  nand (_17691_, _14038_, _26734_);
  nand (_26736_, _17691_, _17690_);
  nand (_17692_, _14792_, _14036_);
  nand (_17693_, _14038_, _26738_);
  nand (_26740_, _17693_, _17692_);
  nand (_17694_, _14795_, _14036_);
  nand (_17695_, _14038_, _26742_);
  nand (_26744_, _17695_, _17694_);
  nand (_17697_, _14799_, _14036_);
  nand (_17698_, _14038_, _26746_);
  nand (_26748_, _17698_, _17697_);
  nand (_17699_, _14802_, _14036_);
  nand (_17700_, _14038_, _26750_);
  nand (_26752_, _17700_, _17699_);
  nand (_17701_, _14805_, _14036_);
  nand (_17702_, _14038_, _26754_);
  nand (_26756_, _17702_, _17701_);
  nand (_17703_, _14808_, _14036_);
  nand (_17705_, _14038_, _26758_);
  nand (_26760_, _17705_, _17703_);
  nand (_17706_, _14029_, _14789_);
  nand (_17707_, _14032_, _26762_);
  nand (_26764_, _17707_, _17706_);
  nand (_17708_, _14792_, _14029_);
  nand (_17709_, _14032_, _26766_);
  nand (_26768_, _17709_, _17708_);
  nand (_17710_, _14795_, _14029_);
  nand (_17711_, _14032_, _26770_);
  nand (_26772_, _17711_, _17710_);
  nand (_17712_, _14799_, _14029_);
  nand (_17713_, _14032_, _26774_);
  nand (_26776_, _17713_, _17712_);
  nand (_17714_, _14802_, _14029_);
  nand (_17715_, _14032_, _26778_);
  nand (_26780_, _17715_, _17714_);
  nand (_17716_, _14805_, _14029_);
  nand (_17717_, _14032_, _26782_);
  nand (_26784_, _17717_, _17716_);
  nand (_17718_, _14808_, _14029_);
  nand (_17719_, _14032_, _26786_);
  nand (_26788_, _17719_, _17718_);
  nand (_17720_, _14025_, _14789_);
  nand (_17721_, _14027_, _26790_);
  nand (_26792_, _17721_, _17720_);
  nand (_17722_, _14792_, _14025_);
  nand (_17723_, _14027_, _26794_);
  nand (_26796_, _17723_, _17722_);
  nand (_17724_, _14795_, _14025_);
  nand (_17726_, _14027_, _26798_);
  nand (_26800_, _17726_, _17724_);
  nand (_17727_, _14799_, _14025_);
  nand (_17728_, _14027_, _26802_);
  nand (_26804_, _17728_, _17727_);
  nand (_17729_, _14802_, _14025_);
  nand (_17730_, _14027_, _26806_);
  nand (_26808_, _17730_, _17729_);
  nand (_17731_, _14805_, _14025_);
  nand (_17732_, _14027_, _26811_);
  nand (_26813_, _17732_, _17731_);
  nand (_17734_, _14808_, _14025_);
  nand (_17735_, _14027_, _26815_);
  nand (_26817_, _17735_, _17734_);
  nand (_17736_, _14021_, _14789_);
  nand (_17737_, _14023_, _26819_);
  nand (_26821_, _17737_, _17736_);
  nand (_17738_, _14792_, _14021_);
  nand (_17739_, _14023_, _26823_);
  nand (_26825_, _17739_, _17738_);
  nand (_17740_, _14795_, _14021_);
  nand (_17741_, _14023_, _26827_);
  nand (_26829_, _17741_, _17740_);
  nand (_17742_, _14799_, _14021_);
  nand (_17743_, _14023_, _26831_);
  nand (_26833_, _17743_, _17742_);
  nand (_17744_, _14802_, _14021_);
  nand (_17745_, _14023_, _26835_);
  nand (_26837_, _17745_, _17744_);
  nand (_17746_, _14805_, _14021_);
  nand (_17747_, _14023_, _26839_);
  nand (_26841_, _17747_, _17746_);
  nand (_17748_, _14808_, _14021_);
  nand (_17749_, _14023_, _26843_);
  nand (_26845_, _17749_, _17748_);
  nand (_17750_, _14017_, _14789_);
  nand (_17751_, _14019_, _26847_);
  nand (_26849_, _17751_, _17750_);
  nand (_17752_, _14792_, _14017_);
  nand (_17753_, _14019_, _26851_);
  nand (_26853_, _17753_, _17752_);
  nand (_17755_, _14795_, _14017_);
  nand (_17756_, _14019_, _26855_);
  nand (_26857_, _17756_, _17755_);
  nand (_17757_, _14799_, _14017_);
  nand (_17758_, _14019_, _26859_);
  nand (_26861_, _17758_, _17757_);
  nand (_17759_, _14802_, _14017_);
  nand (_17760_, _14019_, _26863_);
  nand (_26865_, _17760_, _17759_);
  nand (_17762_, _14805_, _14017_);
  nand (_17763_, _14019_, _26867_);
  nand (_26869_, _17763_, _17762_);
  nand (_17764_, _14808_, _14017_);
  nand (_17765_, _14019_, _26871_);
  nand (_26873_, _17765_, _17764_);
  nand (_17766_, _14013_, _14789_);
  nand (_17767_, _14015_, _26875_);
  nand (_26877_, _17767_, _17766_);
  nand (_17768_, _14792_, _14013_);
  nand (_17769_, _14015_, _26879_);
  nand (_26881_, _17769_, _17768_);
  nand (_17770_, _14795_, _14013_);
  nand (_17771_, _14015_, _26883_);
  nand (_26885_, _17771_, _17770_);
  nand (_17772_, _14799_, _14013_);
  nand (_17773_, _14015_, _26887_);
  nand (_26889_, _17773_, _17772_);
  nand (_17774_, _14802_, _14013_);
  nand (_17775_, _14015_, _26892_);
  nand (_26894_, _17775_, _17774_);
  nand (_17776_, _14805_, _14013_);
  nand (_17777_, _14015_, _26896_);
  nand (_26898_, _17777_, _17776_);
  nand (_17778_, _14808_, _14013_);
  nand (_17779_, _14015_, _26900_);
  nand (_26902_, _17779_, _17778_);
  nand (_17780_, _14009_, _14789_);
  nand (_17781_, _14011_, _26904_);
  nand (_26906_, _17781_, _17780_);
  nand (_17783_, _14792_, _14009_);
  nand (_17784_, _14011_, _26908_);
  nand (_26910_, _17784_, _17783_);
  nand (_17785_, _14795_, _14009_);
  nand (_17786_, _14011_, _26912_);
  nand (_26914_, _17786_, _17785_);
  nand (_17787_, _14799_, _14009_);
  nand (_17788_, _14011_, _26916_);
  nand (_26918_, _17788_, _17787_);
  nand (_17789_, _14802_, _14009_);
  nand (_17791_, _14011_, _26920_);
  nand (_26922_, _17791_, _17789_);
  nand (_17792_, _14805_, _14009_);
  nand (_17793_, _14011_, _26924_);
  nand (_26926_, _17793_, _17792_);
  nand (_17794_, _14808_, _14009_);
  nand (_17795_, _14011_, _26928_);
  nand (_26930_, _17795_, _17794_);
  nand (_17796_, _14005_, _14789_);
  nand (_17797_, _14007_, _26932_);
  nand (_26934_, _17797_, _17796_);
  nand (_17798_, _14792_, _14005_);
  nand (_17799_, _14007_, _26936_);
  nand (_26938_, _17799_, _17798_);
  nand (_17800_, _14795_, _14005_);
  nand (_17801_, _14007_, _26940_);
  nand (_26942_, _17801_, _17800_);
  nand (_17802_, _14799_, _14005_);
  nand (_17803_, _14007_, _26944_);
  nand (_26946_, _17803_, _17802_);
  nand (_17804_, _14802_, _14005_);
  nand (_17805_, _14007_, _26948_);
  nand (_26950_, _17805_, _17804_);
  nand (_17806_, _14805_, _14005_);
  nand (_17807_, _14007_, _26952_);
  nand (_26954_, _17807_, _17806_);
  nand (_17808_, _14808_, _14005_);
  nand (_17809_, _14007_, _26956_);
  nand (_26958_, _17809_, _17808_);
  nand (_17810_, _14001_, _14789_);
  nand (_17812_, _14003_, _26960_);
  nand (_26962_, _17812_, _17810_);
  nand (_17813_, _14792_, _14001_);
  nand (_17814_, _14003_, _26964_);
  nand (_26966_, _17814_, _17813_);
  nand (_17815_, _14795_, _14001_);
  nand (_17816_, _14003_, _26968_);
  nand (_26970_, _17816_, _17815_);
  nand (_17817_, _14799_, _14001_);
  nand (_17818_, _14003_, _26973_);
  nand (_26975_, _17818_, _17817_);
  nand (_17820_, _14802_, _14001_);
  nand (_17821_, _14003_, _26977_);
  nand (_26979_, _17821_, _17820_);
  nand (_17822_, _14805_, _14001_);
  nand (_17823_, _14003_, _26981_);
  nand (_26983_, _17823_, _17822_);
  nand (_17824_, _14808_, _14001_);
  nand (_17825_, _14003_, _26985_);
  nand (_26987_, _17825_, _17824_);
  nand (_17826_, _13996_, _14789_);
  nand (_17827_, _13999_, _26989_);
  nand (_26991_, _17827_, _17826_);
  nand (_17828_, _14792_, _13996_);
  nand (_17829_, _13999_, _26993_);
  nand (_26995_, _17829_, _17828_);
  nand (_17830_, _14795_, _13996_);
  nand (_17831_, _13999_, _26997_);
  nand (_26999_, _17831_, _17830_);
  nand (_17832_, _14799_, _13996_);
  nand (_17833_, _13999_, _27001_);
  nand (_27003_, _17833_, _17832_);
  nand (_17834_, _14802_, _13996_);
  nand (_17835_, _13999_, _27005_);
  nand (_27007_, _17835_, _17834_);
  nand (_17836_, _14805_, _13996_);
  nand (_17837_, _13999_, _27009_);
  nand (_27011_, _17837_, _17836_);
  nand (_17838_, _14808_, _13996_);
  nand (_17839_, _13999_, _27013_);
  nand (_27015_, _17839_, _17838_);
  nand (_17841_, _13992_, _14789_);
  nand (_17842_, _13994_, _27017_);
  nand (_27019_, _17842_, _17841_);
  nand (_17843_, _14792_, _13992_);
  nand (_17844_, _13994_, _27021_);
  nand (_27023_, _17844_, _17843_);
  nand (_17845_, _14795_, _13992_);
  nand (_17846_, _13994_, _27025_);
  nand (_27027_, _17846_, _17845_);
  nand (_17848_, _14799_, _13992_);
  nand (_17849_, _13994_, _27029_);
  nand (_27031_, _17849_, _17848_);
  nand (_17850_, _14802_, _13992_);
  nand (_17851_, _13994_, _27033_);
  nand (_27035_, _17851_, _17850_);
  nand (_17852_, _14805_, _13992_);
  nand (_17853_, _13994_, _27037_);
  nand (_27039_, _17853_, _17852_);
  nand (_17854_, _14808_, _13992_);
  nand (_17855_, _13994_, _27041_);
  nand (_27043_, _17855_, _17854_);
  nand (_17856_, _13988_, _14789_);
  nand (_17857_, _13990_, _27045_);
  nand (_27047_, _17857_, _17856_);
  nand (_17858_, _14792_, _13988_);
  nand (_17859_, _13990_, _27049_);
  nand (_27051_, _17859_, _17858_);
  nand (_17860_, _14795_, _13988_);
  nand (_17861_, _13990_, _27054_);
  nand (_27056_, _17861_, _17860_);
  nand (_17862_, _14799_, _13988_);
  nand (_17863_, _13990_, _27058_);
  nand (_27060_, _17863_, _17862_);
  nand (_17864_, _14802_, _13988_);
  nand (_17865_, _13990_, _27062_);
  nand (_27064_, _17865_, _17864_);
  nand (_17866_, _14805_, _13988_);
  nand (_17867_, _13990_, _27066_);
  nand (_27068_, _17867_, _17866_);
  nand (_17869_, _14808_, _13988_);
  nand (_17870_, _13990_, _27070_);
  nand (_27072_, _17870_, _17869_);
  nand (_17871_, _13984_, _14789_);
  nand (_17872_, _13986_, _27074_);
  nand (_27076_, _17872_, _17871_);
  nand (_17873_, _14792_, _13984_);
  nand (_17874_, _13986_, _27078_);
  nand (_27080_, _17874_, _17873_);
  nand (_17875_, _14795_, _13984_);
  nand (_17877_, _13986_, _27082_);
  nand (_27084_, _17877_, _17875_);
  nand (_17878_, _14799_, _13984_);
  nand (_17879_, _13986_, _27086_);
  nand (_27088_, _17879_, _17878_);
  nand (_17880_, _14802_, _13984_);
  nand (_17881_, _13986_, _27090_);
  nand (_27092_, _17881_, _17880_);
  nand (_17882_, _14805_, _13984_);
  nand (_17883_, _13986_, _27094_);
  nand (_27096_, _17883_, _17882_);
  nand (_17884_, _14808_, _13984_);
  nand (_17885_, _13986_, _27098_);
  nand (_27100_, _17885_, _17884_);
  nand (_17886_, _13980_, _14789_);
  nand (_17887_, _13982_, _27102_);
  nand (_27104_, _17887_, _17886_);
  nand (_17888_, _14792_, _13980_);
  nand (_17889_, _13982_, _27106_);
  nand (_27108_, _17889_, _17888_);
  nand (_17890_, _14795_, _13980_);
  nand (_17891_, _13982_, _27110_);
  nand (_27112_, _17891_, _17890_);
  nand (_17892_, _14799_, _13980_);
  nand (_17893_, _13982_, _27114_);
  nand (_27116_, _17893_, _17892_);
  nand (_17894_, _14802_, _13980_);
  nand (_17895_, _13982_, _27118_);
  nand (_27120_, _17895_, _17894_);
  nand (_17896_, _14805_, _13980_);
  nand (_17898_, _13982_, _27122_);
  nand (_27124_, _17898_, _17896_);
  nand (_17899_, _14808_, _13980_);
  nand (_17900_, _13982_, _27126_);
  nand (_27128_, _17900_, _17899_);
  nand (_17901_, _13976_, _14789_);
  nand (_17902_, _13978_, _27130_);
  nand (_27132_, _17902_, _17901_);
  nand (_17903_, _14792_, _13976_);
  nand (_17904_, _13978_, _27135_);
  nand (_27137_, _17904_, _17903_);
  nand (_17906_, _14795_, _13976_);
  nand (_17907_, _13978_, _27139_);
  nand (_27141_, _17907_, _17906_);
  nand (_17908_, _14799_, _13976_);
  nand (_17909_, _13978_, _27143_);
  nand (_27145_, _17909_, _17908_);
  nand (_17910_, _14802_, _13976_);
  nand (_17911_, _13978_, _27147_);
  nand (_27149_, _17911_, _17910_);
  nand (_17912_, _14805_, _13976_);
  nand (_17913_, _13978_, _27151_);
  nand (_27153_, _17913_, _17912_);
  nand (_17914_, _14808_, _13976_);
  nand (_17915_, _13978_, _27155_);
  nand (_27157_, _17915_, _17914_);
  nand (_17916_, _13972_, _14789_);
  nand (_17917_, _13974_, _27159_);
  nand (_27161_, _17917_, _17916_);
  nand (_17918_, _14792_, _13972_);
  nand (_17919_, _13974_, _27163_);
  nand (_27165_, _17919_, _17918_);
  nand (_17920_, _14795_, _13972_);
  nand (_17921_, _13974_, _27167_);
  nand (_27169_, _17921_, _17920_);
  nand (_17922_, _14799_, _13972_);
  nand (_17923_, _13974_, _27171_);
  nand (_27173_, _17923_, _17922_);
  nand (_17924_, _14802_, _13972_);
  nand (_17925_, _13974_, _27175_);
  nand (_27177_, _17925_, _17924_);
  nand (_17927_, _14805_, _13972_);
  nand (_17928_, _13974_, _27179_);
  nand (_27181_, _17928_, _17927_);
  nand (_17929_, _14808_, _13972_);
  nand (_17930_, _13974_, _27183_);
  nand (_27185_, _17930_, _17929_);
  nand (_17931_, _13968_, _14789_);
  nand (_17932_, _13970_, _27187_);
  nand (_27189_, _17932_, _17931_);
  nand (_17934_, _14792_, _13968_);
  nand (_17935_, _13970_, _27191_);
  nand (_27193_, _17935_, _17934_);
  nand (_17936_, _14795_, _13968_);
  nand (_17937_, _13970_, _27195_);
  nand (_27197_, _17937_, _17936_);
  nand (_17938_, _14799_, _13968_);
  nand (_17939_, _13970_, _27199_);
  nand (_27201_, _17939_, _17938_);
  nand (_17940_, _14802_, _13968_);
  nand (_17941_, _13970_, _27203_);
  nand (_27205_, _17941_, _17940_);
  nand (_17942_, _14805_, _13968_);
  nand (_17943_, _13970_, _27207_);
  nand (_27209_, _17943_, _17942_);
  nand (_17944_, _14808_, _13968_);
  nand (_17945_, _13970_, _27211_);
  nand (_27213_, _17945_, _17944_);
  nand (_17946_, _13959_, _14789_);
  nand (_17947_, _13961_, _27216_);
  nand (_27218_, _17947_, _17946_);
  nand (_17948_, _14792_, _13959_);
  nand (_17949_, _13961_, _27220_);
  nand (_27222_, _17949_, _17948_);
  nand (_17950_, _14795_, _13959_);
  nand (_17951_, _13961_, _27224_);
  nand (_27226_, _17951_, _17950_);
  nand (_17952_, _14799_, _13959_);
  nand (_17953_, _13961_, _27228_);
  nand (_27230_, _17953_, _17952_);
  nand (_17955_, _14802_, _13959_);
  nand (_17956_, _13961_, _27232_);
  nand (_27234_, _17956_, _17955_);
  nand (_17957_, _14805_, _13959_);
  nand (_17958_, _13961_, _27236_);
  nand (_27238_, _17958_, _17957_);
  nand (_17959_, _14808_, _13959_);
  nand (_17960_, _13961_, _27240_);
  nand (_27242_, _17960_, _17959_);
  nand (_17961_, _13955_, _14789_);
  nand (_17963_, _13957_, _27244_);
  nand (_27246_, _17963_, _17961_);
  nand (_17964_, _14792_, _13955_);
  nand (_17965_, _13957_, _27248_);
  nand (_27250_, _17965_, _17964_);
  nand (_17966_, _14795_, _13955_);
  nand (_17967_, _13957_, _27252_);
  nand (_27254_, _17967_, _17966_);
  nand (_17968_, _14799_, _13955_);
  nand (_17969_, _13957_, _27256_);
  nand (_27258_, _17969_, _17968_);
  nand (_17970_, _14802_, _13955_);
  nand (_17971_, _13957_, _27260_);
  nand (_27262_, _17971_, _17970_);
  nand (_17972_, _14805_, _13955_);
  nand (_17973_, _13957_, _27264_);
  nand (_27266_, _17973_, _17972_);
  nand (_17974_, _14808_, _13955_);
  nand (_17975_, _13957_, _27268_);
  nand (_27270_, _17975_, _17974_);
  nand (_17977_, _13951_, _14789_);
  nand (_17978_, _13953_, _27272_);
  nand (_27274_, _17978_, _17977_);
  nand (_17979_, _14792_, _13951_);
  nand (_17980_, _13953_, _27276_);
  nand (_27278_, _17980_, _17979_);
  nand (_17981_, _14795_, _13951_);
  nand (_17982_, _13953_, _27280_);
  nand (_27282_, _17982_, _17981_);
  nand (_17983_, _14799_, _13951_);
  nand (_17985_, _13953_, _27284_);
  nand (_27286_, _17985_, _17983_);
  nand (_17986_, _14802_, _13951_);
  nand (_17987_, _13953_, _27288_);
  nand (_27290_, _17987_, _17986_);
  nand (_17988_, _14805_, _13951_);
  nand (_17989_, _13953_, _27292_);
  nand (_27294_, _17989_, _17988_);
  nand (_17990_, _14808_, _13951_);
  nand (_17991_, _13953_, _27297_);
  nand (_27299_, _17991_, _17990_);
  nand (_17993_, _13947_, _14789_);
  nand (_17994_, _13949_, _27301_);
  nand (_27303_, _17994_, _17993_);
  nand (_17995_, _14792_, _13947_);
  nand (_17996_, _13949_, _27305_);
  nand (_27307_, _17996_, _17995_);
  nand (_17997_, _14795_, _13947_);
  nand (_17998_, _13949_, _27309_);
  nand (_27311_, _17998_, _17997_);
  nand (_17999_, _14799_, _13947_);
  nand (_18000_, _13949_, _27313_);
  nand (_27315_, _18000_, _17999_);
  nand (_18001_, _14802_, _13947_);
  nand (_18002_, _13949_, _27317_);
  nand (_27319_, _18002_, _18001_);
  nand (_18003_, _14805_, _13947_);
  nand (_18004_, _13949_, _27321_);
  nand (_27323_, _18004_, _18003_);
  nand (_18005_, _14808_, _13947_);
  nand (_18006_, _13949_, _27325_);
  nand (_27327_, _18006_, _18005_);
  nand (_18007_, _13943_, _14789_);
  nand (_18008_, _13945_, _27329_);
  nand (_27331_, _18008_, _18007_);
  nand (_18009_, _14792_, _13943_);
  nand (_18010_, _13945_, _27333_);
  nand (_27335_, _18010_, _18009_);
  nand (_18011_, _14795_, _13943_);
  nand (_18012_, _13945_, _27337_);
  nand (_27339_, _18012_, _18011_);
  nand (_18014_, _14799_, _13943_);
  nand (_18015_, _13945_, _27341_);
  nand (_27343_, _18015_, _18014_);
  nand (_18016_, _14802_, _13943_);
  nand (_18017_, _13945_, _27345_);
  nand (_27347_, _18017_, _18016_);
  nand (_18018_, _14805_, _13943_);
  nand (_18019_, _13945_, _27349_);
  nand (_27351_, _18019_, _18018_);
  nand (_18021_, _14808_, _13943_);
  nand (_18022_, _13945_, _27353_);
  nand (_27355_, _18022_, _18021_);
  nand (_18023_, _13939_, _14789_);
  nand (_18024_, _13941_, _27357_);
  nand (_27359_, _18024_, _18023_);
  nand (_18025_, _14792_, _13939_);
  nand (_18026_, _13941_, _27361_);
  nand (_27363_, _18026_, _18025_);
  nand (_18027_, _14795_, _13939_);
  nand (_18028_, _13941_, _27365_);
  nand (_27367_, _18028_, _18027_);
  nand (_18029_, _14799_, _13939_);
  nand (_18030_, _13941_, _27369_);
  nand (_27371_, _18030_, _18029_);
  nand (_18031_, _14802_, _13939_);
  nand (_18032_, _13941_, _27373_);
  nand (_27375_, _18032_, _18031_);
  nand (_18033_, _14805_, _13939_);
  nand (_18034_, _13941_, _27378_);
  nand (_27380_, _18034_, _18033_);
  nand (_18035_, _14808_, _13939_);
  nand (_18036_, _13941_, _27382_);
  nand (_27384_, _18036_, _18035_);
  nand (_18037_, _13935_, _14789_);
  nand (_18038_, _13937_, _27386_);
  nand (_27388_, _18038_, _18037_);
  nand (_18039_, _14792_, _13935_);
  nand (_18040_, _13937_, _27390_);
  nand (_27392_, _18040_, _18039_);
  nand (_18042_, _14795_, _13935_);
  nand (_18043_, _13937_, _27394_);
  nand (_27396_, _18043_, _18042_);
  nand (_18044_, _14799_, _13935_);
  nand (_18045_, _13937_, _27398_);
  nand (_27400_, _18045_, _18044_);
  nand (_18046_, _14802_, _13935_);
  nand (_18047_, _13937_, _27402_);
  nand (_27404_, _18047_, _18046_);
  nand (_18048_, _14805_, _13935_);
  nand (_18050_, _13937_, _27406_);
  nand (_27408_, _18050_, _18048_);
  nand (_18051_, _14808_, _13935_);
  nand (_18052_, _13937_, _27410_);
  nand (_27412_, _18052_, _18051_);
  nand (_18053_, _13930_, _14789_);
  nand (_18054_, _13933_, _27414_);
  nand (_27416_, _18054_, _18053_);
  nand (_18055_, _14792_, _13930_);
  nand (_18056_, _13933_, _27418_);
  nand (_27420_, _18056_, _18055_);
  nand (_18057_, _14795_, _13930_);
  nand (_18058_, _13933_, _27422_);
  nand (_27424_, _18058_, _18057_);
  nand (_18059_, _14799_, _13930_);
  nand (_18060_, _13933_, _27426_);
  nand (_27428_, _18060_, _18059_);
  nand (_18061_, _14802_, _13930_);
  nand (_18062_, _13933_, _27430_);
  nand (_27432_, _18062_, _18061_);
  nand (_18063_, _14805_, _13930_);
  nand (_18064_, _13933_, _27434_);
  nand (_27436_, _18064_, _18063_);
  nand (_18065_, _14808_, _13930_);
  nand (_18066_, _13933_, _27438_);
  nand (_27440_, _18066_, _18065_);
  nand (_18067_, _13926_, _14789_);
  nand (_18068_, _13928_, _27442_);
  nand (_27444_, _18068_, _18067_);
  nand (_18069_, _14792_, _13926_);
  nand (_18070_, _13928_, _27446_);
  nand (_27448_, _18070_, _18069_);
  nand (_18071_, _14795_, _13926_);
  nand (_18072_, _13928_, _27450_);
  nand (_27452_, _18072_, _18071_);
  nand (_18073_, _14799_, _13926_);
  nand (_18074_, _13928_, _27454_);
  nand (_27456_, _18074_, _18073_);
  nand (_18075_, _14802_, _13926_);
  nand (_18076_, _13928_, _27459_);
  nand (_27461_, _18076_, _18075_);
  nand (_18078_, _14805_, _13926_);
  nand (_18079_, _13928_, _27463_);
  nand (_27465_, _18079_, _18078_);
  nand (_18080_, _14808_, _13926_);
  nand (_18081_, _13928_, _27467_);
  nand (_27469_, _18081_, _18080_);
  nand (_18082_, _13922_, _14789_);
  nand (_18083_, _13924_, _27471_);
  nand (_27473_, _18083_, _18082_);
  nand (_18085_, _14792_, _13922_);
  nand (_18086_, _13924_, _27475_);
  nand (_27477_, _18086_, _18085_);
  nand (_18087_, _14795_, _13922_);
  nand (_18088_, _13924_, _27479_);
  nand (_27481_, _18088_, _18087_);
  nand (_18089_, _14799_, _13922_);
  nand (_18090_, _13924_, _27483_);
  nand (_27485_, _18090_, _18089_);
  nand (_18091_, _14802_, _13922_);
  nand (_18092_, _13924_, _27487_);
  nand (_27489_, _18092_, _18091_);
  nand (_18093_, _14805_, _13922_);
  nand (_18094_, _13924_, _27491_);
  nand (_27493_, _18094_, _18093_);
  nand (_18095_, _14808_, _13922_);
  nand (_18096_, _13924_, _27495_);
  nand (_27497_, _18096_, _18095_);
  nand (_18097_, _13906_, _14789_);
  nand (_18098_, _13908_, _27499_);
  nand (_27501_, _18098_, _18097_);
  nand (_18099_, _14792_, _13906_);
  nand (_18100_, _13908_, _27503_);
  nand (_27505_, _18100_, _18099_);
  nand (_18101_, _14795_, _13906_);
  nand (_18102_, _13908_, _27507_);
  nand (_27509_, _18102_, _18101_);
  nand (_18103_, _14799_, _13906_);
  nand (_18104_, _13908_, _27511_);
  nand (_27513_, _18104_, _18103_);
  nand (_18106_, _14802_, _13906_);
  nand (_18107_, _13908_, _27515_);
  nand (_27517_, _18107_, _18106_);
  nand (_18108_, _14805_, _13906_);
  nand (_18109_, _13908_, _27519_);
  nand (_27521_, _18109_, _18108_);
  nand (_18110_, _14808_, _13906_);
  nand (_18111_, _13908_, _27523_);
  nand (_27525_, _18111_, _18110_);
  nand (_18112_, _13902_, _14789_);
  nand (_18114_, _13904_, _27527_);
  nand (_27529_, _18114_, _18112_);
  nand (_18115_, _14792_, _13902_);
  nand (_18116_, _13904_, _27531_);
  nand (_27533_, _18116_, _18115_);
  nand (_18117_, _14795_, _13902_);
  nand (_18118_, _13904_, _27535_);
  nand (_27537_, _18118_, _18117_);
  nand (_18119_, _14799_, _13902_);
  nand (_18120_, _13904_, _27541_);
  nand (_27543_, _18120_, _18119_);
  nand (_18121_, _14802_, _13902_);
  nand (_18122_, _13904_, _27545_);
  nand (_27547_, _18122_, _18121_);
  nand (_18123_, _14805_, _13902_);
  nand (_18124_, _13904_, _27549_);
  nand (_27551_, _18124_, _18123_);
  nand (_18125_, _14808_, _13902_);
  nand (_18126_, _13904_, _27553_);
  nand (_27555_, _18126_, _18125_);
  nand (_18127_, _13897_, _14789_);
  nand (_18128_, _13900_, _27557_);
  nand (_27559_, _18128_, _18127_);
  nand (_18129_, _14792_, _13897_);
  nand (_18130_, _13900_, _27561_);
  nand (_27563_, _18130_, _18129_);
  nand (_18131_, _14795_, _13897_);
  nand (_18132_, _13900_, _27565_);
  nand (_27567_, _18132_, _18131_);
  nand (_18133_, _14799_, _13897_);
  nand (_18135_, _13900_, _27569_);
  nand (_27571_, _18135_, _18133_);
  nand (_18136_, _14802_, _13897_);
  nand (_18137_, _13900_, _27573_);
  nand (_27575_, _18137_, _18136_);
  nand (_18138_, _14805_, _13897_);
  nand (_18139_, _13900_, _27577_);
  nand (_27579_, _18139_, _18138_);
  nand (_18140_, _14808_, _13897_);
  nand (_18141_, _13900_, _27581_);
  nand (_27583_, _18141_, _18140_);
  nand (_18143_, _13889_, _14789_);
  nand (_18144_, _13891_, _27585_);
  nand (_27587_, _18144_, _18143_);
  nand (_18145_, _14792_, _13889_);
  nand (_18146_, _13891_, _27589_);
  nand (_27591_, _18146_, _18145_);
  nand (_18147_, _14795_, _13889_);
  nand (_18148_, _13891_, _27593_);
  nand (_27595_, _18148_, _18147_);
  nand (_18149_, _14799_, _13889_);
  nand (_18150_, _13891_, _27597_);
  nand (_27599_, _18150_, _18149_);
  nand (_18151_, _14802_, _13889_);
  nand (_18152_, _13891_, _27601_);
  nand (_27603_, _18152_, _18151_);
  nand (_18153_, _14805_, _13889_);
  nand (_18154_, _13891_, _27605_);
  nand (_27607_, _18154_, _18153_);
  nand (_18155_, _14808_, _13889_);
  nand (_18156_, _13891_, _27609_);
  nand (_27611_, _18156_, _18155_);
  nand (_18157_, _13885_, _14789_);
  nand (_18158_, _13887_, _27613_);
  nand (_27615_, _18158_, _18157_);
  nand (_18159_, _14792_, _13885_);
  nand (_18160_, _13887_, _27617_);
  nand (_27619_, _18160_, _18159_);
  nand (_18161_, _14795_, _13885_);
  nand (_18162_, _13887_, _27622_);
  nand (_27624_, _18162_, _18161_);
  nand (_18164_, _14799_, _13885_);
  nand (_18165_, _13887_, _27626_);
  nand (_27628_, _18165_, _18164_);
  nand (_18166_, _14802_, _13885_);
  nand (_18167_, _13887_, _27630_);
  nand (_27632_, _18167_, _18166_);
  nand (_18168_, _14805_, _13885_);
  nand (_18169_, _13887_, _27634_);
  nand (_27636_, _18169_, _18168_);
  nand (_18171_, _14808_, _13885_);
  nand (_18172_, _13887_, _27638_);
  nand (_27640_, _18172_, _18171_);
  nand (_18173_, _13881_, _14789_);
  nand (_18174_, _13883_, _27642_);
  nand (_27644_, _18174_, _18173_);
  nand (_18175_, _14792_, _13881_);
  nand (_18176_, _13883_, _27646_);
  nand (_27648_, _18176_, _18175_);
  nand (_18177_, _14795_, _13881_);
  nand (_18178_, _13883_, _27650_);
  nand (_27652_, _18178_, _18177_);
  nand (_18179_, _14799_, _13881_);
  nand (_18180_, _13883_, _27654_);
  nand (_27656_, _18180_, _18179_);
  nand (_18181_, _14802_, _13881_);
  nand (_18182_, _13883_, _27658_);
  nand (_27660_, _18182_, _18181_);
  nand (_18183_, _14805_, _13881_);
  nand (_18184_, _13883_, _27662_);
  nand (_27664_, _18184_, _18183_);
  nand (_18185_, _14808_, _13881_);
  nand (_18186_, _13883_, _27666_);
  nand (_27668_, _18186_, _18185_);
  nand (_18187_, _13873_, _14789_);
  nand (_18188_, _13875_, _27670_);
  nand (_27672_, _18188_, _18187_);
  nand (_18189_, _14792_, _13873_);
  nand (_18190_, _13875_, _27674_);
  nand (_27676_, _18190_, _18189_);
  nand (_18192_, _14795_, _13873_);
  nand (_18193_, _13875_, _27678_);
  nand (_27680_, _18193_, _18192_);
  nand (_18194_, _14799_, _13873_);
  nand (_18195_, _13875_, _27682_);
  nand (_27684_, _18195_, _18194_);
  nand (_18196_, _14802_, _13873_);
  nand (_18197_, _13875_, _27686_);
  nand (_27688_, _18197_, _18196_);
  nand (_18198_, _14805_, _13873_);
  nand (_18200_, _13875_, _27690_);
  nand (_27692_, _18200_, _18198_);
  nand (_18201_, _14808_, _13873_);
  nand (_18202_, _13875_, _27694_);
  nand (_27696_, _18202_, _18201_);
  nand (_18203_, _13868_, _14789_);
  nand (_18204_, _13870_, _27698_);
  nand (_27700_, _18204_, _18203_);
  nand (_18205_, _14792_, _13868_);
  nand (_18206_, _13870_, _27703_);
  nand (_27705_, _18206_, _18205_);
  nand (_18207_, _14795_, _13868_);
  nand (_18208_, _13870_, _27707_);
  nand (_27709_, _18208_, _18207_);
  nand (_18209_, _14799_, _13868_);
  nand (_18210_, _13870_, _27711_);
  nand (_27713_, _18210_, _18209_);
  nand (_18211_, _14802_, _13868_);
  nand (_18212_, _13870_, _27715_);
  nand (_27717_, _18212_, _18211_);
  nand (_18213_, _14805_, _13868_);
  nand (_18214_, _13870_, _27719_);
  nand (_27721_, _18214_, _18213_);
  nand (_18215_, _14808_, _13868_);
  nand (_18216_, _13870_, _27723_);
  nand (_27725_, _18216_, _18215_);
  nand (_18217_, _13864_, _14789_);
  nand (_18218_, _13866_, _27727_);
  nand (_27729_, _18218_, _18217_);
  nand (_18219_, _14792_, _13864_);
  nand (_18221_, _13866_, _27731_);
  nand (_27733_, _18221_, _18219_);
  nand (_18222_, _14795_, _13864_);
  nand (_18223_, _13866_, _27735_);
  nand (_27737_, _18223_, _18222_);
  nand (_18224_, _14799_, _13864_);
  nand (_18225_, _13866_, _27739_);
  nand (_27741_, _18225_, _18224_);
  nand (_18226_, _14802_, _13864_);
  nand (_18227_, _13866_, _27743_);
  nand (_27745_, _18227_, _18226_);
  nand (_18229_, _14805_, _13864_);
  nand (_18230_, _13866_, _27747_);
  nand (_27749_, _18230_, _18229_);
  nand (_18231_, _14808_, _13864_);
  nand (_18232_, _13866_, _27751_);
  nand (_27753_, _18232_, _18231_);
  nand (_18233_, _13859_, _14789_);
  nand (_18234_, _13861_, _27755_);
  nand (_27757_, _18234_, _18233_);
  nand (_18235_, _14792_, _13859_);
  nand (_18236_, _13861_, _27759_);
  nand (_27761_, _18236_, _18235_);
  nand (_18237_, _14795_, _13859_);
  nand (_18238_, _13861_, _27763_);
  nand (_27765_, _18238_, _18237_);
  nand (_18239_, _14799_, _13859_);
  nand (_18240_, _13861_, _27767_);
  nand (_27769_, _18240_, _18239_);
  nand (_18241_, _14802_, _13859_);
  nand (_18242_, _13861_, _27771_);
  nand (_27773_, _18242_, _18241_);
  nand (_18243_, _14805_, _13859_);
  nand (_18244_, _13861_, _27775_);
  nand (_27777_, _18244_, _18243_);
  nand (_18245_, _14808_, _13859_);
  nand (_18246_, _13861_, _27779_);
  nand (_27781_, _18246_, _18245_);
  nand (_18247_, _13855_, _14789_);
  nand (_18248_, _13857_, _27784_);
  nand (_27786_, _18248_, _18247_);
  nand (_18250_, _14792_, _13855_);
  nand (_18251_, _13857_, _27788_);
  nand (_27790_, _18251_, _18250_);
  nand (_18252_, _14795_, _13855_);
  nand (_18253_, _13857_, _27792_);
  nand (_27794_, _18253_, _18252_);
  nand (_18254_, _14799_, _13855_);
  nand (_18255_, _13857_, _27796_);
  nand (_27798_, _18255_, _18254_);
  nand (_18257_, _14802_, _13855_);
  nand (_18258_, _13857_, _27800_);
  nand (_27802_, _18258_, _18257_);
  nand (_18259_, _14805_, _13855_);
  nand (_18260_, _13857_, _27804_);
  nand (_27806_, _18260_, _18259_);
  nand (_18261_, _14808_, _13855_);
  nand (_18262_, _13857_, _27808_);
  nand (_27810_, _18262_, _18261_);
  nand (_18263_, _13851_, _14789_);
  nand (_18265_, _13853_, _27812_);
  nand (_27814_, _18265_, _18263_);
  nand (_18266_, _14792_, _13851_);
  nand (_18267_, _13853_, _27816_);
  nand (_27818_, _18267_, _18266_);
  nand (_18268_, _14795_, _13851_);
  nand (_18269_, _13853_, _27820_);
  nand (_27822_, _18269_, _18268_);
  nand (_18270_, _14799_, _13851_);
  nand (_18271_, _13853_, _27824_);
  nand (_27826_, _18271_, _18270_);
  nand (_18272_, _14802_, _13851_);
  nand (_18273_, _13853_, _27828_);
  nand (_27830_, _18273_, _18272_);
  nand (_18274_, _14805_, _13851_);
  nand (_18275_, _13853_, _27832_);
  nand (_27834_, _18275_, _18274_);
  nand (_18276_, _14808_, _13851_);
  nand (_18277_, _13853_, _27836_);
  nand (_27838_, _18277_, _18276_);
  nand (_18279_, _13847_, _14789_);
  nand (_18280_, _13849_, _27840_);
  nand (_27842_, _18280_, _18279_);
  nand (_18281_, _14792_, _13847_);
  nand (_18282_, _13849_, _27844_);
  nand (_27846_, _18282_, _18281_);
  nand (_18283_, _14795_, _13847_);
  nand (_18284_, _13849_, _27848_);
  nand (_27850_, _18284_, _18283_);
  nand (_18285_, _14799_, _13847_);
  nand (_18287_, _13849_, _27852_);
  nand (_27854_, _18287_, _18285_);
  nand (_18288_, _14802_, _13847_);
  nand (_18289_, _13849_, _27856_);
  nand (_27858_, _18289_, _18288_);
  nand (_18290_, _14805_, _13847_);
  nand (_18291_, _13849_, _27860_);
  nand (_27862_, _18291_, _18290_);
  nand (_18292_, _14808_, _13847_);
  nand (_18293_, _13849_, _27865_);
  nand (_27867_, _18293_, _18292_);
  nand (_18294_, _13843_, _14789_);
  nand (_18295_, _13845_, _27869_);
  nand (_27871_, _18295_, _18294_);
  nand (_18296_, _14792_, _13843_);
  nand (_18297_, _13845_, _27873_);
  nand (_27875_, _18297_, _18296_);
  nand (_18298_, _14795_, _13843_);
  nand (_18299_, _13845_, _27877_);
  nand (_27879_, _18299_, _18298_);
  nand (_18300_, _14799_, _13843_);
  nand (_18301_, _13845_, _27881_);
  nand (_27883_, _18301_, _18300_);
  nand (_18302_, _14802_, _13843_);
  nand (_18303_, _13845_, _27885_);
  nand (_27887_, _18303_, _18302_);
  nand (_18304_, _14805_, _13843_);
  nand (_18305_, _13845_, _27889_);
  nand (_27891_, _18305_, _18304_);
  nand (_18306_, _14808_, _13843_);
  nand (_18308_, _13845_, _27893_);
  nand (_27895_, _18308_, _18306_);
  nand (_18309_, _13835_, _14789_);
  nand (_18310_, _13837_, _27897_);
  nand (_27899_, _18310_, _18309_);
  nand (_18311_, _14792_, _13835_);
  nand (_18312_, _13837_, _27901_);
  nand (_27903_, _18312_, _18311_);
  nand (_18313_, _14795_, _13835_);
  nand (_18314_, _13837_, _27905_);
  nand (_27907_, _18314_, _18313_);
  nand (_18316_, _14799_, _13835_);
  nand (_18317_, _13837_, _27909_);
  nand (_27911_, _18317_, _18316_);
  nand (_18318_, _14802_, _13835_);
  nand (_18319_, _13837_, _27913_);
  nand (_27915_, _18319_, _18318_);
  nand (_18320_, _14805_, _13835_);
  nand (_18321_, _13837_, _27917_);
  nand (_27919_, _18321_, _18320_);
  nand (_18322_, _14808_, _13835_);
  nand (_18323_, _13837_, _27921_);
  nand (_27923_, _18323_, _18322_);
  nand (_18324_, _13826_, _14789_);
  nand (_18325_, _13828_, _27925_);
  nand (_27927_, _18325_, _18324_);
  nand (_18326_, _14792_, _13826_);
  nand (_18327_, _13828_, _27929_);
  nand (_27931_, _18327_, _18326_);
  nand (_18328_, _14795_, _13826_);
  nand (_18329_, _13828_, _27933_);
  nand (_27935_, _18329_, _18328_);
  nand (_18330_, _14799_, _13826_);
  nand (_18331_, _13828_, _27937_);
  nand (_27939_, _18331_, _18330_);
  nand (_18332_, _14802_, _13826_);
  nand (_18333_, _13828_, _27941_);
  nand (_27943_, _18333_, _18332_);
  nand (_18334_, _14805_, _13826_);
  nand (_18335_, _13828_, _27946_);
  nand (_27948_, _18335_, _18334_);
  nand (_18337_, _14808_, _13826_);
  nand (_18338_, _13828_, _27950_);
  nand (_27952_, _18338_, _18337_);
  nand (_18339_, _13813_, _14789_);
  nand (_18340_, _13815_, _27954_);
  nand (_27956_, _18340_, _18339_);
  nand (_18341_, _14792_, _13813_);
  nand (_18342_, _13815_, _27958_);
  nand (_27960_, _18342_, _18341_);
  nand (_18344_, _14795_, _13813_);
  nand (_18345_, _13815_, _27962_);
  nand (_27964_, _18345_, _18344_);
  nand (_18346_, _14799_, _13813_);
  nand (_18347_, _13815_, _27966_);
  nand (_27968_, _18347_, _18346_);
  nand (_18348_, _14802_, _13813_);
  nand (_18349_, _13815_, _27970_);
  nand (_27972_, _18349_, _18348_);
  nand (_18350_, _14805_, _13813_);
  nand (_18351_, _13815_, _27974_);
  nand (_27976_, _18351_, _18350_);
  nand (_18352_, _14808_, _13813_);
  nand (_18353_, _13815_, _27978_);
  nand (_27980_, _18353_, _18352_);
  nand (_18354_, _13809_, _14789_);
  nand (_18355_, _13811_, _27982_);
  nand (_27984_, _18355_, _18354_);
  nand (_18356_, _14792_, _13809_);
  nand (_18357_, _13811_, _27986_);
  nand (_27988_, _18357_, _18356_);
  nand (_18358_, _14795_, _13809_);
  nand (_18359_, _13811_, _27990_);
  nand (_27992_, _18359_, _18358_);
  nand (_18360_, _14799_, _13809_);
  nand (_18361_, _13811_, _27994_);
  nand (_27996_, _18361_, _18360_);
  nand (_18362_, _14802_, _13809_);
  nand (_18363_, _13811_, _27998_);
  nand (_28000_, _18363_, _18362_);
  nand (_18365_, _14805_, _13809_);
  nand (_18366_, _13811_, _28002_);
  nand (_28004_, _18366_, _18365_);
  nand (_18367_, _14808_, _13809_);
  nand (_18368_, _13811_, _28006_);
  nand (_28008_, _18368_, _18367_);
  nand (_18369_, _13805_, _14789_);
  nand (_18370_, _13807_, _28010_);
  nand (_28012_, _18370_, _18369_);
  nand (_18371_, _14792_, _13805_);
  nand (_18373_, _13807_, _28014_);
  nand (_28016_, _18373_, _18371_);
  nand (_18374_, _14795_, _13805_);
  nand (_18375_, _13807_, _28018_);
  nand (_28020_, _18375_, _18374_);
  nand (_18376_, _14799_, _13805_);
  nand (_18377_, _13807_, _28022_);
  nand (_28024_, _18377_, _18376_);
  nand (_18378_, _14802_, _13805_);
  nand (_18379_, _13807_, _28027_);
  nand (_28029_, _18379_, _18378_);
  nand (_18380_, _14805_, _13805_);
  nand (_18381_, _13807_, _28031_);
  nand (_28033_, _18381_, _18380_);
  nand (_18382_, _14808_, _13805_);
  nand (_18383_, _13807_, _28035_);
  nand (_28037_, _18383_, _18382_);
  nand (_18384_, _13801_, _14789_);
  nand (_18385_, _13803_, _28039_);
  nand (_28041_, _18385_, _18384_);
  nand (_18386_, _14792_, _13801_);
  nand (_18387_, _13803_, _28043_);
  nand (_28045_, _18387_, _18386_);
  nand (_18388_, _14795_, _13801_);
  nand (_18389_, _13803_, _28047_);
  nand (_28049_, _18389_, _18388_);
  nand (_18390_, _14799_, _13801_);
  nand (_18391_, _13803_, _28051_);
  nand (_28053_, _18391_, _18390_);
  nand (_18392_, _14802_, _13801_);
  nand (_18394_, _13803_, _28055_);
  nand (_28057_, _18394_, _18392_);
  nand (_18395_, _14805_, _13801_);
  nand (_18396_, _13803_, _28059_);
  nand (_28061_, _18396_, _18395_);
  nand (_18397_, _14808_, _13801_);
  nand (_18398_, _13803_, _28063_);
  nand (_28065_, _18398_, _18397_);
  nand (_18399_, _13711_, _14789_);
  nand (_18400_, _13713_, _28067_);
  nand (_28069_, _18400_, _18399_);
  nand (_18402_, _14792_, _13711_);
  nand (_18403_, _13713_, _28071_);
  nand (_28073_, _18403_, _18402_);
  nand (_18404_, _14795_, _13711_);
  nand (_18405_, _13713_, _28075_);
  nand (_28077_, _18405_, _18404_);
  nand (_18406_, _14799_, _13711_);
  nand (_18407_, _13713_, _28079_);
  nand (_28081_, _18407_, _18406_);
  nand (_18408_, _14802_, _13711_);
  nand (_18409_, _13713_, _28083_);
  nand (_28085_, _18409_, _18408_);
  nand (_18410_, _14805_, _13711_);
  nand (_18411_, _13713_, _28087_);
  nand (_28089_, _18411_, _18410_);
  nand (_18412_, _14808_, _13711_);
  nand (_18413_, _13713_, _28091_);
  nand (_28093_, _18413_, _18412_);
  nand (_18414_, _13705_, _14789_);
  nand (_18415_, _13707_, _28095_);
  nand (_28097_, _18415_, _18414_);
  nand (_18416_, _14792_, _13705_);
  nand (_18417_, _13707_, _28099_);
  nand (_28101_, _18417_, _18416_);
  nand (_18418_, _14795_, _13705_);
  nand (_18419_, _13707_, _28103_);
  nand (_28105_, _18419_, _18418_);
  nand (_18420_, _14799_, _13705_);
  nand (_18421_, _13707_, _28108_);
  nand (_28110_, _18421_, _18420_);
  nand (_18423_, _14802_, _13705_);
  nand (_18424_, _13707_, _28112_);
  nand (_28114_, _18424_, _18423_);
  nand (_18425_, _14805_, _13705_);
  nand (_18426_, _13707_, _28116_);
  nand (_28118_, _18426_, _18425_);
  nand (_18427_, _14808_, _13705_);
  nand (_18428_, _13707_, _28120_);
  nand (_28122_, _18428_, _18427_);
  nand (_18430_, _13699_, _14789_);
  nand (_18431_, _13701_, _28124_);
  nand (_28126_, _18431_, _18430_);
  nand (_18432_, _14792_, _13699_);
  nand (_18433_, _13701_, _28128_);
  nand (_28130_, _18433_, _18432_);
  nand (_18434_, _14795_, _13699_);
  nand (_18435_, _13701_, _28132_);
  nand (_28134_, _18435_, _18434_);
  nand (_18436_, _14799_, _13699_);
  nand (_18437_, _13701_, _28136_);
  nand (_28138_, _18437_, _18436_);
  nand (_18438_, _14802_, _13699_);
  nand (_18439_, _13701_, _28140_);
  nand (_28142_, _18439_, _18438_);
  nand (_18440_, _14805_, _13699_);
  nand (_18441_, _13701_, _28144_);
  nand (_28146_, _18441_, _18440_);
  nand (_18442_, _14808_, _13699_);
  nand (_18443_, _13701_, _28148_);
  nand (_28150_, _18443_, _18442_);
  nand (_18444_, _13689_, _14789_);
  nand (_18445_, _13691_, _28152_);
  nand (_28154_, _18445_, _18444_);
  nand (_18446_, _14792_, _13689_);
  nand (_18447_, _13691_, _28156_);
  nand (_28158_, _18447_, _18446_);
  nand (_18448_, _14795_, _13689_);
  nand (_18449_, _13691_, _28160_);
  nand (_28162_, _18449_, _18448_);
  nand (_18451_, _14799_, _13689_);
  nand (_18452_, _13691_, _28164_);
  nand (_28166_, _18452_, _18451_);
  nand (_18453_, _14802_, _13689_);
  nand (_18454_, _13691_, _28168_);
  nand (_28170_, _18454_, _18453_);
  nand (_18455_, _14805_, _13689_);
  nand (_18456_, _13691_, _28172_);
  nand (_28174_, _18456_, _18455_);
  nand (_18457_, _14808_, _13689_);
  nand (_18459_, _13691_, _28176_);
  nand (_28178_, _18459_, _18457_);
  nand (_18460_, _13683_, _14789_);
  nand (_18461_, _13685_, _28180_);
  nand (_28182_, _18461_, _18460_);
  nand (_18462_, _14792_, _13683_);
  nand (_18463_, _13685_, _28184_);
  nand (_28186_, _18463_, _18462_);
  nand (_18464_, _14795_, _13683_);
  nand (_18465_, _13685_, _28189_);
  nand (_28191_, _18465_, _18464_);
  nand (_18466_, _14799_, _13683_);
  nand (_18467_, _13685_, _28193_);
  nand (_28195_, _18467_, _18466_);
  nand (_18468_, _14802_, _13683_);
  nand (_18469_, _13685_, _28197_);
  nand (_28199_, _18469_, _18468_);
  nand (_18470_, _14805_, _13683_);
  nand (_18471_, _13685_, _28201_);
  nand (_28203_, _18471_, _18470_);
  nand (_18472_, _14808_, _13683_);
  nand (_18473_, _13685_, _28205_);
  nand (_28207_, _18473_, _18472_);
  nand (_18474_, _13784_, _14789_);
  nand (_18475_, _13786_, _28209_);
  nand (_28211_, _18475_, _18474_);
  nand (_18476_, _14792_, _13784_);
  nand (_18477_, _13786_, _28213_);
  nand (_28215_, _18477_, _18476_);
  nand (_18478_, _14795_, _13784_);
  nand (_18480_, _13786_, _28217_);
  nand (_28219_, _18480_, _18478_);
  nand (_18481_, _14799_, _13784_);
  nand (_18482_, _13786_, _28221_);
  nand (_28223_, _18482_, _18481_);
  nand (_18483_, _14802_, _13784_);
  nand (_18484_, _13786_, _28225_);
  nand (_28227_, _18484_, _18483_);
  nand (_18485_, _14805_, _13784_);
  nand (_18486_, _13786_, _28229_);
  nand (_28231_, _18486_, _18485_);
  nand (_18488_, _14808_, _13784_);
  nand (_18489_, _13786_, _28233_);
  nand (_28235_, _18489_, _18488_);
  nand (_18490_, _13677_, _14789_);
  nand (_18491_, _13679_, _28237_);
  nand (_28239_, _18491_, _18490_);
  nand (_18492_, _14792_, _13677_);
  nand (_18493_, _13679_, _28241_);
  nand (_28243_, _18493_, _18492_);
  nand (_18494_, _14795_, _13677_);
  nand (_18495_, _13679_, _28245_);
  nand (_28247_, _18495_, _18494_);
  nand (_18496_, _14799_, _13677_);
  nand (_18497_, _13679_, _28249_);
  nand (_28251_, _18497_, _18496_);
  nand (_18498_, _14802_, _13677_);
  nand (_18499_, _13679_, _28253_);
  nand (_28255_, _18499_, _18498_);
  nand (_18500_, _14805_, _13677_);
  nand (_18501_, _13679_, _28257_);
  nand (_28259_, _18501_, _18500_);
  nand (_18502_, _14808_, _13677_);
  nand (_18503_, _13679_, _28261_);
  nand (_28263_, _18503_, _18502_);
  nand (_18504_, _13671_, _14789_);
  nand (_18505_, _13673_, _28265_);
  nand (_28267_, _18505_, _18504_);
  nand (_18506_, _14792_, _13671_);
  nand (_18507_, _13673_, _28270_);
  nand (_28272_, _18507_, _18506_);
  nand (_18509_, _14795_, _13671_);
  nand (_18510_, _13673_, _28274_);
  nand (_28276_, _18510_, _18509_);
  nand (_18511_, _14799_, _13671_);
  nand (_18512_, _13673_, _28278_);
  nand (_28280_, _18512_, _18511_);
  nand (_18513_, _14802_, _13671_);
  nand (_18514_, _13673_, _28282_);
  nand (_28284_, _18514_, _18513_);
  nand (_18516_, _14805_, _13671_);
  nand (_18517_, _13673_, _28286_);
  nand (_28288_, _18517_, _18516_);
  nand (_18518_, _14808_, _13671_);
  nand (_18519_, _13673_, _28290_);
  nand (_28292_, _18519_, _18518_);
  nand (_18520_, _13660_, _14789_);
  nand (_18521_, _13662_, _28294_);
  nand (_28296_, _18521_, _18520_);
  nand (_18522_, _14792_, _13660_);
  nand (_18523_, _13662_, _28298_);
  nand (_28300_, _18523_, _18522_);
  nand (_18524_, _14795_, _13660_);
  nand (_18525_, _13662_, _28302_);
  nand (_28304_, _18525_, _18524_);
  nand (_18526_, _14799_, _13660_);
  nand (_18527_, _13662_, _28306_);
  nand (_28308_, _18527_, _18526_);
  nand (_18528_, _14802_, _13660_);
  nand (_18529_, _13662_, _28310_);
  nand (_28312_, _18529_, _18528_);
  nand (_18530_, _14805_, _13660_);
  nand (_18531_, _13662_, _28314_);
  nand (_28316_, _18531_, _18530_);
  nand (_18532_, _14808_, _13660_);
  nand (_18533_, _13662_, _28318_);
  nand (_28320_, _18533_, _18532_);
  nand (_18534_, _13788_, _14789_);
  nand (_18535_, _13790_, _28322_);
  nand (_28324_, _18535_, _18534_);
  nand (_18536_, _14792_, _13788_);
  nand (_18537_, _13790_, _28326_);
  nand (_28328_, _18537_, _18536_);
  nand (_18538_, _14795_, _13788_);
  nand (_18539_, _13790_, _28330_);
  nand (_28332_, _18539_, _18538_);
  nand (_18540_, _14799_, _13788_);
  nand (_18541_, _13790_, _28334_);
  nand (_28336_, _18541_, _18540_);
  nand (_18542_, _14802_, _13788_);
  nand (_18544_, _13790_, _28338_);
  nand (_28340_, _18544_, _18542_);
  nand (_18545_, _14805_, _13788_);
  nand (_18546_, _13790_, _28342_);
  nand (_28344_, _18546_, _18545_);
  nand (_18547_, _14808_, _13788_);
  nand (_18548_, _13790_, _28346_);
  nand (_28348_, _18548_, _18547_);
  nand (_18549_, _13651_, _14789_);
  nand (_18550_, _13653_, _28352_);
  nand (_28354_, _18550_, _18549_);
  nand (_18553_, _14792_, _13651_);
  nand (_18554_, _13653_, _28356_);
  nand (_28358_, _18554_, _18553_);
  nand (_18555_, _14795_, _13651_);
  nand (_18556_, _13653_, _28360_);
  nand (_28362_, _18556_, _18555_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _33880_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _33880_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _33880_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _33880_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _33880_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _33880_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _33880_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _33880_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _33904_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _33904_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _33904_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _33904_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _33904_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _33904_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _33904_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _33904_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _33900_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _33900_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _33900_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _33900_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _33900_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _33900_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _33900_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _33900_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _33896_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _33896_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _33896_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _33896_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _33896_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _33896_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _33896_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _33896_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _33892_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _33892_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _33892_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _33892_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _33892_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _33892_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _33892_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _33892_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _33888_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _33888_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _33888_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _33888_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _33888_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _33888_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _33888_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _33888_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _33884_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _33884_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _33884_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _33884_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _33884_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _33884_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _33884_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _33884_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _33940_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _33940_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _33940_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _33940_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _33940_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _33940_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _33940_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _33940_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _33936_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _33936_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _33936_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _33936_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _33936_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _33936_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _33936_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _33936_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _33932_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _33932_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _33932_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _33932_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _33932_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _33932_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _33932_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _33932_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _33928_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _33928_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _33928_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _33928_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _33928_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _33928_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _33928_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _33928_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _33924_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _33924_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _33924_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _33924_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _33924_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _33924_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _33924_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _33924_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _33920_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _33920_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _33920_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _33920_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _33920_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _33920_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _33920_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _33920_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _33916_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _33916_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _33916_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _33916_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _33916_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _33916_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _33916_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _33916_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _33912_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _33912_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _33912_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _33912_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _33912_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _33912_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _33912_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _33912_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _33908_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _33908_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _33908_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _33908_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _33908_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _33908_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _33908_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _33908_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _33955_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _33505_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _33505_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _33505_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _33505_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _33505_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _33505_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _33505_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _33505_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _33505_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _33505_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _33505_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _33505_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _33505_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _33505_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _33505_[15]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _32981_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _32980_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _32982_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _32983_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _32984_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _32985_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _32986_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _32979_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _32987_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _32988_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _32989_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _32990_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _32991_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _32992_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _32993_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _32994_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _32964_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _32963_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _32965_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _32966_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _32967_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _32968_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _32969_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _32970_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _32971_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _32972_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _32973_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _32974_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _32975_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _32976_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _32977_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _32978_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _32997_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _32998_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _32999_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _33000_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _33001_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _33002_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _33003_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _32995_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _33004_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _33005_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _33006_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _33007_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _33008_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _33009_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _33010_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _32996_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _33011_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _33012_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _33013_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _33014_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _33015_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _33016_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _33017_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _33041_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _33042_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _33020_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _33047_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _33046_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _33021_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _33045_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _33022_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _33044_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _33043_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _33048_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _33051_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _33050_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _33049_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _33040_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _33023_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _33024_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _33039_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _33025_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _33038_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _33026_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _33037_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _33036_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _33027_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _33018_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _33019_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _33028_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _33052_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _33029_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _33053_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _33033_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _33035_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _33030_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _33034_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _33031_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _33032_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _33255_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _33256_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _33257_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _33258_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _33259_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _33260_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _33261_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _33232_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _33262_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _33263_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _33264_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _33265_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _33266_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _33267_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _33268_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _33217_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _33269_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _33270_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _33271_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _33272_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _33273_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _33274_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _33275_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _33218_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _33276_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _33277_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _33278_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _33279_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _33280_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _33231_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _33230_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _33219_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _33229_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _33228_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _33227_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _33226_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _33225_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _33224_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _33239_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _33220_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _33240_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _33243_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _33244_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _33247_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _33248_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _33234_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _33235_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _33221_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _33236_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _33237_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _33238_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _33241_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _33242_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _33245_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _33246_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _33222_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _33249_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _33250_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _33251_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _33252_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _33253_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _33254_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _33233_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _33223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _35657_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _35657_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _35657_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _35657_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _35657_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _35657_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _35657_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _35657_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _35657_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _35657_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _35657_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _35657_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _35657_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _35657_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _35657_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _35657_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _35658_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _35658_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _35658_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _35658_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _35658_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _35658_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _35658_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _35658_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _35658_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _35658_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _35658_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _35658_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _35658_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _35658_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _35658_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _35658_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _33056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _33167_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _33168_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _33169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _33170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _33057_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _33171_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _33172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _33173_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _33174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _33175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _33176_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _33177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _33058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _33059_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _33060_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _33178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _33179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _33180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _33181_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _33182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _33183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _33184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _33185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _33186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _33187_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _33188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _33189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _33190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _33191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _33192_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _33061_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _33193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _33194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _33195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _33196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _33197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _33198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _33199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _33200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _33201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _33202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _33203_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _33063_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _33098_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _33097_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _33096_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _33062_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _33064_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _33065_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _33066_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _33095_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _33094_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _33092_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _33093_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _33108_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _33104_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _33146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _33067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _33122_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _33166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _33068_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _33069_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _33070_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _33159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _33139_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _33142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _33163_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _33150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _33145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _33148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _33071_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _33072_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _33073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _33147_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _33152_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _33151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _33074_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _33105_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _33107_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _33106_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _33164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _33114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _33111_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _33090_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _33121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _33128_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _33125_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _33124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _33135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _33149_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _33054_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _33086_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _33134_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _33087_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _33088_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _33102_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _33120_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _33083_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _33143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _33119_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _33126_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _33161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _33115_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _33157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _33133_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _33110_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _33113_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _33109_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _33075_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _33158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _33155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _33136_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _33137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _33117_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _33055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _33081_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _33082_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _33141_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _33131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _33116_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _33154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _33129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _33138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _33144_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _33091_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _33130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _33132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _33162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _33156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _33084_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _33153_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _33089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _33112_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _33140_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _33160_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _33165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _33118_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _33127_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _33101_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _33103_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _33076_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _33077_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _33078_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _33079_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _33123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _33100_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _33085_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _33099_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _33080_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _33205_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _33208_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _33209_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _33210_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _33211_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _33212_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _33213_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _33214_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _33206_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _33207_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _33215_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _33216_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _33204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _37411_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _37411_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _37411_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _37411_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _37411_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _37411_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _37411_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _37411_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _37410_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _37410_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _37410_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _37410_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _37410_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _37410_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _37410_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _37410_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _37409_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _37409_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _37409_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _37409_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _37409_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _37409_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _37409_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _37409_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _37408_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _37408_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _37408_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _37408_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _37408_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _37408_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _37408_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _37408_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _37407_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _37407_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _37407_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _37407_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _37407_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _37407_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _37407_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _37407_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _37406_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _37406_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _37406_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _37406_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _37406_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _37406_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _37406_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _37406_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _37405_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _37405_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _37405_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _37405_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _37405_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _37405_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _37405_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _37405_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _37404_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _37404_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _37404_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _37404_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _37404_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _37404_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _37404_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _37404_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _37403_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _37403_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _37403_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _37403_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _37403_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _37403_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _37403_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _37403_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _37401_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _37401_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _37401_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _37401_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _37401_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _37401_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _37401_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _37401_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _37400_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _37400_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _37400_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _37400_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _37400_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _37400_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _37400_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _37400_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _37399_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _37399_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _37399_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _37399_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _37399_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _37399_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _37399_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _37399_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _37398_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _37398_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _37398_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _37398_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _37398_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _37398_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _37398_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _37398_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _37397_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _37397_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _37397_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _37397_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _37397_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _37397_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _37397_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _37397_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _37396_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _37396_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _37396_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _37396_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _37396_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _37396_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _37396_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _37396_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _37395_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _37395_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _37395_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _37395_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _37395_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _37395_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _37395_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _37395_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _37394_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _37394_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _37394_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _37394_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _37394_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _37394_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _37394_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _37394_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _37393_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _37393_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _37393_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _37393_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _37393_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _37393_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _37393_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _37393_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _37392_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _37392_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _37392_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _37392_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _37392_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _37392_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _37392_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _37392_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _37390_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _37390_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _37390_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _37390_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _37390_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _37390_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _37390_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _37390_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _37389_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _37389_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _37389_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _37389_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _37389_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _37389_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _37389_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _37389_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _37388_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _37388_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _37388_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _37388_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _37388_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _37388_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _37388_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _37388_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _37387_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _37387_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _37387_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _37387_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _37387_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _37387_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _37387_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _37387_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _37386_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _37386_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _37386_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _37386_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _37386_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _37386_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _37386_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _37386_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _37385_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _37385_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _37385_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _37385_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _37385_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _37385_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _37385_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _37385_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _37384_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _37384_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _37384_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _37384_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _37384_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _37384_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _37384_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _37384_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _37383_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _37383_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _37383_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _37383_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _37383_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _37383_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _37383_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _37383_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _37382_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _37382_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _37382_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _37382_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _37382_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _37382_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _37382_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _37382_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _37381_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _37381_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _37381_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _37381_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _37381_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _37381_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _37381_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _37381_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _37379_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _37379_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _37379_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _37379_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _37379_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _37379_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _37379_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _37379_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _37378_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _37378_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _37378_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _37378_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _37378_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _37378_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _37378_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _37378_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _37377_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _37377_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _37377_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _37377_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _37377_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _37377_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _37377_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _37377_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _37376_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _37376_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _37376_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _37376_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _37376_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _37376_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _37376_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _37376_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _37375_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _37375_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _37375_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _37375_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _37375_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _37375_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _37375_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _37375_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _37374_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _37374_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _37374_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _37374_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _37374_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _37374_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _37374_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _37374_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _37373_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _37373_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _37373_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _37373_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _37373_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _37373_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _37373_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _37373_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _37372_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _37372_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _37372_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _37372_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _37372_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _37372_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _37372_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _37372_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _37371_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _37371_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _37371_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _37371_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _37371_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _37371_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _37371_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _37371_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _37370_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _37370_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _37370_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _37370_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _37370_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _37370_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _37370_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _37370_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _37368_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _37368_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _37368_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _37368_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _37368_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _37368_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _37368_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _37368_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _37367_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _37367_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _37367_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _37367_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _37367_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _37367_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _37367_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _37367_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _37366_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _37366_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _37366_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _37366_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _37366_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _37366_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _37366_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _37366_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _37365_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _37365_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _37365_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _37365_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _37365_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _37365_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _37365_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _37365_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _37364_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _37364_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _37364_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _37364_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _37364_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _37364_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _37364_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _37364_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _37363_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _37363_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _37363_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _37363_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _37363_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _37363_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _37363_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _37363_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _37362_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _37362_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _37362_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _37362_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _37362_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _37362_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _37362_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _37362_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _37361_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _37361_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _37361_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _37361_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _37361_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _37361_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _37361_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _37361_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _37360_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _37360_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _37360_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _37360_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _37360_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _37360_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _37360_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _37360_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _37359_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _37359_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _37359_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _37359_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _37359_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _37359_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _37359_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _37359_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _37357_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _37357_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _37357_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _37357_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _37357_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _37357_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _37357_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _37357_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _37303_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _37303_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _37303_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _37303_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _37303_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _37303_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _37303_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _37303_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _37412_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _37412_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _37412_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _37412_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _37412_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _37412_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _37412_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _37412_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _37416_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _37416_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _37416_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _37416_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _37416_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _37416_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _37416_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _37416_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _37415_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _37415_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _37415_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _37415_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _37415_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _37415_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _37415_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _37415_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _37414_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _37414_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _37414_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _37414_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _37414_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _37414_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _37414_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _37414_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _37347_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _37347_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _37347_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _37347_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _37347_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _37347_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _37347_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _37347_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _37346_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _37346_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _37346_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _37346_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _37346_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _37346_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _37346_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _37346_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _37345_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _37345_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _37345_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _37345_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _37345_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _37345_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _37345_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _37345_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _37344_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _37344_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _37344_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _37344_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _37344_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _37344_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _37344_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _37344_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _37343_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _37343_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _37343_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _37343_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _37343_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _37343_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _37343_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _37343_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _37342_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _37342_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _37342_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _37342_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _37342_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _37342_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _37342_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _37342_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _37341_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _37341_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _37341_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _37341_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _37341_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _37341_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _37341_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _37341_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _37340_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _37340_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _37340_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _37340_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _37340_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _37340_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _37340_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _37340_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _37339_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _37339_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _37339_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _37339_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _37339_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _37339_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _37339_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _37339_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _37338_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _37338_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _37338_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _37338_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _37338_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _37338_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _37338_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _37338_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _37337_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _37337_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _37337_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _37337_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _37337_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _37337_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _37337_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _37337_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _37336_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _37336_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _37336_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _37336_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _37336_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _37336_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _37336_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _37336_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _37335_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _37335_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _37335_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _37335_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _37335_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _37335_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _37335_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _37335_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _37334_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _37334_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _37334_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _37334_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _37334_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _37334_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _37334_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _37334_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _37358_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _37358_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _37358_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _37358_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _37358_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _37358_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _37358_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _37358_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _37331_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _37331_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _37331_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _37331_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _37331_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _37331_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _37331_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _37331_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _37418_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _37418_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _37418_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _37418_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _37418_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _37418_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _37418_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _37418_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _37380_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _37380_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _37380_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _37380_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _37380_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _37380_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _37380_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _37380_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _37369_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _37369_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _37369_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _37369_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _37369_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _37369_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _37369_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _37369_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _37413_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _37413_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _37413_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _37413_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _37413_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _37413_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _37413_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _37413_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _37402_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _37402_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _37402_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _37402_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _37402_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _37402_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _37402_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _37402_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _37391_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _37391_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _37391_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _37391_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _37391_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _37391_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _37391_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _37391_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _37206_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _37206_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _37206_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _37206_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _37206_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _37206_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _37206_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _37206_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _37417_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _37417_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _37417_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _37417_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _37417_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _37417_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _37417_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _37417_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _37226_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _37226_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _37226_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _37226_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _37226_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _37226_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _37226_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _37226_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _37217_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _37217_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _37217_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _37217_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _37217_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _37217_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _37217_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _37217_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _37355_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _37355_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _37355_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _37355_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _37355_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _37355_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _37355_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _37355_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _37354_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _37354_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _37354_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _37354_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _37354_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _37354_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _37354_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _37354_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _37353_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _37353_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _37353_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _37353_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _37353_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _37353_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _37353_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _37353_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _37352_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _37352_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _37352_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _37352_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _37352_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _37352_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _37352_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _37352_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _37351_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _37351_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _37351_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _37351_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _37351_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _37351_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _37351_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _37351_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _37350_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _37350_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _37350_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _37350_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _37350_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _37350_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _37350_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _37350_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _37349_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _37349_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _37349_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _37349_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _37349_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _37349_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _37349_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _37349_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _37348_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _37348_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _37348_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _37348_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _37348_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _37348_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _37348_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _37348_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _37218_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _37218_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _37218_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _37218_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _37218_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _37218_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _37218_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _37218_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _37302_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _37302_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _37302_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _37302_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _37302_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _37302_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _37302_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _37302_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _37301_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _37301_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _37301_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _37301_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _37301_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _37301_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _37301_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _37301_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _37300_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _37300_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _37300_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _37300_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _37300_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _37300_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _37300_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _37300_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _37299_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _37299_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _37299_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _37299_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _37299_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _37299_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _37299_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _37299_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _37298_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _37298_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _37298_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _37298_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _37298_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _37298_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _37298_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _37298_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _37297_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _37297_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _37297_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _37297_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _37297_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _37297_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _37297_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _37297_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _37296_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _37296_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _37296_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _37296_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _37296_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _37296_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _37296_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _37296_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _37295_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _37295_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _37295_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _37295_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _37295_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _37295_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _37295_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _37295_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _37294_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _37294_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _37294_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _37294_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _37294_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _37294_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _37294_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _37294_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _37293_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _37293_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _37293_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _37293_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _37293_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _37293_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _37293_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _37293_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _37292_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _37292_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _37292_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _37292_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _37292_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _37292_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _37292_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _37292_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _37291_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _37291_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _37291_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _37291_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _37291_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _37291_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _37291_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _37291_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _37290_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _37290_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _37290_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _37290_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _37290_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _37290_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _37290_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _37290_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _37289_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _37289_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _37289_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _37289_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _37289_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _37289_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _37289_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _37289_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _37288_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _37288_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _37288_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _37288_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _37288_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _37288_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _37288_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _37288_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _37287_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _37287_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _37287_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _37287_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _37287_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _37287_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _37287_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _37287_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _37286_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _37286_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _37286_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _37286_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _37286_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _37286_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _37286_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _37286_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _37285_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _37285_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _37285_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _37285_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _37285_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _37285_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _37285_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _37285_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _37284_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _37284_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _37284_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _37284_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _37284_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _37284_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _37284_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _37284_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _37283_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _37283_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _37283_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _37283_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _37283_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _37283_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _37283_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _37283_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _37282_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _37282_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _37282_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _37282_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _37282_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _37282_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _37282_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _37282_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _37281_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _37281_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _37281_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _37281_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _37281_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _37281_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _37281_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _37281_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _37280_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _37280_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _37280_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _37280_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _37280_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _37280_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _37280_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _37280_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _37279_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _37279_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _37279_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _37279_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _37279_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _37279_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _37279_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _37279_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _37278_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _37278_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _37278_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _37278_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _37278_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _37278_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _37278_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _37278_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _37277_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _37277_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _37277_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _37277_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _37277_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _37277_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _37277_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _37277_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _37276_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _37276_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _37276_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _37276_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _37276_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _37276_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _37276_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _37276_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _37275_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _37275_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _37275_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _37275_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _37275_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _37275_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _37275_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _37275_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _37274_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _37274_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _37274_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _37274_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _37274_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _37274_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _37274_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _37274_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _37273_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _37273_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _37273_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _37273_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _37273_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _37273_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _37273_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _37273_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _37272_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _37272_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _37272_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _37272_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _37272_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _37272_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _37272_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _37272_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _37271_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _37271_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _37271_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _37271_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _37271_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _37271_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _37271_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _37271_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _37270_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _37270_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _37270_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _37270_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _37270_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _37270_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _37270_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _37270_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _37269_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _37269_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _37269_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _37269_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _37269_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _37269_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _37269_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _37269_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _37268_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _37268_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _37268_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _37268_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _37268_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _37268_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _37268_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _37268_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _37267_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _37267_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _37267_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _37267_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _37267_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _37267_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _37267_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _37267_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _37266_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _37266_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _37266_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _37266_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _37266_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _37266_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _37266_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _37266_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _37265_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _37265_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _37265_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _37265_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _37265_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _37265_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _37265_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _37265_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _37264_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _37264_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _37264_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _37264_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _37264_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _37264_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _37264_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _37264_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _37263_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _37263_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _37263_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _37263_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _37263_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _37263_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _37263_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _37263_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _37262_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _37262_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _37262_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _37262_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _37262_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _37262_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _37262_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _37262_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _37261_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _37261_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _37261_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _37261_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _37261_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _37261_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _37261_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _37261_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _37260_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _37260_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _37260_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _37260_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _37260_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _37260_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _37260_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _37260_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _37259_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _37259_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _37259_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _37259_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _37259_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _37259_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _37259_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _37259_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _37258_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _37258_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _37258_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _37258_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _37258_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _37258_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _37258_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _37258_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _37257_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _37257_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _37257_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _37257_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _37257_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _37257_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _37257_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _37257_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _37256_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _37256_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _37256_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _37256_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _37256_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _37256_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _37256_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _37256_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _37255_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _37255_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _37255_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _37255_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _37255_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _37255_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _37255_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _37255_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _37254_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _37254_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _37254_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _37254_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _37254_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _37254_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _37254_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _37254_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _37253_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _37253_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _37253_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _37253_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _37253_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _37253_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _37253_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _37253_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _37252_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _37252_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _37252_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _37252_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _37252_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _37252_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _37252_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _37252_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _37251_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _37251_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _37251_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _37251_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _37251_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _37251_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _37251_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _37251_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _37250_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _37250_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _37250_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _37250_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _37250_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _37250_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _37250_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _37250_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _37249_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _37249_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _37249_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _37249_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _37249_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _37249_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _37249_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _37249_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _37248_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _37248_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _37248_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _37248_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _37248_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _37248_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _37248_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _37248_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _37247_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _37247_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _37247_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _37247_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _37247_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _37247_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _37247_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _37247_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _37246_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _37246_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _37246_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _37246_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _37246_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _37246_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _37246_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _37246_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _37245_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _37245_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _37245_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _37245_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _37245_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _37245_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _37245_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _37245_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _37244_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _37244_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _37244_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _37244_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _37244_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _37244_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _37244_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _37244_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _37243_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _37243_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _37243_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _37243_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _37243_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _37243_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _37243_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _37243_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _37242_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _37242_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _37242_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _37242_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _37242_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _37242_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _37242_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _37242_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _37241_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _37241_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _37241_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _37241_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _37241_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _37241_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _37241_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _37241_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _37240_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _37240_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _37240_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _37240_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _37240_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _37240_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _37240_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _37240_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _37239_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _37239_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _37239_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _37239_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _37239_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _37239_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _37239_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _37239_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _37238_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _37238_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _37238_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _37238_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _37238_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _37238_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _37238_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _37238_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _37237_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _37237_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _37237_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _37237_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _37237_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _37237_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _37237_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _37237_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _37236_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _37236_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _37236_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _37236_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _37236_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _37236_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _37236_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _37236_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _37235_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _37235_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _37235_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _37235_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _37235_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _37235_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _37235_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _37235_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _37234_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _37234_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _37234_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _37234_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _37234_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _37234_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _37234_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _37234_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _37233_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _37233_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _37233_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _37233_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _37233_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _37233_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _37233_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _37233_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _37232_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _37232_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _37232_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _37232_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _37232_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _37232_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _37232_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _37232_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _37231_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _37231_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _37231_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _37231_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _37231_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _37231_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _37231_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _37231_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _37230_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _37230_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _37230_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _37230_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _37230_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _37230_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _37230_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _37230_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _37229_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _37229_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _37229_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _37229_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _37229_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _37229_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _37229_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _37229_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _37228_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _37228_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _37228_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _37228_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _37228_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _37228_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _37228_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _37228_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _37227_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _37227_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _37227_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _37227_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _37227_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _37227_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _37227_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _37227_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _37225_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _37225_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _37225_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _37225_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _37225_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _37225_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _37225_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _37225_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _37224_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _37224_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _37224_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _37224_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _37224_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _37224_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _37224_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _37224_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _37223_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _37223_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _37223_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _37223_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _37223_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _37223_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _37223_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _37223_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _37222_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _37222_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _37222_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _37222_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _37222_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _37222_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _37222_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _37222_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _37221_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _37221_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _37221_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _37221_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _37221_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _37221_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _37221_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _37221_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _37220_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _37220_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _37220_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _37220_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _37220_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _37220_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _37220_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _37220_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _37219_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _37219_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _37219_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _37219_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _37219_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _37219_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _37219_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _37219_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _37333_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _37333_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _37333_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _37333_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _37333_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _37333_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _37333_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _37333_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _37332_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _37332_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _37332_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _37332_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _37332_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _37332_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _37332_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _37332_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _37215_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _37215_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _37215_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _37215_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _37215_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _37215_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _37215_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _37215_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _37214_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _37214_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _37214_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _37214_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _37214_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _37214_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _37214_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _37214_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _37213_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _37213_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _37213_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _37213_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _37213_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _37213_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _37213_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _37213_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _37212_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _37212_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _37212_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _37212_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _37212_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _37212_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _37212_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _37212_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _37211_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _37211_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _37211_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _37211_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _37211_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _37211_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _37211_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _37211_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _37210_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _37210_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _37210_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _37210_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _37210_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _37210_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _37210_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _37210_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _37209_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _37209_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _37209_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _37209_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _37209_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _37209_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _37209_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _37209_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _37208_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _37208_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _37208_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _37208_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _37208_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _37208_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _37208_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _37208_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _37207_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _37207_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _37207_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _37207_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _37207_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _37207_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _37207_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _37207_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _37205_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _37205_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _37205_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _37205_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _37205_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _37205_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _37205_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _37205_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _37204_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _37204_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _37204_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _37204_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _37204_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _37204_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _37204_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _37204_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _37203_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _37203_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _37203_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _37203_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _37203_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _37203_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _37203_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _37203_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _37202_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _37202_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _37202_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _37202_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _37202_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _37202_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _37202_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _37202_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _37201_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _37201_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _37201_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _37201_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _37201_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _37201_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _37201_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _37201_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _37200_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _37200_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _37200_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _37200_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _37200_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _37200_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _37200_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _37200_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _37199_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _37199_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _37199_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _37199_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _37199_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _37199_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _37199_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _37199_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _37198_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _37198_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _37198_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _37198_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _37198_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _37198_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _37198_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _37198_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _37197_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _37197_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _37197_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _37197_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _37197_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _37197_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _37197_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _37197_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _37196_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _37196_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _37196_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _37196_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _37196_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _37196_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _37196_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _37196_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _37194_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _37194_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _37194_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _37194_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _37194_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _37194_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _37194_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _37194_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _37193_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _37193_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _37193_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _37193_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _37193_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _37193_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _37193_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _37193_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _37192_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _37192_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _37192_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _37192_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _37192_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _37192_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _37192_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _37192_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _37191_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _37191_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _37191_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _37191_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _37191_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _37191_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _37191_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _37191_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _37190_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _37190_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _37190_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _37190_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _37190_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _37190_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _37190_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _37190_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _37189_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _37189_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _37189_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _37189_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _37189_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _37189_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _37189_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _37189_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _37188_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _37188_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _37188_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _37188_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _37188_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _37188_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _37188_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _37188_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _37187_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _37187_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _37187_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _37187_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _37187_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _37187_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _37187_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _37187_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _37186_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _37186_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _37186_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _37186_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _37186_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _37186_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _37186_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _37186_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _37185_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _37185_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _37185_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _37185_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _37185_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _37185_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _37185_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _37185_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _37183_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _37183_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _37183_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _37183_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _37183_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _37183_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _37183_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _37183_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _37182_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _37182_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _37182_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _37182_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _37182_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _37182_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _37182_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _37182_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _37181_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _37181_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _37181_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _37181_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _37181_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _37181_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _37181_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _37181_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _37180_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _37180_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _37180_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _37180_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _37180_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _37180_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _37180_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _37180_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _37179_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _37179_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _37179_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _37179_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _37179_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _37179_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _37179_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _37179_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _37178_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _37178_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _37178_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _37178_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _37178_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _37178_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _37178_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _37178_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _37177_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _37177_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _37177_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _37177_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _37177_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _37177_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _37177_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _37177_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _37176_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _37176_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _37176_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _37176_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _37176_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _37176_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _37176_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _37176_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _37175_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _37175_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _37175_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _37175_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _37175_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _37175_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _37175_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _37175_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _37174_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _37174_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _37174_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _37174_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _37174_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _37174_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _37174_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _37174_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _37172_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _37172_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _37172_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _37172_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _37172_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _37172_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _37172_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _37172_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _37171_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _37171_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _37171_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _37171_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _37171_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _37171_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _37171_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _37171_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _37170_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _37170_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _37170_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _37170_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _37170_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _37170_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _37170_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _37170_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _37169_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _37169_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _37169_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _37169_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _37169_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _37169_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _37169_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _37169_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _37168_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _37168_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _37168_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _37168_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _37168_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _37168_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _37168_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _37168_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _37167_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _37167_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _37167_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _37167_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _37167_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _37167_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _37167_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _37167_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _37166_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _37166_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _37166_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _37166_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _37166_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _37166_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _37166_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _37166_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _37165_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _37165_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _37165_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _37165_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _37165_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _37165_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _37165_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _37165_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _37164_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _37164_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _37164_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _37164_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _37164_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _37164_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _37164_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _37164_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _37163_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _37163_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _37163_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _37163_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _37163_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _37163_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _37163_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _37163_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _37329_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _37329_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _37329_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _37329_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _37329_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _37329_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _37329_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _37329_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _37328_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _37328_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _37328_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _37328_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _37328_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _37328_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _37328_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _37328_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _37327_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _37327_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _37327_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _37327_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _37327_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _37327_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _37327_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _37327_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _37326_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _37326_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _37326_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _37326_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _37326_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _37326_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _37326_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _37326_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _37325_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _37325_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _37325_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _37325_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _37325_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _37325_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _37325_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _37325_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _37324_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _37324_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _37324_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _37324_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _37324_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _37324_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _37324_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _37324_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _37323_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _37323_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _37323_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _37323_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _37323_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _37323_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _37323_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _37323_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _37322_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _37322_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _37322_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _37322_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _37322_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _37322_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _37322_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _37322_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _37321_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _37321_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _37321_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _37321_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _37321_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _37321_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _37321_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _37321_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _37320_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _37320_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _37320_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _37320_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _37320_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _37320_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _37320_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _37320_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _37319_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _37319_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _37319_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _37319_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _37319_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _37319_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _37319_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _37319_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _37318_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _37318_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _37318_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _37318_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _37318_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _37318_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _37318_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _37318_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _37317_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _37317_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _37317_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _37317_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _37317_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _37317_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _37317_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _37317_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _37316_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _37316_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _37316_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _37316_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _37316_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _37316_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _37316_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _37316_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _37315_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _37315_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _37315_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _37315_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _37315_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _37315_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _37315_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _37315_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _37314_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _37314_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _37314_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _37314_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _37314_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _37314_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _37314_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _37314_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _37313_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _37313_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _37313_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _37313_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _37313_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _37313_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _37313_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _37313_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _37312_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _37312_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _37312_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _37312_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _37312_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _37312_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _37312_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _37312_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _37311_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _37311_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _37311_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _37311_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _37311_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _37311_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _37311_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _37311_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _37310_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _37310_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _37310_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _37310_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _37310_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _37310_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _37310_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _37310_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _37309_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _37309_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _37309_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _37309_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _37309_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _37309_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _37309_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _37309_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _37308_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _37308_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _37308_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _37308_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _37308_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _37308_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _37308_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _37308_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _37307_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _37307_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _37307_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _37307_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _37307_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _37307_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _37307_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _37307_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _37306_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _37306_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _37306_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _37306_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _37306_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _37306_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _37306_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _37306_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _37305_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _37305_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _37305_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _37305_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _37305_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _37305_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _37305_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _37305_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _37304_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _37304_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _37304_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _37304_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _37304_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _37304_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _37304_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _37304_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _37356_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _37356_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _37356_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _37356_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _37356_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _37356_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _37356_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _37356_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _37216_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _37216_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _37216_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _37216_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _37216_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _37216_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _37216_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _37216_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _37195_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _37195_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _37195_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _37195_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _37195_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _37195_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _37195_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _37195_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _37184_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _37184_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _37184_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _37184_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _37184_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _37184_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _37184_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _37184_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _37173_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _37173_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _37173_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _37173_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _37173_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _37173_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _37173_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _37173_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _37330_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _37330_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _37330_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _37330_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _37330_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _37330_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _37330_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _37330_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _32679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _32678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _32677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _32676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _32675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _32673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _32674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _32744_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , _33297_);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _33282_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _33287_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _33288_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _33289_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _33283_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _33284_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _33285_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _33290_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _33291_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _33292_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _33293_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _33294_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _33295_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _33296_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _33286_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _32956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _32957_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _32958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _32959_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _32960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _32961_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _32962_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _32955_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _32954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _32953_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _32952_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _32951_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _32950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _32949_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _32948_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _32947_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _32721_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _32727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _32728_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _32734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _32733_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _32732_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _32731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _32720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _32730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _32729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _32726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _32725_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _32724_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _32723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _32722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _32719_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _32795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _32791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _32790_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _32808_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _32806_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _32807_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _32811_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _32816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _32815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _32812_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _32792_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _32810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _32793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _32794_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _32809_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _32805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _32796_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _32804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _32813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _32797_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _32814_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _32834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _32798_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _32799_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _32800_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _32801_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _32833_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _32832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _32831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _32802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _32830_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _32829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _32828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _32827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _32826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _32825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _32824_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _32803_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _32823_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _32821_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _32822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _32820_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _32819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _32818_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _32817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _33281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _32707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _32704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _32706_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _32705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _32703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _32688_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _32689_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _32686_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _32691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _32690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _32692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _32694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _32693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _32696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _32695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _32687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _32700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _32701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _32702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _32685_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _32684_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _32683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _32682_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _32680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _32711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _32710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _32709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _32708_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _32699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _32698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _32697_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _32681_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _32718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _32717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _32716_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _32715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _32714_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _32713_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _32712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _32736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _32737_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _32738_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _32739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _32740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _32741_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _32742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _32743_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _32735_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _32748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _32749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _32755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _32756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _32757_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _32758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _32759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _32760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _32761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _32750_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _32762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _32763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _32764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _32765_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _32766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _32767_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _32768_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _32751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _32752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _32753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _32769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _32770_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _32771_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _32772_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _32773_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _32774_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _32775_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _32754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _32776_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _32777_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _32778_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _32779_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _32780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _32781_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _32782_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _32746_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _32745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _32783_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _32784_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _32785_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _32786_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _32787_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _32788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _32789_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _32747_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _32902_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _32903_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _32907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _32901_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _32926_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _32927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _32929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _32936_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _32937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _32938_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _32939_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _32904_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _32940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _32941_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _32942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _32943_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _32944_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _32945_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _32946_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _32905_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _32906_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _32912_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _32913_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _32914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _32915_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _32916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _32917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _32918_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _32908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _32919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _32920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _32921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _32922_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _32923_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _32924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _32925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _32909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _32910_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _32928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _32930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _32931_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _32932_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _32933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _32934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _32935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _32911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _32858_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _32843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _32840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _32839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _32838_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _32887_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _32850_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _32891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _32888_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _32900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _32857_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _32893_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _32894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _32846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _32856_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _32855_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _32854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _32849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _32842_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _32847_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _32866_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _32886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _32863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _32864_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _32865_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _32874_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _32875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _32878_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _32884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _32885_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _32835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _32836_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _32837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _32841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _32844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _32892_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _32897_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _32899_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _32848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _32845_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _32859_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _32860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _32861_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _32862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _32867_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _32868_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _32869_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _32870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _32871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _32851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _32872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _32873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _32876_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _32877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _32879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _32880_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _32881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _32852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _32882_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _32883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _32889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _32890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _32895_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _32896_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _32898_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _32853_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rmw , \oc8051_top_1.oc8051_decoder1.rmw );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.bank_sel [0], \oc8051_top_1.oc8051_memory_interface1.rn [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.bank_sel [1], \oc8051_top_1.oc8051_memory_interface1.rn [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_sfr [0], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_sfr [1], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [0], \oc8051_top_1.oc8051_memory_interface1.des_acc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [1], \oc8051_top_1.oc8051_memory_interface1.des_acc [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [2], \oc8051_top_1.oc8051_memory_interface1.des_acc [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [3], \oc8051_top_1.oc8051_memory_interface1.des_acc [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [4], \oc8051_top_1.oc8051_memory_interface1.des_acc [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [5], \oc8051_top_1.oc8051_memory_interface1.des_acc [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [6], \oc8051_top_1.oc8051_memory_interface1.des_acc [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [7], \oc8051_top_1.oc8051_memory_interface1.des_acc [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [0], \oc8051_top_1.oc8051_memory_interface1.des2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [1], \oc8051_top_1.oc8051_memory_interface1.des2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [2], \oc8051_top_1.oc8051_memory_interface1.des2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [3], \oc8051_top_1.oc8051_memory_interface1.des2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [4], \oc8051_top_1.oc8051_memory_interface1.des2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [5], \oc8051_top_1.oc8051_memory_interface1.des2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [6], \oc8051_top_1.oc8051_memory_interface1.des2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [7], \oc8051_top_1.oc8051_memory_interface1.des2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_rd_sel [0], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_rd_sel [1], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_rd_sel [2], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [0], \oc8051_top_1.oc8051_memory_interface1.sp [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [1], \oc8051_top_1.oc8051_memory_interface1.sp [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [2], \oc8051_top_1.oc8051_memory_interface1.sp [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [3], \oc8051_top_1.oc8051_memory_interface1.sp [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [4], \oc8051_top_1.oc8051_memory_interface1.sp [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [5], \oc8051_top_1.oc8051_memory_interface1.sp [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [6], \oc8051_top_1.oc8051_memory_interface1.sp [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_out [7], \oc8051_top_1.oc8051_memory_interface1.sp [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.bit_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.bit_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [0], \oc8051_top_1.oc8051_memory_interface1.des_acc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [1], \oc8051_top_1.oc8051_memory_interface1.des_acc [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [2], \oc8051_top_1.oc8051_memory_interface1.des_acc [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [3], \oc8051_top_1.oc8051_memory_interface1.des_acc [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [4], \oc8051_top_1.oc8051_memory_interface1.des_acc [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [5], \oc8051_top_1.oc8051_memory_interface1.des_acc [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [6], \oc8051_top_1.oc8051_memory_interface1.des_acc [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [7], \oc8051_top_1.oc8051_memory_interface1.des_acc [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_sfr [0], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_sfr [1], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [0], \oc8051_top_1.oc8051_memory_interface1.des_acc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [1], \oc8051_top_1.oc8051_memory_interface1.des_acc [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [2], \oc8051_top_1.oc8051_memory_interface1.des_acc [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [3], \oc8051_top_1.oc8051_memory_interface1.des_acc [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [4], \oc8051_top_1.oc8051_memory_interface1.des_acc [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [5], \oc8051_top_1.oc8051_memory_interface1.des_acc [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [6], \oc8051_top_1.oc8051_memory_interface1.des_acc [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [7], \oc8051_top_1.oc8051_memory_interface1.des_acc [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [0], \oc8051_top_1.oc8051_memory_interface1.des2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [1], \oc8051_top_1.oc8051_memory_interface1.des2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [2], \oc8051_top_1.oc8051_memory_interface1.des2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [3], \oc8051_top_1.oc8051_memory_interface1.des2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [4], \oc8051_top_1.oc8051_memory_interface1.des2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [5], \oc8051_top_1.oc8051_memory_interface1.des2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [6], \oc8051_top_1.oc8051_memory_interface1.des2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [7], \oc8051_top_1.oc8051_memory_interface1.des2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.enable , \oc8051_top_1.oc8051_alu1.enable_mul );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src1 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [6]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.src2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 [11], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 [12], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 [13], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 [14], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result1 [15], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [2], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [3], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [4], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [5], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [6], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [6]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [7], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [8], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [9], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [10], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [11], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [12], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [13], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [14], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.mul_result [15], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.shifted [0], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.shifted [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.enable , \oc8051_top_1.oc8051_alu1.enable_div );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem0 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [14], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [15], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [0], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [6]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [8], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [9], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [8]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [10], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [9]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [11], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [10]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [12], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [11]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [13], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [12]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [14], \oc8051_top_1.oc8051_alu1.oc8051_div1.cmp0 [13]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.cmp1 [15], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rem_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcCy , \oc8051_top_1.oc8051_cy_select1.data_out );
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.bit_in , \oc8051_top_1.oc8051_cy_select1.data_in );
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.op_code [0], \oc8051_top_1.oc8051_decoder1.alu_op_o [0]);
  buf(\oc8051_top_1.oc8051_alu1.op_code [1], \oc8051_top_1.oc8051_decoder1.alu_op_o [1]);
  buf(\oc8051_top_1.oc8051_alu1.op_code [2], \oc8051_top_1.oc8051_decoder1.alu_op_o [2]);
  buf(\oc8051_top_1.oc8051_alu1.op_code [3], \oc8051_top_1.oc8051_decoder1.alu_op_o [3]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.src1 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [2]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [3]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [4]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [5]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [6]);
  buf(\oc8051_top_1.oc8051_alu1.src2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [0], \oc8051_top_1.oc8051_alu_src_sel1.src3 [0]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [1], \oc8051_top_1.oc8051_alu_src_sel1.src3 [1]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [2], \oc8051_top_1.oc8051_alu_src_sel1.src3 [2]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [3], \oc8051_top_1.oc8051_alu_src_sel1.src3 [3]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [4], \oc8051_top_1.oc8051_alu_src_sel1.src3 [4]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [5], \oc8051_top_1.oc8051_alu_src_sel1.src3 [5]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [6], \oc8051_top_1.oc8051_alu_src_sel1.src3 [6]);
  buf(\oc8051_top_1.oc8051_alu1.src3 [7], \oc8051_top_1.oc8051_alu_src_sel1.src3 [7]);
  buf(\oc8051_top_1.oc8051_alu1.desCy , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_alu1.desAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in );
  buf(\oc8051_top_1.oc8051_alu1.desOv , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in );
  buf(\oc8051_top_1.oc8051_alu1.des1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_alu1.des1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_alu1.des1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_alu1.des1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_alu1.des1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_alu1.des1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_alu1.des1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_alu1.des1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [0], \oc8051_top_1.oc8051_memory_interface1.des2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [1], \oc8051_top_1.oc8051_memory_interface1.des2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [2], \oc8051_top_1.oc8051_memory_interface1.des2 [2]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [3], \oc8051_top_1.oc8051_memory_interface1.des2 [3]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [4], \oc8051_top_1.oc8051_memory_interface1.des2 [4]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [5], \oc8051_top_1.oc8051_memory_interface1.des2 [5]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [6], \oc8051_top_1.oc8051_memory_interface1.des2 [6]);
  buf(\oc8051_top_1.oc8051_alu1.des2 [7], \oc8051_top_1.oc8051_memory_interface1.des2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [0], \oc8051_top_1.oc8051_memory_interface1.des_acc [0]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [1], \oc8051_top_1.oc8051_memory_interface1.des_acc [1]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [2], \oc8051_top_1.oc8051_memory_interface1.des_acc [2]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [3], \oc8051_top_1.oc8051_memory_interface1.des_acc [3]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [4], \oc8051_top_1.oc8051_memory_interface1.des_acc [4]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [5], \oc8051_top_1.oc8051_memory_interface1.des_acc [5]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [6], \oc8051_top_1.oc8051_memory_interface1.des_acc [6]);
  buf(\oc8051_top_1.oc8051_alu1.des_acc [7], \oc8051_top_1.oc8051_memory_interface1.des_acc [7]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [0], \oc8051_top_1.oc8051_comp1.des [0]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [1], \oc8051_top_1.oc8051_comp1.des [1]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [2], \oc8051_top_1.oc8051_comp1.des [2]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [3], \oc8051_top_1.oc8051_comp1.des [3]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [4], \oc8051_top_1.oc8051_comp1.des [4]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [5], \oc8051_top_1.oc8051_comp1.des [5]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [6], \oc8051_top_1.oc8051_comp1.des [6]);
  buf(\oc8051_top_1.oc8051_alu1.sub_result [7], \oc8051_top_1.oc8051_comp1.des [7]);
  buf(\oc8051_top_1.oc8051_alu1.add1 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.add1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.add1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.add1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.add1 [4], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.add2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.add2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [2]);
  buf(\oc8051_top_1.oc8051_alu1.add2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [3]);
  buf(\oc8051_top_1.oc8051_alu1.add2 [4], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add3 [0], \oc8051_top_1.oc8051_cy_select1.data_out );
  buf(\oc8051_top_1.oc8051_alu1.add3 [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add3 [2], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add3 [3], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add3 [4], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add4 [4], \oc8051_top_1.oc8051_alu1.add7 [0]);
  buf(\oc8051_top_1.oc8051_alu1.add5 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.add5 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.add5 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.add5 [3], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add6 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [4]);
  buf(\oc8051_top_1.oc8051_alu1.add6 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [5]);
  buf(\oc8051_top_1.oc8051_alu1.add6 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [6]);
  buf(\oc8051_top_1.oc8051_alu1.add6 [3], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add7 [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add7 [2], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add7 [3], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.add9 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.add9 [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.adda [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.adda [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.addb [0], \oc8051_top_1.oc8051_alu1.add8 [3]);
  buf(\oc8051_top_1.oc8051_alu1.addb [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub1 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.sub1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.sub1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.sub1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.sub1 [4], 1'b1);
  buf(\oc8051_top_1.oc8051_alu1.sub2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.sub2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.sub2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [2]);
  buf(\oc8051_top_1.oc8051_alu1.sub2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [3]);
  buf(\oc8051_top_1.oc8051_alu1.sub2 [4], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub3 [0], \oc8051_top_1.oc8051_cy_select1.data_out );
  buf(\oc8051_top_1.oc8051_alu1.sub3 [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub3 [2], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub3 [3], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub3 [4], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub4 [0], \oc8051_top_1.oc8051_comp1.des [0]);
  buf(\oc8051_top_1.oc8051_alu1.sub4 [1], \oc8051_top_1.oc8051_comp1.des [1]);
  buf(\oc8051_top_1.oc8051_alu1.sub4 [2], \oc8051_top_1.oc8051_comp1.des [2]);
  buf(\oc8051_top_1.oc8051_alu1.sub4 [3], \oc8051_top_1.oc8051_comp1.des [3]);
  buf(\oc8051_top_1.oc8051_alu1.sub5 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.sub5 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.sub5 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.sub5 [3], 1'b1);
  buf(\oc8051_top_1.oc8051_alu1.sub6 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [4]);
  buf(\oc8051_top_1.oc8051_alu1.sub6 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [5]);
  buf(\oc8051_top_1.oc8051_alu1.sub6 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [6]);
  buf(\oc8051_top_1.oc8051_alu1.sub6 [3], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub7 [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub7 [2], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub7 [3], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.sub8 [0], \oc8051_top_1.oc8051_comp1.des [4]);
  buf(\oc8051_top_1.oc8051_alu1.sub8 [1], \oc8051_top_1.oc8051_comp1.des [5]);
  buf(\oc8051_top_1.oc8051_alu1.sub8 [2], \oc8051_top_1.oc8051_comp1.des [6]);
  buf(\oc8051_top_1.oc8051_alu1.sub9 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.sub9 [1], 1'b1);
  buf(\oc8051_top_1.oc8051_alu1.suba [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.suba [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.subb [1], 1'b0);
  buf(\oc8051_top_1.oc8051_alu1.subc [0], \oc8051_top_1.oc8051_comp1.des [7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [2], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [3], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [4], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [5], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [6], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [7], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_mul1.des2 [7]);
  buf(\oc8051_top_1.oc8051_alu1.mulOv , \oc8051_top_1.oc8051_alu1.oc8051_mul1.desOv );
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [5]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [6]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.des1 [7]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.divOv , \oc8051_top_1.oc8051_alu1.oc8051_div1.desOv );
  buf(\oc8051_top_1.oc8051_alu1.dec [0], \oc8051_top_1.oc8051_alu1.inc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rd , \oc8051_top_1.oc8051_decoder1.rd );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [0], \oc8051_top_1.oc8051_memory_interface1.iram_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [1], \oc8051_top_1.oc8051_memory_interface1.iram_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [2], \oc8051_top_1.oc8051_memory_interface1.iram_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [3], \oc8051_top_1.oc8051_memory_interface1.iram_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [4], \oc8051_top_1.oc8051_memory_interface1.iram_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [5], \oc8051_top_1.oc8051_memory_interface1.iram_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [6], \oc8051_top_1.oc8051_memory_interface1.iram_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.ram [7], \oc8051_top_1.oc8051_memory_interface1.iram_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [0], \oc8051_top_1.oc8051_decoder1.op_in [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [1], \oc8051_top_1.oc8051_decoder1.op_in [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [2], \oc8051_top_1.oc8051_decoder1.op_in [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [3], \oc8051_top_1.oc8051_decoder1.op_in [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [4], \oc8051_top_1.oc8051_decoder1.op_in [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [5], \oc8051_top_1.oc8051_decoder1.op_in [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [6], \oc8051_top_1.oc8051_decoder1.op_in [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op1 [7], \oc8051_top_1.oc8051_decoder1.op_in [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [0], \oc8051_top_1.oc8051_memory_interface1.op2_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [1], \oc8051_top_1.oc8051_memory_interface1.op2_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [2], \oc8051_top_1.oc8051_memory_interface1.op2_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [3], \oc8051_top_1.oc8051_memory_interface1.op2_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [4], \oc8051_top_1.oc8051_memory_interface1.op2_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [5], \oc8051_top_1.oc8051_memory_interface1.op2_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [6], \oc8051_top_1.oc8051_memory_interface1.op2_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2 [7], \oc8051_top_1.oc8051_memory_interface1.op2_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [0], \oc8051_top_1.oc8051_memory_interface1.op3_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [1], \oc8051_top_1.oc8051_memory_interface1.op3_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [2], \oc8051_top_1.oc8051_memory_interface1.op3_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [3], \oc8051_top_1.oc8051_memory_interface1.op3_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [4], \oc8051_top_1.oc8051_memory_interface1.op3_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [5], \oc8051_top_1.oc8051_memory_interface1.op3_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [6], \oc8051_top_1.oc8051_memory_interface1.op3_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3 [7], \oc8051_top_1.oc8051_memory_interface1.op3_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src1 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.src2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.wr_o , \oc8051_top_1.wr_o );
  buf(\oc8051_top_1.oc8051_decoder1.pc_wr , \oc8051_top_1.pc_wr );
  buf(\oc8051_top_1.oc8051_decoder1.op1_c [0], \oc8051_top_1.oc8051_decoder1.op_cur [0]);
  buf(\oc8051_top_1.oc8051_decoder1.op1_c [1], \oc8051_top_1.oc8051_decoder1.op_cur [1]);
  buf(\oc8051_top_1.oc8051_decoder1.op1_c [2], \oc8051_top_1.oc8051_decoder1.op_cur [2]);
  buf(\oc8051_top_1.oc8051_comp1.sel [0], \oc8051_top_1.oc8051_decoder1.comp_sel [0]);
  buf(\oc8051_top_1.oc8051_comp1.sel [1], \oc8051_top_1.oc8051_decoder1.comp_sel [1]);
  buf(\oc8051_top_1.oc8051_comp1.b_in , \oc8051_top_1.oc8051_cy_select1.data_in );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_comp1.eq , \oc8051_top_1.oc8051_decoder1.eq );
  buf(\oc8051_top_1.oc8051_comp1.eq_r , \oc8051_top_1.oc8051_decoder1.eq );
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_i , \oc8051_top_1.wr_o );
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_bit_i , \oc8051_top_1.oc8051_decoder1.bit_addr );
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [2], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [3], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [4], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [5], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [6], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sp_w [7], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_out , \oc8051_top_1.oc8051_cy_select1.data_in );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_wait , \oc8051_top_1.oc8051_decoder1.mem_wait );
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_o , \oc8051_top_1.wr_o );
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_bit_o , \oc8051_top_1.oc8051_decoder1.bit_addr );
  buf(\oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff );
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [4], cxrom_addr[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [5], cxrom_addr[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [6], cxrom_addr[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [7], cxrom_addr[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [8], cxrom_addr[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [9], cxrom_addr[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [10], cxrom_addr[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [11], cxrom_addr[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [12], cxrom_addr[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [13], cxrom_addr[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [14], cxrom_addr[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.iadr_o [15], cxrom_addr[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_rom_sel , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_sel [0], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_sel [1], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_sel [2], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rn [0], \oc8051_top_1.oc8051_decoder1.op_cur [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rn [1], \oc8051_top_1.oc8051_decoder1.op_cur [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rn [2], \oc8051_top_1.oc8051_decoder1.op_cur [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [0], \oc8051_top_1.oc8051_ram_top1.rd_addr [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [1], \oc8051_top_1.oc8051_ram_top1.rd_addr [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [2], \oc8051_top_1.oc8051_ram_top1.rd_addr [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [3], \oc8051_top_1.oc8051_ram_top1.rd_addr [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [4], \oc8051_top_1.oc8051_ram_top1.rd_addr [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [5], \oc8051_top_1.oc8051_ram_top1.rd_addr [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [6], \oc8051_top_1.oc8051_ram_top1.rd_addr [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rd_addr [7], \oc8051_top_1.oc8051_ram_top1.rd_addr [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [0], \oc8051_top_1.oc8051_memory_interface1.op2_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [1], \oc8051_top_1.oc8051_memory_interface1.op2_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [2], \oc8051_top_1.oc8051_memory_interface1.op2_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [3], \oc8051_top_1.oc8051_memory_interface1.op2_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [4], \oc8051_top_1.oc8051_memory_interface1.op2_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [5], \oc8051_top_1.oc8051_memory_interface1.op2_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [6], \oc8051_top_1.oc8051_memory_interface1.op2_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm [7], \oc8051_top_1.oc8051_memory_interface1.op2_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [0], \oc8051_top_1.oc8051_memory_interface1.op3_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [1], \oc8051_top_1.oc8051_memory_interface1.op3_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [2], \oc8051_top_1.oc8051_memory_interface1.op3_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [3], \oc8051_top_1.oc8051_memory_interface1.op3_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [4], \oc8051_top_1.oc8051_memory_interface1.op3_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [5], \oc8051_top_1.oc8051_memory_interface1.op3_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [6], \oc8051_top_1.oc8051_memory_interface1.op3_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2 [7], \oc8051_top_1.oc8051_memory_interface1.op3_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.intr , \oc8051_top_1.oc8051_sfr1.oc8051_int1.intr );
  buf(\oc8051_top_1.oc8051_memory_interface1.rd , \oc8051_top_1.oc8051_decoder1.rd );
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [0], \oc8051_top_1.oc8051_decoder1.op_in [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [1], \oc8051_top_1.oc8051_decoder1.op_in [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [2], \oc8051_top_1.oc8051_decoder1.op_in [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [3], \oc8051_top_1.oc8051_decoder1.op_in [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [4], \oc8051_top_1.oc8051_decoder1.op_in [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [5], \oc8051_top_1.oc8051_decoder1.op_in [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [6], \oc8051_top_1.oc8051_decoder1.op_in [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op1_out [7], \oc8051_top_1.oc8051_decoder1.op_in [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_wr_sel [0], \oc8051_top_1.oc8051_decoder1.pc_sel [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_wr_sel [1], \oc8051_top_1.oc8051_decoder1.pc_sel [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_wr_sel [2], \oc8051_top_1.oc8051_decoder1.pc_sel [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [0], \oc8051_top_1.oc8051_memory_interface1.des_acc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [1], \oc8051_top_1.oc8051_memory_interface1.des_acc [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [2], \oc8051_top_1.oc8051_memory_interface1.des_acc [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [3], \oc8051_top_1.oc8051_memory_interface1.des_acc [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [4], \oc8051_top_1.oc8051_memory_interface1.des_acc [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [5], \oc8051_top_1.oc8051_memory_interface1.des_acc [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [6], \oc8051_top_1.oc8051_memory_interface1.des_acc [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [7], \oc8051_top_1.oc8051_memory_interface1.des_acc [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [8], \oc8051_top_1.oc8051_memory_interface1.des2 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [9], \oc8051_top_1.oc8051_memory_interface1.des2 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [10], \oc8051_top_1.oc8051_memory_interface1.des2 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [11], \oc8051_top_1.oc8051_memory_interface1.des2 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [12], \oc8051_top_1.oc8051_memory_interface1.des2 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [13], \oc8051_top_1.oc8051_memory_interface1.des2 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [14], \oc8051_top_1.oc8051_memory_interface1.des2 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [15], \oc8051_top_1.oc8051_memory_interface1.des2 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.bank [0], \oc8051_top_1.oc8051_memory_interface1.rn [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.bank [1], \oc8051_top_1.oc8051_memory_interface1.rn [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.wr , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr );
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr , \oc8051_top_1.oc8051_decoder1.bit_addr );
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_data_out , \oc8051_top_1.oc8051_memory_interface1.bit_in );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [0], \oc8051_top_1.oc8051_memory_interface1.in_ram [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [1], \oc8051_top_1.oc8051_memory_interface1.in_ram [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [2], \oc8051_top_1.oc8051_memory_interface1.in_ram [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [3], \oc8051_top_1.oc8051_memory_interface1.in_ram [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [4], \oc8051_top_1.oc8051_memory_interface1.in_ram [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [5], \oc8051_top_1.oc8051_memory_interface1.in_ram [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [6], \oc8051_top_1.oc8051_memory_interface1.in_ram [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data [7], \oc8051_top_1.oc8051_memory_interface1.in_ram [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_data [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_addr_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_addr [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_addr_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr , \oc8051_top_1.wr_o );
  buf(\oc8051_top_1.oc8051_indi_addr1.sel , \oc8051_top_1.oc8051_decoder1.op_cur [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit , \oc8051_top_1.oc8051_decoder1.bit_addr );
  buf(\oc8051_top_1.oc8051_indi_addr1.bank [0], \oc8051_top_1.oc8051_memory_interface1.rn [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.bank [1], \oc8051_top_1.oc8051_memory_interface1.rn [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_addr [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [0], \oc8051_top_1.oc8051_memory_interface1.ri [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [1], \oc8051_top_1.oc8051_memory_interface1.ri [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [2], \oc8051_top_1.oc8051_memory_interface1.ri [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [3], \oc8051_top_1.oc8051_memory_interface1.ri [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [4], \oc8051_top_1.oc8051_memory_interface1.ri [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [5], \oc8051_top_1.oc8051_memory_interface1.ri [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [6], \oc8051_top_1.oc8051_memory_interface1.ri [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.ri_out [7], \oc8051_top_1.oc8051_memory_interface1.ri [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.we , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr );
  buf(\oc8051_top_1.oc8051_sfr1.bit_in , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.oc8051_sfr1.desAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in );
  buf(\oc8051_top_1.oc8051_sfr1.desOv , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in );
  buf(\oc8051_top_1.oc8051_sfr1.rmw , \oc8051_top_1.oc8051_decoder1.rmw );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit , \oc8051_top_1.oc8051_decoder1.bit_addr );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.wr_sfr [0], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [0]);
  buf(\oc8051_top_1.oc8051_sfr1.wr_sfr [1], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [1]);
  buf(\oc8051_top_1.oc8051_sfr1.comp_sel [0], \oc8051_top_1.oc8051_decoder1.comp_sel [0]);
  buf(\oc8051_top_1.oc8051_sfr1.comp_sel [1], \oc8051_top_1.oc8051_decoder1.comp_sel [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ram_rd_sel [0], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ram_rd_sel [1], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ram_rd_sel [2], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [2]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [0], \oc8051_top_1.oc8051_ram_top1.rd_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [1], \oc8051_top_1.oc8051_ram_top1.rd_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [2], \oc8051_top_1.oc8051_ram_top1.rd_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [3], \oc8051_top_1.oc8051_ram_top1.rd_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [4], \oc8051_top_1.oc8051_ram_top1.rd_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [5], \oc8051_top_1.oc8051_ram_top1.rd_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [6], \oc8051_top_1.oc8051_ram_top1.rd_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.adr0 [7], \oc8051_top_1.oc8051_ram_top1.rd_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.oc8051_sfr1.adr1 [7], \oc8051_top_1.wr_addr [7]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [0], \oc8051_top_1.oc8051_memory_interface1.des_acc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [1], \oc8051_top_1.oc8051_memory_interface1.des_acc [1]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [2], \oc8051_top_1.oc8051_memory_interface1.des_acc [2]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [3], \oc8051_top_1.oc8051_memory_interface1.des_acc [3]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [4], \oc8051_top_1.oc8051_memory_interface1.des_acc [4]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [5], \oc8051_top_1.oc8051_memory_interface1.des_acc [5]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [6], \oc8051_top_1.oc8051_memory_interface1.des_acc [6]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [7], \oc8051_top_1.oc8051_memory_interface1.des_acc [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [0], \oc8051_top_1.oc8051_memory_interface1.des2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [1], \oc8051_top_1.oc8051_memory_interface1.des2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [2], \oc8051_top_1.oc8051_memory_interface1.des2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [3], \oc8051_top_1.oc8051_memory_interface1.des2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [4], \oc8051_top_1.oc8051_memory_interface1.des2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [5], \oc8051_top_1.oc8051_memory_interface1.des2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [6], \oc8051_top_1.oc8051_memory_interface1.des2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [7], \oc8051_top_1.oc8051_memory_interface1.des2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.intr , \oc8051_top_1.oc8051_sfr1.oc8051_int1.intr );
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.comp_wait , \oc8051_top_1.comp_wait );
  buf(\oc8051_top_1.oc8051_sfr1.bank_sel [0], \oc8051_top_1.oc8051_memory_interface1.rn [3]);
  buf(\oc8051_top_1.oc8051_sfr1.bank_sel [1], \oc8051_top_1.oc8051_memory_interface1.rn [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [0], \oc8051_top_1.oc8051_memory_interface1.sp [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [1], \oc8051_top_1.oc8051_memory_interface1.sp [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [2], \oc8051_top_1.oc8051_memory_interface1.sp [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [3], \oc8051_top_1.oc8051_memory_interface1.sp [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [4], \oc8051_top_1.oc8051_memory_interface1.sp [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [5], \oc8051_top_1.oc8051_memory_interface1.sp [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [6], \oc8051_top_1.oc8051_memory_interface1.sp [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sp [7], \oc8051_top_1.oc8051_memory_interface1.sp [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [2], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [3], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [4], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [5], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [6], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sp_w [7], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_data [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_data [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_data [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_data [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.p , \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p );
  buf(\oc8051_top_1.oc8051_sfr1.uart_int , \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tc2_int , \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p );
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [0], \oc8051_top_1.oc8051_memory_interface1.iadr_o [0]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [1], \oc8051_top_1.oc8051_memory_interface1.iadr_o [1]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [2], \oc8051_top_1.oc8051_memory_interface1.iadr_o [2]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [3], \oc8051_top_1.oc8051_memory_interface1.iadr_o [3]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [4], cxrom_addr[4]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [5], cxrom_addr[5]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [6], cxrom_addr[6]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [7], cxrom_addr[7]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [8], cxrom_addr[8]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [9], cxrom_addr[9]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [10], cxrom_addr[10]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [11], cxrom_addr[11]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [12], cxrom_addr[12]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [13], cxrom_addr[13]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [14], cxrom_addr[14]);
  buf(\oc8051_symbolic_cxrom1.cxrom_addr [15], cxrom_addr[15]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.op_valid , op_valid);
  buf(\oc8051_symbolic_cxrom1.op_out [0], op_out[0]);
  buf(\oc8051_symbolic_cxrom1.op_out [1], op_out[1]);
  buf(\oc8051_symbolic_cxrom1.op_out [2], op_out[2]);
  buf(\oc8051_symbolic_cxrom1.op_out [3], op_out[3]);
  buf(\oc8051_symbolic_cxrom1.op_out [4], op_out[4]);
  buf(\oc8051_symbolic_cxrom1.op_out [5], op_out[5]);
  buf(\oc8051_symbolic_cxrom1.op_out [6], op_out[6]);
  buf(\oc8051_symbolic_cxrom1.op_out [7], op_out[7]);
  buf(\oc8051_symbolic_cxrom1.addr0 [0], \oc8051_top_1.oc8051_memory_interface1.iadr_o [0]);
  buf(\oc8051_symbolic_cxrom1.addr0 [1], \oc8051_top_1.oc8051_memory_interface1.iadr_o [1]);
  buf(\oc8051_symbolic_cxrom1.addr0 [2], \oc8051_top_1.oc8051_memory_interface1.iadr_o [2]);
  buf(\oc8051_symbolic_cxrom1.addr0 [3], \oc8051_top_1.oc8051_memory_interface1.iadr_o [3]);
  buf(\oc8051_symbolic_cxrom1.addr2 [0], \oc8051_top_1.oc8051_memory_interface1.iadr_o [0]);
  buf(\oc8051_symbolic_cxrom1.addr3 [0], \oc8051_symbolic_cxrom1.addr1 [0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc13 [0], \oc8051_symbolic_cxrom1.pc11 [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc23 [0], \oc8051_symbolic_cxrom1.pc21 [0]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.cxrom_addr [0], \oc8051_top_1.oc8051_memory_interface1.iadr_o [0]);
  buf(\oc8051_top_1.cxrom_addr [1], \oc8051_top_1.oc8051_memory_interface1.iadr_o [1]);
  buf(\oc8051_top_1.cxrom_addr [2], \oc8051_top_1.oc8051_memory_interface1.iadr_o [2]);
  buf(\oc8051_top_1.cxrom_addr [3], \oc8051_top_1.oc8051_memory_interface1.iadr_o [3]);
  buf(\oc8051_top_1.cxrom_addr [4], cxrom_addr[4]);
  buf(\oc8051_top_1.cxrom_addr [5], cxrom_addr[5]);
  buf(\oc8051_top_1.cxrom_addr [6], cxrom_addr[6]);
  buf(\oc8051_top_1.cxrom_addr [7], cxrom_addr[7]);
  buf(\oc8051_top_1.cxrom_addr [8], cxrom_addr[8]);
  buf(\oc8051_top_1.cxrom_addr [9], cxrom_addr[9]);
  buf(\oc8051_top_1.cxrom_addr [10], cxrom_addr[10]);
  buf(\oc8051_top_1.cxrom_addr [11], cxrom_addr[11]);
  buf(\oc8051_top_1.cxrom_addr [12], cxrom_addr[12]);
  buf(\oc8051_top_1.cxrom_addr [13], cxrom_addr[13]);
  buf(\oc8051_top_1.cxrom_addr [14], cxrom_addr[14]);
  buf(\oc8051_top_1.cxrom_addr [15], cxrom_addr[15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.ri [0], \oc8051_top_1.oc8051_memory_interface1.ri [0]);
  buf(\oc8051_top_1.ri [1], \oc8051_top_1.oc8051_memory_interface1.ri [1]);
  buf(\oc8051_top_1.ri [2], \oc8051_top_1.oc8051_memory_interface1.ri [2]);
  buf(\oc8051_top_1.ri [3], \oc8051_top_1.oc8051_memory_interface1.ri [3]);
  buf(\oc8051_top_1.ri [4], \oc8051_top_1.oc8051_memory_interface1.ri [4]);
  buf(\oc8051_top_1.ri [5], \oc8051_top_1.oc8051_memory_interface1.ri [5]);
  buf(\oc8051_top_1.ri [6], \oc8051_top_1.oc8051_memory_interface1.ri [6]);
  buf(\oc8051_top_1.ri [7], \oc8051_top_1.oc8051_memory_interface1.ri [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.sub_result [0], \oc8051_top_1.oc8051_comp1.des [0]);
  buf(\oc8051_top_1.sub_result [1], \oc8051_top_1.oc8051_comp1.des [1]);
  buf(\oc8051_top_1.sub_result [2], \oc8051_top_1.oc8051_comp1.des [2]);
  buf(\oc8051_top_1.sub_result [3], \oc8051_top_1.oc8051_comp1.des [3]);
  buf(\oc8051_top_1.sub_result [4], \oc8051_top_1.oc8051_comp1.des [4]);
  buf(\oc8051_top_1.sub_result [5], \oc8051_top_1.oc8051_comp1.des [5]);
  buf(\oc8051_top_1.sub_result [6], \oc8051_top_1.oc8051_comp1.des [6]);
  buf(\oc8051_top_1.sub_result [7], \oc8051_top_1.oc8051_comp1.des [7]);
  buf(\oc8051_top_1.iadr_o [0], \oc8051_top_1.oc8051_memory_interface1.iadr_o [0]);
  buf(\oc8051_top_1.iadr_o [1], \oc8051_top_1.oc8051_memory_interface1.iadr_o [1]);
  buf(\oc8051_top_1.iadr_o [2], \oc8051_top_1.oc8051_memory_interface1.iadr_o [2]);
  buf(\oc8051_top_1.iadr_o [3], \oc8051_top_1.oc8051_memory_interface1.iadr_o [3]);
  buf(\oc8051_top_1.iadr_o [4], cxrom_addr[4]);
  buf(\oc8051_top_1.iadr_o [5], cxrom_addr[5]);
  buf(\oc8051_top_1.iadr_o [6], cxrom_addr[6]);
  buf(\oc8051_top_1.iadr_o [7], cxrom_addr[7]);
  buf(\oc8051_top_1.iadr_o [8], cxrom_addr[8]);
  buf(\oc8051_top_1.iadr_o [9], cxrom_addr[9]);
  buf(\oc8051_top_1.iadr_o [10], cxrom_addr[10]);
  buf(\oc8051_top_1.iadr_o [11], cxrom_addr[11]);
  buf(\oc8051_top_1.iadr_o [12], cxrom_addr[12]);
  buf(\oc8051_top_1.iadr_o [13], cxrom_addr[13]);
  buf(\oc8051_top_1.iadr_o [14], cxrom_addr[14]);
  buf(\oc8051_top_1.iadr_o [15], cxrom_addr[15]);
  buf(\oc8051_top_1.sp [0], \oc8051_top_1.oc8051_memory_interface1.sp [0]);
  buf(\oc8051_top_1.sp [1], \oc8051_top_1.oc8051_memory_interface1.sp [1]);
  buf(\oc8051_top_1.sp [2], \oc8051_top_1.oc8051_memory_interface1.sp [2]);
  buf(\oc8051_top_1.sp [3], \oc8051_top_1.oc8051_memory_interface1.sp [3]);
  buf(\oc8051_top_1.sp [4], \oc8051_top_1.oc8051_memory_interface1.sp [4]);
  buf(\oc8051_top_1.sp [5], \oc8051_top_1.oc8051_memory_interface1.sp [5]);
  buf(\oc8051_top_1.sp [6], \oc8051_top_1.oc8051_memory_interface1.sp [6]);
  buf(\oc8051_top_1.sp [7], \oc8051_top_1.oc8051_memory_interface1.sp [7]);
  buf(\oc8051_top_1.sp_w [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [0]);
  buf(\oc8051_top_1.sp_w [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [1]);
  buf(\oc8051_top_1.sp_w [2], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [2]);
  buf(\oc8051_top_1.sp_w [3], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [3]);
  buf(\oc8051_top_1.sp_w [4], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [4]);
  buf(\oc8051_top_1.sp_w [5], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [5]);
  buf(\oc8051_top_1.sp_w [6], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [6]);
  buf(\oc8051_top_1.sp_w [7], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp_w [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.wr_sfr [0], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [0]);
  buf(\oc8051_top_1.wr_sfr [1], \oc8051_top_1.oc8051_decoder1.wr_sfr_o [1]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.ram_rd_sel [0], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [0]);
  buf(\oc8051_top_1.ram_rd_sel [1], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [1]);
  buf(\oc8051_top_1.ram_rd_sel [2], \oc8051_top_1.oc8051_decoder1.ram_rd_sel_o [2]);
  buf(\oc8051_top_1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [0]);
  buf(\oc8051_top_1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [1]);
  buf(\oc8051_top_1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel_o [2]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.ram_data [0], \oc8051_top_1.oc8051_memory_interface1.in_ram [0]);
  buf(\oc8051_top_1.ram_data [1], \oc8051_top_1.oc8051_memory_interface1.in_ram [1]);
  buf(\oc8051_top_1.ram_data [2], \oc8051_top_1.oc8051_memory_interface1.in_ram [2]);
  buf(\oc8051_top_1.ram_data [3], \oc8051_top_1.oc8051_memory_interface1.in_ram [3]);
  buf(\oc8051_top_1.ram_data [4], \oc8051_top_1.oc8051_memory_interface1.in_ram [4]);
  buf(\oc8051_top_1.ram_data [5], \oc8051_top_1.oc8051_memory_interface1.in_ram [5]);
  buf(\oc8051_top_1.ram_data [6], \oc8051_top_1.oc8051_memory_interface1.in_ram [6]);
  buf(\oc8051_top_1.ram_data [7], \oc8051_top_1.oc8051_memory_interface1.in_ram [7]);
  buf(\oc8051_top_1.ram_out [0], \oc8051_top_1.oc8051_memory_interface1.iram_out [0]);
  buf(\oc8051_top_1.ram_out [1], \oc8051_top_1.oc8051_memory_interface1.iram_out [1]);
  buf(\oc8051_top_1.ram_out [2], \oc8051_top_1.oc8051_memory_interface1.iram_out [2]);
  buf(\oc8051_top_1.ram_out [3], \oc8051_top_1.oc8051_memory_interface1.iram_out [3]);
  buf(\oc8051_top_1.ram_out [4], \oc8051_top_1.oc8051_memory_interface1.iram_out [4]);
  buf(\oc8051_top_1.ram_out [5], \oc8051_top_1.oc8051_memory_interface1.iram_out [5]);
  buf(\oc8051_top_1.ram_out [6], \oc8051_top_1.oc8051_memory_interface1.iram_out [6]);
  buf(\oc8051_top_1.ram_out [7], \oc8051_top_1.oc8051_memory_interface1.iram_out [7]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.wr_dat [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.wr_dat [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.wr_dat [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.wr_dat [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.wr_dat [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.wr_dat [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.wr_dat [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.wr_dat [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.wr_addr [0], \oc8051_top_1.oc8051_memory_interface1.wr_addr [0]);
  buf(\oc8051_top_1.wr_addr [1], \oc8051_top_1.oc8051_memory_interface1.wr_addr [1]);
  buf(\oc8051_top_1.wr_addr [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [2]);
  buf(\oc8051_top_1.wr_addr [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_addr [3]);
  buf(\oc8051_top_1.wr_addr [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_addr [4]);
  buf(\oc8051_top_1.wr_addr [5], \oc8051_top_1.oc8051_memory_interface1.wr_addr [5]);
  buf(\oc8051_top_1.wr_addr [6], \oc8051_top_1.oc8051_memory_interface1.wr_addr [6]);
  buf(\oc8051_top_1.rd_addr [0], \oc8051_top_1.oc8051_ram_top1.rd_addr [0]);
  buf(\oc8051_top_1.rd_addr [1], \oc8051_top_1.oc8051_ram_top1.rd_addr [1]);
  buf(\oc8051_top_1.rd_addr [2], \oc8051_top_1.oc8051_ram_top1.rd_addr [2]);
  buf(\oc8051_top_1.rd_addr [3], \oc8051_top_1.oc8051_ram_top1.rd_addr [3]);
  buf(\oc8051_top_1.rd_addr [4], \oc8051_top_1.oc8051_ram_top1.rd_addr [4]);
  buf(\oc8051_top_1.rd_addr [5], \oc8051_top_1.oc8051_ram_top1.rd_addr [5]);
  buf(\oc8051_top_1.rd_addr [6], \oc8051_top_1.oc8051_ram_top1.rd_addr [6]);
  buf(\oc8051_top_1.rd_addr [7], \oc8051_top_1.oc8051_ram_top1.rd_addr [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.bank_sel [0], \oc8051_top_1.oc8051_memory_interface1.rn [3]);
  buf(\oc8051_top_1.bank_sel [1], \oc8051_top_1.oc8051_memory_interface1.rn [4]);
  buf(\oc8051_top_1.idat_i [0], \oc8051_top_1.oc8051_memory_interface1.idat_i [0]);
  buf(\oc8051_top_1.idat_i [1], \oc8051_top_1.oc8051_memory_interface1.idat_i [1]);
  buf(\oc8051_top_1.idat_i [2], \oc8051_top_1.oc8051_memory_interface1.idat_i [2]);
  buf(\oc8051_top_1.idat_i [3], \oc8051_top_1.oc8051_memory_interface1.idat_i [3]);
  buf(\oc8051_top_1.idat_i [4], \oc8051_top_1.oc8051_memory_interface1.idat_i [4]);
  buf(\oc8051_top_1.idat_i [5], \oc8051_top_1.oc8051_memory_interface1.idat_i [5]);
  buf(\oc8051_top_1.idat_i [6], \oc8051_top_1.oc8051_memory_interface1.idat_i [6]);
  buf(\oc8051_top_1.idat_i [7], \oc8051_top_1.oc8051_memory_interface1.idat_i [7]);
  buf(\oc8051_top_1.idat_i [8], \oc8051_top_1.oc8051_memory_interface1.idat_i [8]);
  buf(\oc8051_top_1.idat_i [9], \oc8051_top_1.oc8051_memory_interface1.idat_i [9]);
  buf(\oc8051_top_1.idat_i [10], \oc8051_top_1.oc8051_memory_interface1.idat_i [10]);
  buf(\oc8051_top_1.idat_i [11], \oc8051_top_1.oc8051_memory_interface1.idat_i [11]);
  buf(\oc8051_top_1.idat_i [12], \oc8051_top_1.oc8051_memory_interface1.idat_i [12]);
  buf(\oc8051_top_1.idat_i [13], \oc8051_top_1.oc8051_memory_interface1.idat_i [13]);
  buf(\oc8051_top_1.idat_i [14], \oc8051_top_1.oc8051_memory_interface1.idat_i [14]);
  buf(\oc8051_top_1.idat_i [15], \oc8051_top_1.oc8051_memory_interface1.idat_i [15]);
  buf(\oc8051_top_1.idat_i [16], \oc8051_top_1.oc8051_memory_interface1.idat_i [16]);
  buf(\oc8051_top_1.idat_i [17], \oc8051_top_1.oc8051_memory_interface1.idat_i [17]);
  buf(\oc8051_top_1.idat_i [18], \oc8051_top_1.oc8051_memory_interface1.idat_i [18]);
  buf(\oc8051_top_1.idat_i [19], \oc8051_top_1.oc8051_memory_interface1.idat_i [19]);
  buf(\oc8051_top_1.idat_i [20], \oc8051_top_1.oc8051_memory_interface1.idat_i [20]);
  buf(\oc8051_top_1.idat_i [21], \oc8051_top_1.oc8051_memory_interface1.idat_i [21]);
  buf(\oc8051_top_1.idat_i [22], \oc8051_top_1.oc8051_memory_interface1.idat_i [22]);
  buf(\oc8051_top_1.idat_i [23], \oc8051_top_1.oc8051_memory_interface1.idat_i [23]);
  buf(\oc8051_top_1.idat_i [24], \oc8051_top_1.oc8051_memory_interface1.idat_i [24]);
  buf(\oc8051_top_1.idat_i [25], \oc8051_top_1.oc8051_memory_interface1.idat_i [25]);
  buf(\oc8051_top_1.idat_i [26], \oc8051_top_1.oc8051_memory_interface1.idat_i [26]);
  buf(\oc8051_top_1.idat_i [27], \oc8051_top_1.oc8051_memory_interface1.idat_i [27]);
  buf(\oc8051_top_1.idat_i [28], \oc8051_top_1.oc8051_memory_interface1.idat_i [28]);
  buf(\oc8051_top_1.idat_i [29], \oc8051_top_1.oc8051_memory_interface1.idat_i [29]);
  buf(\oc8051_top_1.idat_i [30], \oc8051_top_1.oc8051_memory_interface1.idat_i [30]);
  buf(\oc8051_top_1.idat_i [31], \oc8051_top_1.oc8051_memory_interface1.idat_i [31]);
  buf(\oc8051_top_1.rmw , \oc8051_top_1.oc8051_decoder1.rmw );
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.intr , \oc8051_top_1.oc8051_sfr1.oc8051_int1.intr );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_wait , \oc8051_top_1.oc8051_decoder1.mem_wait );
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.alu_op [0], \oc8051_top_1.oc8051_decoder1.alu_op_o [0]);
  buf(\oc8051_top_1.alu_op [1], \oc8051_top_1.oc8051_decoder1.alu_op_o [1]);
  buf(\oc8051_top_1.alu_op [2], \oc8051_top_1.oc8051_decoder1.alu_op_o [2]);
  buf(\oc8051_top_1.alu_op [3], \oc8051_top_1.oc8051_decoder1.alu_op_o [3]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.src1 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [0]);
  buf(\oc8051_top_1.src1 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [1]);
  buf(\oc8051_top_1.src1 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [2]);
  buf(\oc8051_top_1.src1 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [3]);
  buf(\oc8051_top_1.src1 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [4]);
  buf(\oc8051_top_1.src1 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [5]);
  buf(\oc8051_top_1.src1 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [6]);
  buf(\oc8051_top_1.src1 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src1 [7]);
  buf(\oc8051_top_1.src2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [0]);
  buf(\oc8051_top_1.src2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [1]);
  buf(\oc8051_top_1.src2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [2]);
  buf(\oc8051_top_1.src2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [3]);
  buf(\oc8051_top_1.src2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [4]);
  buf(\oc8051_top_1.src2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [5]);
  buf(\oc8051_top_1.src2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [6]);
  buf(\oc8051_top_1.src2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.src2 [7]);
  buf(\oc8051_top_1.src3 [0], \oc8051_top_1.oc8051_alu_src_sel1.src3 [0]);
  buf(\oc8051_top_1.src3 [1], \oc8051_top_1.oc8051_alu_src_sel1.src3 [1]);
  buf(\oc8051_top_1.src3 [2], \oc8051_top_1.oc8051_alu_src_sel1.src3 [2]);
  buf(\oc8051_top_1.src3 [3], \oc8051_top_1.oc8051_alu_src_sel1.src3 [3]);
  buf(\oc8051_top_1.src3 [4], \oc8051_top_1.oc8051_alu_src_sel1.src3 [4]);
  buf(\oc8051_top_1.src3 [5], \oc8051_top_1.oc8051_alu_src_sel1.src3 [5]);
  buf(\oc8051_top_1.src3 [6], \oc8051_top_1.oc8051_alu_src_sel1.src3 [6]);
  buf(\oc8051_top_1.src3 [7], \oc8051_top_1.oc8051_alu_src_sel1.src3 [7]);
  buf(\oc8051_top_1.des_acc [0], \oc8051_top_1.oc8051_memory_interface1.des_acc [0]);
  buf(\oc8051_top_1.des_acc [1], \oc8051_top_1.oc8051_memory_interface1.des_acc [1]);
  buf(\oc8051_top_1.des_acc [2], \oc8051_top_1.oc8051_memory_interface1.des_acc [2]);
  buf(\oc8051_top_1.des_acc [3], \oc8051_top_1.oc8051_memory_interface1.des_acc [3]);
  buf(\oc8051_top_1.des_acc [4], \oc8051_top_1.oc8051_memory_interface1.des_acc [4]);
  buf(\oc8051_top_1.des_acc [5], \oc8051_top_1.oc8051_memory_interface1.des_acc [5]);
  buf(\oc8051_top_1.des_acc [6], \oc8051_top_1.oc8051_memory_interface1.des_acc [6]);
  buf(\oc8051_top_1.des_acc [7], \oc8051_top_1.oc8051_memory_interface1.des_acc [7]);
  buf(\oc8051_top_1.des1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0]);
  buf(\oc8051_top_1.des1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1]);
  buf(\oc8051_top_1.des1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2]);
  buf(\oc8051_top_1.des1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3]);
  buf(\oc8051_top_1.des1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4]);
  buf(\oc8051_top_1.des1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5]);
  buf(\oc8051_top_1.des1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6]);
  buf(\oc8051_top_1.des1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7]);
  buf(\oc8051_top_1.des2 [0], \oc8051_top_1.oc8051_memory_interface1.des2 [0]);
  buf(\oc8051_top_1.des2 [1], \oc8051_top_1.oc8051_memory_interface1.des2 [1]);
  buf(\oc8051_top_1.des2 [2], \oc8051_top_1.oc8051_memory_interface1.des2 [2]);
  buf(\oc8051_top_1.des2 [3], \oc8051_top_1.oc8051_memory_interface1.des2 [3]);
  buf(\oc8051_top_1.des2 [4], \oc8051_top_1.oc8051_memory_interface1.des2 [4]);
  buf(\oc8051_top_1.des2 [5], \oc8051_top_1.oc8051_memory_interface1.des2 [5]);
  buf(\oc8051_top_1.des2 [6], \oc8051_top_1.oc8051_memory_interface1.des2 [6]);
  buf(\oc8051_top_1.des2 [7], \oc8051_top_1.oc8051_memory_interface1.des2 [7]);
  buf(\oc8051_top_1.desCy , \oc8051_top_1.oc8051_ram_top1.bit_data_in );
  buf(\oc8051_top_1.desAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in );
  buf(\oc8051_top_1.desOv , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in );
  buf(\oc8051_top_1.alu_cy , \oc8051_top_1.oc8051_cy_select1.data_out );
  buf(\oc8051_top_1.wr , \oc8051_top_1.wr_o );
  buf(\oc8051_top_1.rd , \oc8051_top_1.oc8051_decoder1.rd );
  buf(\oc8051_top_1.pc_wr_sel [0], \oc8051_top_1.oc8051_decoder1.pc_sel [0]);
  buf(\oc8051_top_1.pc_wr_sel [1], \oc8051_top_1.oc8051_decoder1.pc_sel [1]);
  buf(\oc8051_top_1.pc_wr_sel [2], \oc8051_top_1.oc8051_decoder1.pc_sel [2]);
  buf(\oc8051_top_1.op1_n [0], \oc8051_top_1.oc8051_decoder1.op_in [0]);
  buf(\oc8051_top_1.op1_n [1], \oc8051_top_1.oc8051_decoder1.op_in [1]);
  buf(\oc8051_top_1.op1_n [2], \oc8051_top_1.oc8051_decoder1.op_in [2]);
  buf(\oc8051_top_1.op1_n [3], \oc8051_top_1.oc8051_decoder1.op_in [3]);
  buf(\oc8051_top_1.op1_n [4], \oc8051_top_1.oc8051_decoder1.op_in [4]);
  buf(\oc8051_top_1.op1_n [5], \oc8051_top_1.oc8051_decoder1.op_in [5]);
  buf(\oc8051_top_1.op1_n [6], \oc8051_top_1.oc8051_decoder1.op_in [6]);
  buf(\oc8051_top_1.op1_n [7], \oc8051_top_1.oc8051_decoder1.op_in [7]);
  buf(\oc8051_top_1.op2_n [0], \oc8051_top_1.oc8051_memory_interface1.op2_out [0]);
  buf(\oc8051_top_1.op2_n [1], \oc8051_top_1.oc8051_memory_interface1.op2_out [1]);
  buf(\oc8051_top_1.op2_n [2], \oc8051_top_1.oc8051_memory_interface1.op2_out [2]);
  buf(\oc8051_top_1.op2_n [3], \oc8051_top_1.oc8051_memory_interface1.op2_out [3]);
  buf(\oc8051_top_1.op2_n [4], \oc8051_top_1.oc8051_memory_interface1.op2_out [4]);
  buf(\oc8051_top_1.op2_n [5], \oc8051_top_1.oc8051_memory_interface1.op2_out [5]);
  buf(\oc8051_top_1.op2_n [6], \oc8051_top_1.oc8051_memory_interface1.op2_out [6]);
  buf(\oc8051_top_1.op2_n [7], \oc8051_top_1.oc8051_memory_interface1.op2_out [7]);
  buf(\oc8051_top_1.op3_n [0], \oc8051_top_1.oc8051_memory_interface1.op3_out [0]);
  buf(\oc8051_top_1.op3_n [1], \oc8051_top_1.oc8051_memory_interface1.op3_out [1]);
  buf(\oc8051_top_1.op3_n [2], \oc8051_top_1.oc8051_memory_interface1.op3_out [2]);
  buf(\oc8051_top_1.op3_n [3], \oc8051_top_1.oc8051_memory_interface1.op3_out [3]);
  buf(\oc8051_top_1.op3_n [4], \oc8051_top_1.oc8051_memory_interface1.op3_out [4]);
  buf(\oc8051_top_1.op3_n [5], \oc8051_top_1.oc8051_memory_interface1.op3_out [5]);
  buf(\oc8051_top_1.op3_n [6], \oc8051_top_1.oc8051_memory_interface1.op3_out [6]);
  buf(\oc8051_top_1.op3_n [7], \oc8051_top_1.oc8051_memory_interface1.op3_out [7]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.comp_sel [0], \oc8051_top_1.oc8051_decoder1.comp_sel [0]);
  buf(\oc8051_top_1.comp_sel [1], \oc8051_top_1.oc8051_decoder1.comp_sel [1]);
  buf(\oc8051_top_1.eq , \oc8051_top_1.oc8051_decoder1.eq );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wr_ind , \oc8051_top_1.oc8051_memory_interface1.wr_ind );
  buf(\oc8051_top_1.op1_cur [0], \oc8051_top_1.oc8051_decoder1.op_cur [0]);
  buf(\oc8051_top_1.op1_cur [1], \oc8051_top_1.oc8051_decoder1.op_cur [1]);
  buf(\oc8051_top_1.op1_cur [2], \oc8051_top_1.oc8051_decoder1.op_cur [2]);
  buf(\oc8051_top_1.bit_addr , \oc8051_top_1.oc8051_decoder1.bit_addr );
  buf(\oc8051_top_1.bit_data , \oc8051_top_1.oc8051_memory_interface1.bit_in );
  buf(\oc8051_top_1.bit_out , \oc8051_top_1.oc8051_cy_select1.data_in );
  buf(\oc8051_top_1.bit_addr_o , \oc8051_top_1.oc8051_decoder1.bit_addr );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.iack_i , \oc8051_top_1.oc8051_memory_interface1.iack_i );
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(cxrom_addr[0], \oc8051_top_1.oc8051_memory_interface1.iadr_o [0]);
  buf(cxrom_addr[1], \oc8051_top_1.oc8051_memory_interface1.iadr_o [1]);
  buf(cxrom_addr[2], \oc8051_top_1.oc8051_memory_interface1.iadr_o [2]);
  buf(cxrom_addr[3], \oc8051_top_1.oc8051_memory_interface1.iadr_o [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(_10957_, 1'b0);
  buf(_10625_, 1'b1);
  buf(_33297_, _10625_);
  buf(_23698_, rst);
  buf(_33296_, _29226_);
  buf(_33295_, _02158_);
  buf(_33294_, _06159_);
  buf(_33293_, _10626_);
  buf(_33292_, _14540_);
  buf(_33291_, _17402_);
  buf(_33290_, _20930_);
  buf(_33289_, _23346_);
  buf(_33288_, _23699_);
  buf(_33287_, _24110_);
  buf(_33286_, _24521_);
  buf(_33285_, _24932_);
  buf(_33284_, _25343_);
  buf(_33283_, _25917_);
  buf(_33282_, _26728_);
  buf(_33281_, _27539_);
  buf(_33280_, _28350_);
  buf(_33279_, _28815_);
  buf(_33278_, _29227_);
  buf(_33277_, _29639_);
  buf(_33276_, _30050_);
  buf(_33275_, _30492_);
  buf(_33274_, _30969_);
  buf(_33273_, _00001_);
  buf(_33272_, _00440_);
  buf(_33271_, _00871_);
  buf(_33270_, _01281_);
  buf(_33269_, _01726_);
  buf(_33268_, _02159_);
  buf(_33267_, _02541_);
  buf(_33266_, _02878_);
  buf(_33265_, _03289_);
  buf(_33264_, _03630_);
  buf(_33263_, _04029_);
  buf(_33262_, _04419_);
  buf(_33261_, _04830_);
  buf(_33260_, _05287_);
  buf(_33259_, _05725_);
  buf(_33258_, _06160_);
  buf(_33257_, _06634_);
  buf(_33256_, _07049_);
  buf(_33255_, _07422_);
  buf(_33254_, _07840_);
  buf(_33253_, _08287_);
  buf(_33252_, _08791_);
  buf(_33251_, _09311_);
  buf(_33250_, _09801_);
  buf(_33249_, _10212_);
  buf(_33248_, _10627_);
  buf(_33247_, _11040_);
  buf(_33246_, _11450_);
  buf(_33245_, _11861_);
  buf(_33244_, _12271_);
  buf(_33243_, _12683_);
  buf(_33242_, _13094_);
  buf(_33241_, _13505_);
  buf(_33240_, _13872_);
  buf(_33239_, _14206_);
  buf(_33238_, _14541_);
  buf(_33237_, _14862_);
  buf(_33236_, _15140_);
  buf(_33235_, _15412_);
  buf(_33234_, _15688_);
  buf(_33233_, _15972_);
  buf(_33232_, _16254_);
  buf(_33231_, _16542_);
  buf(_33230_, _16828_);
  buf(_33229_, _17114_);
  buf(_33228_, _17403_);
  buf(_33227_, _17689_);
  buf(_33226_, _17976_);
  buf(_33225_, _18264_);
  buf(_33224_, _18551_);
  buf(_33223_, _18911_);
  buf(_33222_, _19310_);
  buf(_33221_, _19712_);
  buf(_33220_, _20122_);
  buf(_33219_, _20533_);
  buf(_33218_, _20931_);
  buf(_33217_, _21320_);
  buf(_33216_, _21708_);
  buf(_33215_, _22100_);
  buf(_33214_, _22521_);
  buf(_33213_, _22942_);
  buf(_33212_, _23263_);
  buf(_33211_, _23284_);
  buf(_33210_, _23304_);
  buf(_33209_, _23325_);
  buf(_33208_, _23347_);
  buf(_33207_, _23376_);
  buf(_33206_, _23417_);
  buf(_33205_, _23458_);
  buf(_33204_, _23499_);
  buf(_33203_, _23540_);
  buf(_33202_, _23581_);
  buf(_33201_, _23622_);
  buf(_33200_, _23663_);
  buf(_33199_, _23685_);
  buf(_33198_, _23700_);
  buf(_33197_, _23741_);
  buf(_33196_, _23782_);
  buf(_33195_, _23823_);
  buf(_33194_, _23864_);
  buf(_33193_, _23905_);
  buf(_33192_, _23946_);
  buf(_33191_, _23987_);
  buf(_33190_, _24028_);
  buf(_33189_, _24069_);
  buf(_33188_, _24111_);
  buf(_33187_, _24152_);
  buf(_33186_, _24193_);
  buf(_33185_, _24234_);
  buf(_33184_, _24275_);
  buf(_33183_, _24316_);
  buf(_33182_, _24357_);
  buf(_33181_, _24398_);
  buf(_33180_, _24439_);
  buf(_33179_, _24480_);
  buf(_33178_, _24522_);
  buf(_33177_, _24563_);
  buf(_33176_, _24604_);
  buf(_33175_, _24645_);
  buf(_33174_, _24686_);
  buf(_33173_, _24727_);
  buf(_33172_, _24768_);
  buf(_33171_, _24809_);
  buf(_33170_, _24850_);
  buf(_33169_, _24891_);
  buf(_33168_, _24933_);
  buf(_33167_, _24974_);
  buf(_33166_, _25015_);
  buf(_33165_, _25056_);
  buf(_33164_, _25097_);
  buf(_33163_, _25138_);
  buf(_33162_, _25179_);
  buf(_33161_, _25220_);
  buf(_33160_, _25261_);
  buf(_33159_, _25302_);
  buf(_33158_, _25344_);
  buf(_33157_, _25385_);
  buf(_33156_, _25426_);
  buf(_33155_, _25467_);
  buf(_33154_, _25508_);
  buf(_33153_, _25549_);
  buf(_33152_, _25593_);
  buf(_33151_, _25674_);
  buf(_33150_, _25755_);
  buf(_33149_, _25836_);
  buf(_33148_, _25918_);
  buf(_33147_, _25999_);
  buf(_33146_, _26080_);
  buf(_33145_, _26161_);
  buf(_33144_, _26242_);
  buf(_33143_, _26323_);
  buf(_33142_, _26404_);
  buf(_33141_, _26485_);
  buf(_33140_, _26566_);
  buf(_33139_, _26647_);
  buf(_33138_, _26729_);
  buf(_33137_, _26810_);
  buf(_33136_, _26891_);
  buf(_33135_, _26972_);
  buf(_33134_, _27053_);
  buf(_33133_, _27134_);
  buf(_33132_, _27215_);
  buf(_33131_, _27296_);
  buf(_33130_, _27377_);
  buf(_33129_, _27458_);
  buf(_33128_, _27540_);
  buf(_33127_, _27621_);
  buf(_33126_, _27702_);
  buf(_33125_, _27783_);
  buf(_33124_, _27864_);
  buf(_33123_, _27945_);
  buf(_33122_, _28026_);
  buf(_33121_, _28107_);
  buf(_33120_, _28188_);
  buf(_33119_, _28269_);
  buf(_33118_, _28351_);
  buf(_33117_, _28432_);
  buf(_33116_, _28487_);
  buf(_33115_, _28528_);
  buf(_33114_, _28569_);
  buf(_33113_, _28610_);
  buf(_33112_, _28651_);
  buf(_33111_, _28692_);
  buf(_33110_, _28733_);
  buf(_33109_, _28774_);
  buf(_33108_, _28816_);
  buf(_33107_, _28857_);
  buf(_33106_, _28898_);
  buf(_33105_, _28939_);
  buf(_33104_, _28980_);
  buf(_33103_, _29021_);
  buf(_33102_, _29062_);
  buf(_33101_, _29103_);
  buf(_33100_, _29144_);
  buf(_33099_, _29185_);
  buf(_33098_, _29228_);
  buf(_33097_, _29269_);
  buf(_33096_, _29311_);
  buf(_33095_, _29352_);
  buf(_33094_, _29393_);
  buf(_33093_, _29434_);
  buf(_33092_, _29475_);
  buf(_33091_, _29516_);
  buf(_33090_, _29557_);
  buf(_33089_, _29598_);
  buf(_33088_, _29640_);
  buf(_33087_, _29681_);
  buf(_33086_, _29722_);
  buf(_33085_, _29763_);
  buf(_33084_, _29804_);
  buf(_33083_, _29845_);
  buf(_33082_, _29886_);
  buf(_33081_, _29927_);
  buf(_33080_, _29968_);
  buf(_33079_, _30009_);
  buf(_33078_, _30051_);
  buf(_33077_, _30092_);
  buf(_33076_, _30132_);
  buf(_33075_, _30173_);
  buf(_33074_, _30214_);
  buf(_33073_, _30254_);
  buf(_33072_, _30303_);
  buf(_30316_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  buf(_33071_, _30352_);
  buf(_33070_, _30398_);
  buf(_33069_, _30443_);
  buf(_33068_, _30493_);
  buf(_33067_, _30539_);
  buf(_33066_, _30600_);
  buf(_33065_, _30646_);
  buf(_30658_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  buf(_33064_, _30695_);
  buf(_33063_, _30738_);
  buf(_33062_, _30787_);
  buf(_33061_, _30835_);
  buf(_33060_, _30883_);
  buf(_30894_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r );
  buf(_33059_, _30925_);
  buf(_33058_, _30970_);
  buf(_33057_, _31021_);
  buf(_33056_, _31068_);
  buf(_33055_, _31111_);
  buf(_33054_, _31155_);
  buf(_33053_, _31199_);
  buf(_33052_, _31248_);
  buf(_33051_, _31297_);
  buf(_33050_, _31338_);
  buf(_33049_, _31379_);
  buf(_33048_, _00002_);
  buf(_33047_, _00045_);
  buf(_33046_, _00086_);
  buf(_33045_, _00127_);
  buf(_33044_, _00171_);
  buf(_33043_, _00215_);
  buf(_33042_, _00262_);
  buf(_33041_, _00304_);
  buf(_33040_, _00353_);
  buf(_33039_, _00395_);
  buf(_33038_, _00441_);
  buf(_33037_, _00485_);
  buf(_33036_, _00530_);
  buf(_33035_, _00579_);
  buf(_33034_, _00620_);
  buf(_33033_, _00663_);
  buf(_33032_, _00704_);
  buf(_33031_, _00745_);
  buf(_33030_, _00787_);
  buf(_33029_, _00830_);
  buf(_33028_, _00872_);
  buf(_33027_, _00910_);
  buf(_33026_, _00945_);
  buf(_33025_, _00987_);
  buf(_33024_, _01038_);
  buf(_33023_, _01071_);
  buf(_33022_, _01105_);
  buf(_33021_, _01142_);
  buf(_33020_, _01181_);
  buf(_33019_, _01232_);
  buf(_33018_, _01282_);
  buf(_33017_, _01328_);
  buf(_33016_, _01371_);
  buf(_33015_, _01419_);
  buf(_33014_, _01471_);
  buf(_33013_, _01518_);
  buf(_33012_, _01559_);
  buf(_33011_, _01602_);
  buf(_33010_, _01643_);
  buf(_33009_, _01680_);
  buf(_33008_, _01727_);
  buf(_33007_, _01770_);
  buf(_33006_, _01811_);
  buf(_33005_, _01852_);
  buf(_33004_, _01895_);
  buf(_33003_, _01937_);
  buf(_33002_, _01979_);
  buf(_33001_, _02032_);
  buf(_33000_, _02073_);
  buf(_32999_, _02117_);
  buf(_32998_, _02160_);
  buf(_32997_, _02200_);
  buf(_32996_, _02246_);
  buf(_32995_, _02286_);
  buf(_32994_, _02326_);
  buf(_32993_, _02366_);
  buf(_32992_, _02404_);
  buf(_32991_, _02443_);
  buf(_32990_, _02481_);
  buf(_32989_, _02509_);
  buf(_32988_, _02542_);
  buf(_32987_, _02575_);
  buf(_32986_, _02611_);
  buf(_02619_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(_32985_, _02644_);
  buf(_02652_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(_32984_, _02677_);
  buf(_02686_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(_32983_, _02711_);
  buf(_32982_, _02743_);
  buf(_32981_, _02774_);
  buf(_32980_, _02814_);
  buf(_32979_, _02846_);
  buf(_02855_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(_32978_, _02879_);
  buf(_32977_, _02912_);
  buf(_32976_, _02947_);
  buf(_32975_, _02980_);
  buf(_32974_, _03020_);
  buf(_32973_, _03062_);
  buf(_32972_, _03107_);
  buf(_32971_, _03149_);
  buf(_32970_, _03199_);
  buf(_32969_, _03239_);
  buf(_32968_, _03290_);
  buf(_32967_, _03339_);
  buf(_32966_, _03385_);
  buf(_32965_, _03422_);
  buf(_32964_, _03457_);
  buf(_32963_, _03495_);
  buf(_32962_, _03535_);
  buf(_32961_, _03546_);
  buf(_32960_, _03562_);
  buf(_32959_, _03592_);
  buf(_32958_, _03631_);
  buf(_32957_, _03669_);
  buf(_32956_, _03708_);
  buf(_32955_, _03744_);
  buf(_32954_, _03782_);
  buf(_32953_, _03836_);
  buf(_32952_, _03873_);
  buf(_32951_, _03910_);
  buf(_32950_, _03951_);
  buf(_32949_, _03990_);
  buf(_32948_, _04030_);
  buf(_32947_, _04068_);
  buf(_32946_, _04107_);
  buf(_32945_, _04145_);
  buf(_32944_, _04184_);
  buf(_32943_, _04222_);
  buf(_32942_, _04255_);
  buf(_32941_, _04294_);
  buf(_32940_, _04331_);
  buf(_32939_, _04374_);
  buf(_32938_, _04420_);
  buf(_32937_, _04460_);
  buf(_32936_, _04499_);
  buf(_32935_, _04538_);
  buf(_32934_, _04575_);
  buf(_32933_, _04610_);
  buf(_32932_, _04651_);
  buf(_32931_, _04691_);
  buf(_32930_, _04735_);
  buf(_32929_, _04784_);
  buf(_32928_, _04831_);
  buf(_32927_, _04874_);
  buf(_32926_, _04922_);
  buf(_32925_, _04962_);
  buf(_32924_, _04998_);
  buf(_32923_, _05038_);
  buf(_32922_, _05103_);
  buf(_32921_, _05169_);
  buf(_32920_, _05210_);
  buf(_32919_, _05250_);
  buf(_32918_, _05288_);
  buf(_32917_, _05328_);
  buf(_32916_, _05378_);
  buf(_32915_, _05434_);
  buf(_32914_, _05488_);
  buf(_32913_, _05522_);
  buf(_32912_, _05559_);
  buf(_32911_, _05600_);
  buf(_32910_, _05647_);
  buf(_32909_, _05686_);
  buf(_32908_, _05726_);
  buf(_32907_, _05766_);
  buf(_32906_, _05804_);
  buf(_32905_, _05842_);
  buf(_32904_, _05881_);
  buf(_32903_, _05929_);
  buf(_32902_, _05980_);
  buf(_32901_, _06018_);
  buf(_06028_, t2ex_i);
  buf(_32900_, _06070_);
  buf(_32899_, _06112_);
  buf(_32898_, _06161_);
  buf(_32897_, _06206_);
  buf(_32896_, _06246_);
  buf(_32895_, _06283_);
  buf(_32894_, _06324_);
  buf(_32893_, _06366_);
  buf(_32892_, _06417_);
  buf(_32891_, _06463_);
  buf(_32890_, _06514_);
  buf(_32889_, _06575_);
  buf(_32888_, _06635_);
  buf(_32887_, _06676_);
  buf(_32886_, _06718_);
  buf(_32885_, _06759_);
  buf(_32884_, _06800_);
  buf(_32883_, _06841_);
  buf(_32882_, _06882_);
  buf(_32881_, _06923_);
  buf(_32880_, _06966_);
  buf(_32879_, _07008_);
  buf(_32878_, _07050_);
  buf(_32877_, _07091_);
  buf(_32876_, _07132_);
  buf(_32875_, _07161_);
  buf(_32874_, _07196_);
  buf(_32873_, _07230_);
  buf(_32872_, _07269_);
  buf(_32871_, _07307_);
  buf(_32870_, _07346_);
  buf(_32869_, _07383_);
  buf(_32868_, _07423_);
  buf(_32867_, _07461_);
  buf(_32866_, _07498_);
  buf(_32865_, _07537_);
  buf(_32864_, _07583_);
  buf(_32863_, _07623_);
  buf(_32862_, _07664_);
  buf(_32861_, _07707_);
  buf(_32860_, _07752_);
  buf(_32859_, _07795_);
  buf(_32858_, _07841_);
  buf(_32857_, _07887_);
  buf(_32856_, _07933_);
  buf(_32855_, _07974_);
  buf(_32854_, _08024_);
  buf(_32853_, _08072_);
  buf(_32852_, _08114_);
  buf(_32851_, _08156_);
  buf(_32850_, _08199_);
  buf(_32849_, _08243_);
  buf(_32848_, _08288_);
  buf(_32847_, _08332_);
  buf(_32846_, _08378_);
  buf(_32845_, _08444_);
  buf(_32844_, _08508_);
  buf(_32843_, _08572_);
  buf(_32842_, _08616_);
  buf(_32841_, _08657_);
  buf(_32840_, _08698_);
  buf(_32839_, _08750_);
  buf(_32838_, _08792_);
  buf(_32837_, _08845_);
  buf(_32836_, _08897_);
  buf(_32835_, _08959_);
  buf(_32834_, _09014_);
  buf(_32833_, _09071_);
  buf(_32832_, _09112_);
  buf(_32831_, _09158_);
  buf(_32830_, _09208_);
  buf(_32829_, _09259_);
  buf(_32828_, _09312_);
  buf(_32827_, _09361_);
  buf(_32826_, _09415_);
  buf(_32825_, _09463_);
  buf(_32824_, _09516_);
  buf(_32823_, _09566_);
  buf(_32822_, _09617_);
  buf(_32821_, _09672_);
  buf(_32820_, _09719_);
  buf(_32819_, _09760_);
  buf(_32818_, _09802_);
  buf(_32817_, _09843_);
  buf(_32816_, _09884_);
  buf(_32815_, _09925_);
  buf(_32814_, _09966_);
  buf(_32813_, _10007_);
  buf(_32812_, _10048_);
  buf(_32811_, _10089_);
  buf(_32810_, _10130_);
  buf(_32809_, _10171_);
  buf(_32808_, _10213_);
  buf(_32807_, _10255_);
  buf(_32806_, _10298_);
  buf(_32805_, _10339_);
  buf(_32804_, _10380_);
  buf(_32803_, _10421_);
  buf(_32802_, _10461_);
  buf(_32801_, _10502_);
  buf(_32800_, _10543_);
  buf(_32799_, _10584_);
  buf(_32798_, _10628_);
  buf(_32797_, _10669_);
  buf(_32796_, _10710_);
  buf(_32795_, _10751_);
  buf(_10762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(_32794_, _10793_);
  buf(_32793_, _10834_);
  buf(_32792_, _10875_);
  buf(_32791_, _10916_);
  buf(_32790_, _10957_);
  buf(_32789_, _10988_);
  buf(_32788_, _11029_);
  buf(_32787_, _11071_);
  buf(_32786_, _11112_);
  buf(_32785_, _11153_);
  buf(_32784_, _11194_);
  buf(_32783_, _11235_);
  buf(_32782_, _11275_);
  buf(_32781_, _11316_);
  buf(_32780_, _11357_);
  buf(_32779_, _11398_);
  buf(_32778_, _11439_);
  buf(_32777_, _11481_);
  buf(_32776_, _11522_);
  buf(_32775_, _11563_);
  buf(_32774_, _11604_);
  buf(_32773_, _11645_);
  buf(_32772_, _11686_);
  buf(_32771_, _11727_);
  buf(_32770_, _11768_);
  buf(_32769_, _11809_);
  buf(_32768_, _11850_);
  buf(_32767_, _11892_);
  buf(_32766_, _11933_);
  buf(_32765_, _11974_);
  buf(_32764_, _12015_);
  buf(_32763_, _12055_);
  buf(_32762_, _12096_);
  buf(_32761_, _12137_);
  buf(_32760_, _12178_);
  buf(_32759_, _12219_);
  buf(_32758_, _12260_);
  buf(_32757_, _12302_);
  buf(_32756_, _12343_);
  buf(_32755_, _12384_);
  buf(_32754_, _12425_);
  buf(_32753_, _12466_);
  buf(_32752_, _12507_);
  buf(_32751_, _12548_);
  buf(_32750_, _12589_);
  buf(_32749_, _12630_);
  buf(_12641_, t1_i);
  buf(_32748_, _12672_);
  buf(_12684_, t0_i);
  buf(_32747_, _12715_);
  buf(_32746_, _12756_);
  buf(_32745_, _12797_);
  buf(_32744_, _12837_);
  buf(_32743_, _12878_);
  buf(_32742_, _12919_);
  buf(_32741_, _12960_);
  buf(_32740_, _13001_);
  buf(_32739_, _13042_);
  buf(_32738_, _13083_);
  buf(_32737_, _13125_);
  buf(_32736_, _13166_);
  buf(_32735_, _13207_);
  buf(_32734_, _13248_);
  buf(_32733_, _13289_);
  buf(_32732_, _13330_);
  buf(_32731_, _13371_);
  buf(_32730_, _13412_);
  buf(_32729_, _13453_);
  buf(_32728_, _13494_);
  buf(_32727_, _13536_);
  buf(_32726_, _13577_);
  buf(_32725_, _13618_);
  buf(_32724_, _13655_);
  buf(_32723_, _13692_);
  buf(_32722_, _13728_);
  buf(_32721_, _13763_);
  buf(_32720_, _13796_);
  buf(_32719_, _13830_);
  buf(_32718_, _13863_);
  buf(_32717_, _13898_);
  buf(_32716_, _13931_);
  buf(_32715_, _13964_);
  buf(_32714_, _13998_);
  buf(_32713_, _14031_);
  buf(_32712_, _14064_);
  buf(_32711_, _14097_);
  buf(_32710_, _14131_);
  buf(_32709_, _14164_);
  buf(_32708_, _14197_);
  buf(_32707_, _14231_);
  buf(_32706_, _14265_);
  buf(_32705_, _14298_);
  buf(_32704_, _14331_);
  buf(_32703_, _14364_);
  buf(_32702_, _14398_);
  buf(_32701_, _14431_);
  buf(_32700_, _14464_);
  buf(_32699_, _14497_);
  buf(_32698_, _14531_);
  buf(_32697_, _14566_);
  buf(_32696_, _14599_);
  buf(_32695_, _14632_);
  buf(_32694_, _14666_);
  buf(_32693_, _14699_);
  buf(_32692_, _14732_);
  buf(_32691_, _14765_);
  buf(_32690_, _14798_);
  buf(_32689_, _14827_);
  buf(_32688_, _14854_);
  buf(_32687_, _14883_);
  buf(_32686_, _14911_);
  buf(_32685_, _14938_);
  buf(_32684_, _14966_);
  buf(_32683_, _14994_);
  buf(_32682_, _15021_);
  buf(_32681_, _15049_);
  buf(_32680_, _15077_);
  buf(_32679_, _15104_);
  buf(_32678_, _15132_);
  buf(_32677_, _15161_);
  buf(_32676_, _15188_);
  buf(_32675_, _15216_);
  buf(_32674_, _15244_);
  buf(_32673_, _15271_);
  buf(_15473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  buf(_37331_[7], _15488_);
  buf(_15535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  buf(_37358_[7], _15543_);
  buf(_15591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  buf(_37369_[7], _15598_);
  buf(_15633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  buf(_37380_[7], _15640_);
  buf(_15689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  buf(_37391_[7], _15697_);
  buf(_15724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  buf(_37402_[7], _15732_);
  buf(_15760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  buf(_37413_[7], _15767_);
  buf(_15795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  buf(_37417_[7], _15803_);
  buf(_15850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  buf(_37418_[7], _15858_);
  buf(_15886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  buf(_37330_[7], _15893_);
  buf(_15921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  buf(_37173_[7], _15929_);
  buf(_15956_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  buf(_37184_[7], _15964_);
  buf(_15999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  buf(_37195_[7], _16007_);
  buf(_16035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  buf(_37206_[7], _16042_);
  buf(_16070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  buf(_37216_[7], _16078_);
  buf(_16105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  buf(_37217_[7], _16113_);
  buf(_16161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  buf(_37218_[7], _16168_);
  buf(_16189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  buf(_37226_[7], _16197_);
  buf(_16218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  buf(_37356_[7], _16226_);
  buf(_16247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  buf(_37357_[7], _16255_);
  buf(_16276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  buf(_37359_[7], _16284_);
  buf(_16305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  buf(_37360_[7], _16313_);
  buf(_16334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  buf(_37361_[7], _16341_);
  buf(_16362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  buf(_37362_[7], _16370_);
  buf(_16391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  buf(_37363_[7], _16399_);
  buf(_16420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  buf(_37364_[7], _16427_);
  buf(_16448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  buf(_37365_[7], _16456_);
  buf(_16477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  buf(_37366_[7], _16485_);
  buf(_16506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  buf(_37367_[7], _16513_);
  buf(_16534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  buf(_37368_[7], _16543_);
  buf(_16564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  buf(_37370_[7], _16572_);
  buf(_16593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  buf(_37371_[7], _16600_);
  buf(_16648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  buf(_37372_[7], _16656_);
  buf(_16677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  buf(_37373_[7], _16684_);
  buf(_16705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  buf(_37374_[7], _16713_);
  buf(_16734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  buf(_37375_[7], _16742_);
  buf(_16763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  buf(_37376_[7], _16770_);
  buf(_16791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  buf(_37377_[7], _16799_);
  buf(_16820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  buf(_37378_[7], _16829_);
  buf(_16850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  buf(_37379_[7], _16857_);
  buf(_16878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  buf(_37381_[7], _16886_);
  buf(_16907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  buf(_37382_[7], _16915_);
  buf(_16936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  buf(_37383_[7], _16943_);
  buf(_16964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  buf(_37384_[7], _16972_);
  buf(_16993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  buf(_37385_[7], _17001_);
  buf(_17022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  buf(_37386_[7], _17029_);
  buf(_17050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  buf(_37387_[7], _17058_);
  buf(_17079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  buf(_37388_[7], _17087_);
  buf(_17122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  buf(_37389_[7], _17130_);
  buf(_17151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  buf(_37390_[7], _17158_);
  buf(_17179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  buf(_37392_[7], _17187_);
  buf(_17208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  buf(_37393_[7], _17216_);
  buf(_17237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  buf(_37394_[7], _17244_);
  buf(_17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  buf(_37395_[7], _17273_);
  buf(_17294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  buf(_37396_[7], _17302_);
  buf(_17323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  buf(_37397_[7], _17330_);
  buf(_17351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  buf(_37398_[7], _17359_);
  buf(_17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  buf(_37399_[7], _17388_);
  buf(_17411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  buf(_37400_[7], _17418_);
  buf(_17439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  buf(_37401_[7], _17447_);
  buf(_17468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  buf(_37403_[7], _17476_);
  buf(_17497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  buf(_37404_[7], _17504_);
  buf(_17525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  buf(_37405_[7], _17533_);
  buf(_17554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  buf(_37406_[7], _17562_);
  buf(_17609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  buf(_37407_[7], _17617_);
  buf(_17638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  buf(_37408_[7], _17646_);
  buf(_17667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  buf(_37409_[7], _17674_);
  buf(_17696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  buf(_37410_[7], _17704_);
  buf(_17725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  buf(_37411_[7], _17733_);
  buf(_17754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  buf(_37412_[7], _17761_);
  buf(_17782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  buf(_37303_[7], _17790_);
  buf(_17811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  buf(_37304_[7], _17819_);
  buf(_17840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  buf(_37414_[7], _17847_);
  buf(_17868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  buf(_37415_[7], _17876_);
  buf(_17897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  buf(_37416_[7], _17905_);
  buf(_17926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  buf(_37305_[7], _17933_);
  buf(_17954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  buf(_37306_[7], _17962_);
  buf(_17984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  buf(_37307_[7], _17992_);
  buf(_18013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  buf(_37308_[7], _18020_);
  buf(_18041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  buf(_37309_[7], _18049_);
  buf(_18077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  buf(_37310_[7], _18084_);
  buf(_18105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  buf(_37311_[7], _18113_);
  buf(_18134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  buf(_37312_[7], _18142_);
  buf(_18163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  buf(_37313_[7], _18170_);
  buf(_18191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  buf(_37314_[7], _18199_);
  buf(_18220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  buf(_37315_[7], _18228_);
  buf(_18249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  buf(_37316_[7], _18256_);
  buf(_18278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  buf(_37317_[7], _18286_);
  buf(_18307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  buf(_37318_[7], _18315_);
  buf(_18336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  buf(_37319_[7], _18343_);
  buf(_18364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  buf(_37320_[7], _18372_);
  buf(_18393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  buf(_37321_[7], _18401_);
  buf(_18422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  buf(_37322_[7], _18429_);
  buf(_18450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  buf(_37323_[7], _18458_);
  buf(_18479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  buf(_37324_[7], _18487_);
  buf(_18508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  buf(_37325_[7], _18515_);
  buf(_18543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  buf(_37326_[7], _18552_);
  buf(_18573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  buf(_37327_[7], _18580_);
  buf(_18599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  buf(_37328_[7], _18608_);
  buf(_18633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  buf(_37329_[7], _18642_);
  buf(_18667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  buf(_37163_[7], _18676_);
  buf(_18701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  buf(_37164_[7], _18710_);
  buf(_18735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  buf(_37165_[7], _18744_);
  buf(_18775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  buf(_37166_[7], _18786_);
  buf(_18817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  buf(_37167_[7], _18828_);
  buf(_18859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  buf(_37168_[7], _18870_);
  buf(_18900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  buf(_37169_[7], _18912_);
  buf(_18943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  buf(_37170_[7], _18954_);
  buf(_18985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  buf(_37171_[7], _18996_);
  buf(_19026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  buf(_37172_[7], _19037_);
  buf(_19068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  buf(_37174_[7], _19079_);
  buf(_19109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  buf(_37175_[7], _19120_);
  buf(_19161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  buf(_37176_[7], _19171_);
  buf(_19202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  buf(_37177_[7], _19213_);
  buf(_19236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  buf(_37178_[7], _19246_);
  buf(_19272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  buf(_37179_[7], _19281_);
  buf(_19311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  buf(_37180_[7], _19322_);
  buf(_19352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  buf(_37181_[7], _19363_);
  buf(_19392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  buf(_37182_[7], _19403_);
  buf(_19432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  buf(_37183_[7], _19443_);
  buf(_19472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  buf(_37185_[7], _19483_);
  buf(_19512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  buf(_37186_[7], _19523_);
  buf(_19552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  buf(_37187_[7], _19563_);
  buf(_19592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  buf(_37188_[7], _19603_);
  buf(_19632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  buf(_37189_[7], _19643_);
  buf(_19672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  buf(_37190_[7], _19683_);
  buf(_19713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  buf(_37191_[7], _19724_);
  buf(_19754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  buf(_37192_[7], _19764_);
  buf(_19844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  buf(_37193_[7], _19854_);
  buf(_19885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  buf(_37194_[7], _19896_);
  buf(_19926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  buf(_37196_[7], _19937_);
  buf(_19967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  buf(_37197_[7], _19978_);
  buf(_20008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  buf(_37198_[7], _20019_);
  buf(_20050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  buf(_37199_[7], _20060_);
  buf(_20091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  buf(_37200_[7], _20102_);
  buf(_20133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  buf(_37201_[7], _20144_);
  buf(_20174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  buf(_37202_[7], _20185_);
  buf(_20215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  buf(_37203_[7], _20226_);
  buf(_20256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  buf(_37204_[7], _20267_);
  buf(_20298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  buf(_37205_[7], _20308_);
  buf(_20339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  buf(_37207_[7], _20350_);
  buf(_20380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  buf(_37208_[7], _20391_);
  buf(_20421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  buf(_37209_[7], _20432_);
  buf(_20462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  buf(_37210_[7], _20473_);
  buf(_20512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  buf(_37211_[7], _20522_);
  buf(_20553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  buf(_37212_[7], _20563_);
  buf(_20593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  buf(_37213_[7], _20604_);
  buf(_20633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  buf(_37214_[7], _20644_);
  buf(_20674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  buf(_37215_[7], _20684_);
  buf(_20714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  buf(_37332_[7], _20724_);
  buf(_20754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  buf(_37333_[7], _20765_);
  buf(_20793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  buf(_37334_[7], _20804_);
  buf(_20832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  buf(_37335_[7], _20842_);
  buf(_20871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  buf(_37336_[7], _20881_);
  buf(_20909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  buf(_37337_[7], _20920_);
  buf(_20950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  buf(_37338_[7], _20960_);
  buf(_20989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  buf(_37339_[7], _20999_);
  buf(_21028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  buf(_37340_[7], _21038_);
  buf(_21067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  buf(_37341_[7], _21077_);
  buf(_21106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  buf(_37342_[7], _21116_);
  buf(_21154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  buf(_37343_[7], _21164_);
  buf(_21193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  buf(_37344_[7], _21203_);
  buf(_21232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  buf(_37345_[7], _21242_);
  buf(_21271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  buf(_37346_[7], _21281_);
  buf(_21310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  buf(_37347_[7], _21321_);
  buf(_21350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  buf(_37348_[7], _21360_);
  buf(_21388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  buf(_37349_[7], _21399_);
  buf(_21427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  buf(_37350_[7], _21437_);
  buf(_21466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  buf(_37351_[7], _21476_);
  buf(_21504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  buf(_37352_[7], _21515_);
  buf(_21543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  buf(_37353_[7], _21553_);
  buf(_21582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  buf(_37354_[7], _21592_);
  buf(_21620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  buf(_37355_[7], _21631_);
  buf(_21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  buf(_37219_[7], _21669_);
  buf(_21698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  buf(_37220_[7], _21709_);
  buf(_21737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  buf(_37221_[7], _21748_);
  buf(_21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  buf(_37222_[7], _21796_);
  buf(_21825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  buf(_37223_[7], _21835_);
  buf(_21863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  buf(_37224_[7], _21874_);
  buf(_21902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  buf(_37225_[7], _21912_);
  buf(_21941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  buf(_37227_[7], _21951_);
  buf(_21980_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  buf(_37228_[7], _21990_);
  buf(_22018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  buf(_37229_[7], _22029_);
  buf(_22058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  buf(_37230_[7], _22069_);
  buf(_22101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  buf(_37231_[7], _22112_);
  buf(_22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  buf(_37232_[7], _22154_);
  buf(_22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  buf(_37233_[7], _22196_);
  buf(_22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  buf(_37234_[7], _22238_);
  buf(_22269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  buf(_37235_[7], _22280_);
  buf(_22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  buf(_37236_[7], _22322_);
  buf(_22353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  buf(_37237_[7], _22364_);
  buf(_22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  buf(_37238_[7], _22406_);
  buf(_22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  buf(_37239_[7], _22468_);
  buf(_22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  buf(_37240_[7], _22510_);
  buf(_22542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  buf(_37241_[7], _22553_);
  buf(_22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  buf(_37242_[7], _22595_);
  buf(_22626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  buf(_37243_[7], _22637_);
  buf(_22668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  buf(_37244_[7], _22679_);
  buf(_22710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  buf(_37245_[7], _22721_);
  buf(_22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  buf(_37246_[7], _22763_);
  buf(_22794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  buf(_37247_[7], _22805_);
  buf(_22836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  buf(_37248_[7], _22847_);
  buf(_22878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  buf(_37249_[7], _22889_);
  buf(_22920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  buf(_37250_[7], _22931_);
  buf(_22963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  buf(_37251_[7], _22974_);
  buf(_23005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  buf(_37252_[7], _23016_);
  buf(_23047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  buf(_37253_[7], _23058_);
  buf(_23089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  buf(_37254_[7], _23100_);
  buf(_23141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  buf(_37255_[7], _23152_);
  buf(_23183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  buf(_37256_[7], _23194_);
  buf(_23225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  buf(_37257_[7], _23236_);
  buf(_23258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  buf(_37258_[7], _23259_);
  buf(_23260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  buf(_37259_[7], _23261_);
  buf(_23262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  buf(_37260_[7], _23264_);
  buf(_23265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  buf(_37261_[7], _23266_);
  buf(_23267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  buf(_37262_[7], _23268_);
  buf(_23269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  buf(_37263_[7], _23270_);
  buf(_23271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  buf(_37264_[7], _23272_);
  buf(_23273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  buf(_37265_[7], _23274_);
  buf(_23275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  buf(_37266_[7], _23276_);
  buf(_23277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  buf(_37267_[7], _23278_);
  buf(_23279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  buf(_37268_[7], _23280_);
  buf(_23281_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  buf(_37269_[7], _23282_);
  buf(_23283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  buf(_37270_[7], _23285_);
  buf(_23286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  buf(_37271_[7], _23287_);
  buf(_23288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  buf(_37272_[7], _23289_);
  buf(_23290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  buf(_37273_[7], _23291_);
  buf(_23292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  buf(_37274_[7], _23293_);
  buf(_23294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  buf(_37275_[7], _23295_);
  buf(_23296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  buf(_37276_[7], _23297_);
  buf(_23298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  buf(_37277_[7], _23299_);
  buf(_23300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  buf(_37278_[7], _23301_);
  buf(_23302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  buf(_37279_[7], _23303_);
  buf(_23305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  buf(_37280_[7], _23306_);
  buf(_23307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  buf(_37281_[7], _23308_);
  buf(_23309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  buf(_37282_[7], _23310_);
  buf(_23311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  buf(_37283_[7], _23312_);
  buf(_23313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  buf(_37284_[7], _23314_);
  buf(_23315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  buf(_37285_[7], _23316_);
  buf(_23317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  buf(_37286_[7], _23318_);
  buf(_23319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  buf(_37287_[7], _23320_);
  buf(_23321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  buf(_37288_[7], _23322_);
  buf(_23323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  buf(_37289_[7], _23324_);
  buf(_23326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  buf(_37290_[7], _23327_);
  buf(_23328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  buf(_37291_[7], _23329_);
  buf(_23330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  buf(_37292_[7], _23331_);
  buf(_23332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  buf(_37293_[7], _23333_);
  buf(_23334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  buf(_37294_[7], _23335_);
  buf(_23336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  buf(_37295_[7], _23337_);
  buf(_23338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  buf(_37296_[7], _23339_);
  buf(_23340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  buf(_37297_[7], _23341_);
  buf(_23342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  buf(_37298_[7], _23343_);
  buf(_23344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  buf(_37299_[7], _23345_);
  buf(_23348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  buf(_37300_[7], _23349_);
  buf(_23350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  buf(_37301_[7], _23351_);
  buf(_23352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  buf(_37302_[7], _23353_);
  buf(_23354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  buf(_37360_[0], _23355_);
  buf(_23356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  buf(_37360_[1], _23357_);
  buf(_23358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  buf(_37360_[2], _23359_);
  buf(_23360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  buf(_37360_[3], _23361_);
  buf(_23362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  buf(_37360_[4], _23363_);
  buf(_23364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  buf(_37360_[5], _23365_);
  buf(_23366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  buf(_37360_[6], _23367_);
  buf(_23368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  buf(_37359_[0], _23369_);
  buf(_23370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  buf(_37359_[1], _23371_);
  buf(_23372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  buf(_37359_[2], _23373_);
  buf(_23374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  buf(_37359_[3], _23375_);
  buf(_23377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  buf(_37359_[4], _23378_);
  buf(_23379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  buf(_37359_[5], _23380_);
  buf(_23381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  buf(_37359_[6], _23382_);
  buf(_23383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  buf(_37357_[0], _23384_);
  buf(_23385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  buf(_37357_[1], _23386_);
  buf(_23387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  buf(_37357_[2], _23388_);
  buf(_23389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  buf(_37357_[3], _23390_);
  buf(_23391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  buf(_37357_[4], _23392_);
  buf(_23393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  buf(_37357_[5], _23394_);
  buf(_23395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  buf(_37357_[6], _23396_);
  buf(_23397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  buf(_37356_[0], _23398_);
  buf(_23399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  buf(_37356_[1], _23400_);
  buf(_23401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  buf(_37356_[2], _23402_);
  buf(_23403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  buf(_37356_[3], _23404_);
  buf(_23405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  buf(_37356_[4], _23406_);
  buf(_23407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  buf(_37356_[5], _23408_);
  buf(_23409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  buf(_37356_[6], _23410_);
  buf(_23411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  buf(_37226_[0], _23412_);
  buf(_23413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  buf(_37226_[1], _23414_);
  buf(_23415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  buf(_37226_[2], _23416_);
  buf(_23418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  buf(_37226_[3], _23419_);
  buf(_23420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  buf(_37226_[4], _23421_);
  buf(_23422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  buf(_37226_[5], _23423_);
  buf(_23424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  buf(_37226_[6], _23425_);
  buf(_23426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  buf(_37218_[0], _23427_);
  buf(_23428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  buf(_37218_[1], _23429_);
  buf(_23430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  buf(_37218_[2], _23431_);
  buf(_23432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  buf(_37218_[3], _23433_);
  buf(_23434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  buf(_37218_[4], _23435_);
  buf(_23436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  buf(_37218_[5], _23437_);
  buf(_23438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  buf(_37218_[6], _23439_);
  buf(_23440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  buf(_37217_[0], _23441_);
  buf(_23442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  buf(_37217_[1], _23443_);
  buf(_23444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  buf(_37217_[2], _23445_);
  buf(_23446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  buf(_37217_[3], _23447_);
  buf(_23448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  buf(_37217_[4], _23449_);
  buf(_23450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  buf(_37217_[5], _23451_);
  buf(_23452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  buf(_37217_[6], _23453_);
  buf(_23454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  buf(_37216_[0], _23455_);
  buf(_23456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  buf(_37216_[1], _23457_);
  buf(_23459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  buf(_37216_[2], _23460_);
  buf(_23461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  buf(_37216_[3], _23462_);
  buf(_23463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  buf(_37216_[4], _23464_);
  buf(_23465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  buf(_37216_[5], _23466_);
  buf(_23467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  buf(_37216_[6], _23468_);
  buf(_23469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  buf(_37206_[0], _23470_);
  buf(_23471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  buf(_37206_[1], _23472_);
  buf(_23473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  buf(_37206_[2], _23474_);
  buf(_23475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  buf(_37206_[3], _23476_);
  buf(_23477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  buf(_37206_[4], _23478_);
  buf(_23479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  buf(_37206_[5], _23480_);
  buf(_23481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  buf(_37206_[6], _23482_);
  buf(_23483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  buf(_37195_[0], _23484_);
  buf(_23485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  buf(_37195_[1], _23486_);
  buf(_23487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  buf(_37195_[2], _23488_);
  buf(_23489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  buf(_37195_[3], _23490_);
  buf(_23491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  buf(_37195_[4], _23492_);
  buf(_23493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  buf(_37195_[5], _23494_);
  buf(_23495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  buf(_37195_[6], _23496_);
  buf(_23497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  buf(_37184_[0], _23498_);
  buf(_23500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  buf(_37184_[1], _23501_);
  buf(_23502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  buf(_37184_[2], _23503_);
  buf(_23504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  buf(_37184_[3], _23505_);
  buf(_23506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  buf(_37184_[4], _23507_);
  buf(_23508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  buf(_37184_[5], _23509_);
  buf(_23510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  buf(_37184_[6], _23511_);
  buf(_23512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  buf(_37365_[0], _23513_);
  buf(_23514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  buf(_37365_[1], _23515_);
  buf(_23516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  buf(_37365_[2], _23517_);
  buf(_23518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  buf(_37365_[3], _23519_);
  buf(_23520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  buf(_37365_[4], _23521_);
  buf(_23522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  buf(_37365_[5], _23523_);
  buf(_23524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  buf(_37365_[6], _23525_);
  buf(_23526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  buf(_37364_[0], _23527_);
  buf(_23528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  buf(_37364_[1], _23529_);
  buf(_23530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  buf(_37364_[2], _23531_);
  buf(_23532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  buf(_37364_[3], _23533_);
  buf(_23534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  buf(_37364_[4], _23535_);
  buf(_23536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  buf(_37364_[5], _23537_);
  buf(_23538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  buf(_37364_[6], _23539_);
  buf(_23541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  buf(_37371_[0], _23542_);
  buf(_23543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  buf(_37371_[1], _23544_);
  buf(_23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  buf(_37371_[2], _23546_);
  buf(_23547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  buf(_37371_[3], _23548_);
  buf(_23549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  buf(_37371_[4], _23550_);
  buf(_23551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  buf(_37371_[5], _23552_);
  buf(_23553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  buf(_37371_[6], _23554_);
  buf(_23555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  buf(_37373_[0], _23556_);
  buf(_23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  buf(_37373_[1], _23558_);
  buf(_23559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  buf(_37373_[2], _23560_);
  buf(_23561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  buf(_37373_[3], _23562_);
  buf(_23563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  buf(_37373_[4], _23564_);
  buf(_23565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  buf(_37373_[5], _23566_);
  buf(_23567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  buf(_37373_[6], _23568_);
  buf(_23569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  buf(_37375_[0], _23570_);
  buf(_23571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  buf(_37375_[1], _23572_);
  buf(_23573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  buf(_37375_[2], _23574_);
  buf(_23575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  buf(_37375_[3], _23576_);
  buf(_23577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  buf(_37375_[4], _23578_);
  buf(_23579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  buf(_37375_[5], _23580_);
  buf(_23582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  buf(_37375_[6], _23583_);
  buf(_23584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  buf(_37385_[0], _23585_);
  buf(_23586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  buf(_37385_[1], _23587_);
  buf(_23588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  buf(_37385_[2], _23589_);
  buf(_23590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  buf(_37385_[3], _23591_);
  buf(_23592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  buf(_37385_[4], _23593_);
  buf(_23594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  buf(_37385_[5], _23595_);
  buf(_23596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  buf(_37385_[6], _23597_);
  buf(_23598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  buf(_37393_[0], _23599_);
  buf(_23600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  buf(_37393_[1], _23601_);
  buf(_23602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  buf(_37393_[2], _23603_);
  buf(_23604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  buf(_37393_[3], _23605_);
  buf(_23606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  buf(_37393_[4], _23607_);
  buf(_23608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  buf(_37393_[5], _23609_);
  buf(_23610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  buf(_37393_[6], _23611_);
  buf(_23612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  buf(_37395_[0], _23613_);
  buf(_23614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  buf(_37395_[1], _23615_);
  buf(_23616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  buf(_37395_[2], _23617_);
  buf(_23618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  buf(_37395_[3], _23619_);
  buf(_23620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  buf(_37395_[4], _23621_);
  buf(_23623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  buf(_37395_[5], _23624_);
  buf(_23625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  buf(_37395_[6], _23626_);
  buf(_23627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  buf(_37340_[0], _23628_);
  buf(_23629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  buf(_37340_[1], _23630_);
  buf(_23631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  buf(_37340_[2], _23632_);
  buf(_23633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  buf(_37340_[3], _23634_);
  buf(_23635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  buf(_37340_[4], _23636_);
  buf(_23637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  buf(_37340_[5], _23638_);
  buf(_23639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  buf(_37340_[6], _23640_);
  buf(_23641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  buf(_37339_[0], _23642_);
  buf(_23643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  buf(_37339_[1], _23644_);
  buf(_23645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  buf(_37339_[2], _23646_);
  buf(_23647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  buf(_37339_[3], _23648_);
  buf(_23649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  buf(_37339_[4], _23650_);
  buf(_23651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  buf(_37339_[5], _23652_);
  buf(_23653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  buf(_37339_[6], _23654_);
  buf(_23655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  buf(_37341_[0], _23656_);
  buf(_23657_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  buf(_37341_[1], _23658_);
  buf(_23659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  buf(_37341_[2], _23660_);
  buf(_23661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  buf(_37341_[3], _23662_);
  buf(_23664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  buf(_37341_[4], _23665_);
  buf(_23666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  buf(_37341_[5], _23667_);
  buf(_23668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  buf(_37341_[6], _23669_);
  buf(_23670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  buf(_37338_[0], _23671_);
  buf(_23672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  buf(_37338_[1], _23673_);
  buf(_23674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  buf(_37338_[2], _23675_);
  buf(_23676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  buf(_37338_[3], _23677_);
  buf(_23678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  buf(_37338_[4], _23679_);
  buf(_23680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  buf(_37338_[5], _23681_);
  buf(_23682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  buf(_37338_[6], _23683_);
  buf(_23684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(_23686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(_23687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(_23688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(_23689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(_23690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(_23691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(_23692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  buf(_37394_[0], _23693_);
  buf(_23694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  buf(_37394_[1], _23695_);
  buf(_23696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  buf(_37394_[2], _23697_);
  buf(_23701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  buf(_37394_[3], _23702_);
  buf(_23703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  buf(_37394_[4], _23704_);
  buf(_23705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  buf(_37394_[5], _23706_);
  buf(_23707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  buf(_37394_[6], _23708_);
  buf(_23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  buf(_37302_[0], _23710_);
  buf(_23711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  buf(_37302_[1], _23712_);
  buf(_23713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  buf(_37302_[2], _23714_);
  buf(_23715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  buf(_37302_[3], _23716_);
  buf(_23717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  buf(_37302_[4], _23718_);
  buf(_23719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  buf(_37302_[5], _23720_);
  buf(_23721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  buf(_37302_[6], _23722_);
  buf(_23723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  buf(_37301_[0], _23724_);
  buf(_23725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  buf(_37301_[1], _23726_);
  buf(_23727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  buf(_37301_[2], _23728_);
  buf(_23729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  buf(_37301_[3], _23730_);
  buf(_23731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  buf(_37301_[4], _23732_);
  buf(_23733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  buf(_37301_[5], _23734_);
  buf(_23735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  buf(_37301_[6], _23736_);
  buf(_23737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  buf(_37300_[0], _23738_);
  buf(_23739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  buf(_37300_[1], _23740_);
  buf(_23742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  buf(_37300_[2], _23743_);
  buf(_23744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  buf(_37300_[3], _23745_);
  buf(_23746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  buf(_37300_[4], _23747_);
  buf(_23748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  buf(_37300_[5], _23749_);
  buf(_23750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  buf(_37300_[6], _23751_);
  buf(_23752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  buf(_37299_[0], _23753_);
  buf(_23754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  buf(_37299_[1], _23755_);
  buf(_23756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  buf(_37299_[2], _23757_);
  buf(_23758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  buf(_37299_[3], _23759_);
  buf(_23760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  buf(_37299_[4], _23761_);
  buf(_23762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  buf(_37299_[5], _23763_);
  buf(_23764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  buf(_37299_[6], _23765_);
  buf(_23766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  buf(_37298_[0], _23767_);
  buf(_23768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  buf(_37298_[1], _23769_);
  buf(_23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  buf(_37298_[2], _23771_);
  buf(_23772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  buf(_37298_[3], _23773_);
  buf(_23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  buf(_37298_[4], _23775_);
  buf(_23776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  buf(_37298_[5], _23777_);
  buf(_23778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  buf(_37298_[6], _23779_);
  buf(_23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  buf(_37297_[0], _23781_);
  buf(_23783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  buf(_37297_[1], _23784_);
  buf(_23785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  buf(_37297_[2], _23786_);
  buf(_23787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  buf(_37297_[3], _23788_);
  buf(_23789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  buf(_37297_[4], _23790_);
  buf(_23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  buf(_37297_[5], _23792_);
  buf(_23793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  buf(_37297_[6], _23794_);
  buf(_23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  buf(_37296_[0], _23796_);
  buf(_23797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  buf(_37296_[1], _23798_);
  buf(_23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  buf(_37296_[2], _23800_);
  buf(_23801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  buf(_37296_[3], _23802_);
  buf(_23803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  buf(_37296_[4], _23804_);
  buf(_23805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  buf(_37296_[5], _23806_);
  buf(_23807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  buf(_37296_[6], _23808_);
  buf(_23809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  buf(_37295_[0], _23810_);
  buf(_23811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  buf(_37295_[1], _23812_);
  buf(_23813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  buf(_37295_[2], _23814_);
  buf(_23815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  buf(_37295_[3], _23816_);
  buf(_23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  buf(_37295_[4], _23818_);
  buf(_23819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  buf(_37295_[5], _23820_);
  buf(_23821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  buf(_37295_[6], _23822_);
  buf(_23824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  buf(_37294_[0], _23825_);
  buf(_23826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  buf(_37294_[1], _23827_);
  buf(_23828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  buf(_37294_[2], _23829_);
  buf(_23830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  buf(_37294_[3], _23831_);
  buf(_23832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  buf(_37294_[4], _23833_);
  buf(_23834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  buf(_37294_[5], _23835_);
  buf(_23836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  buf(_37294_[6], _23837_);
  buf(_23838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  buf(_37293_[0], _23839_);
  buf(_23840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  buf(_37293_[1], _23841_);
  buf(_23842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  buf(_37293_[2], _23843_);
  buf(_23844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  buf(_37293_[3], _23845_);
  buf(_23846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  buf(_37293_[4], _23847_);
  buf(_23848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  buf(_37293_[5], _23849_);
  buf(_23850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  buf(_37293_[6], _23851_);
  buf(_23852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  buf(_37292_[0], _23853_);
  buf(_23854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  buf(_37292_[1], _23855_);
  buf(_23856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  buf(_37292_[2], _23857_);
  buf(_23858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  buf(_37292_[3], _23859_);
  buf(_23860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  buf(_37292_[4], _23861_);
  buf(_23862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  buf(_37292_[5], _23863_);
  buf(_23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  buf(_37292_[6], _23866_);
  buf(_23867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  buf(_37291_[0], _23868_);
  buf(_23869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  buf(_37291_[1], _23870_);
  buf(_23871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  buf(_37291_[2], _23872_);
  buf(_23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  buf(_37291_[3], _23874_);
  buf(_23875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  buf(_37291_[4], _23876_);
  buf(_23877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  buf(_37291_[5], _23878_);
  buf(_23879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  buf(_37291_[6], _23880_);
  buf(_23881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  buf(_37290_[0], _23882_);
  buf(_23883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  buf(_37290_[1], _23884_);
  buf(_23885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  buf(_37290_[2], _23886_);
  buf(_23887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  buf(_37290_[3], _23888_);
  buf(_23889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  buf(_37290_[4], _23890_);
  buf(_23891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  buf(_37290_[5], _23892_);
  buf(_23893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  buf(_37290_[6], _23894_);
  buf(_23895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  buf(_37289_[0], _23896_);
  buf(_23897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  buf(_37289_[1], _23898_);
  buf(_23899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  buf(_37289_[2], _23900_);
  buf(_23901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  buf(_37289_[3], _23902_);
  buf(_23903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  buf(_37289_[4], _23904_);
  buf(_23906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  buf(_37289_[5], _23907_);
  buf(_23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  buf(_37289_[6], _23909_);
  buf(_23910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  buf(_37288_[0], _23911_);
  buf(_23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  buf(_37288_[1], _23913_);
  buf(_23914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  buf(_37288_[2], _23915_);
  buf(_23916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  buf(_37288_[3], _23917_);
  buf(_23918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  buf(_37288_[4], _23919_);
  buf(_23920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  buf(_37288_[5], _23921_);
  buf(_23922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  buf(_37288_[6], _23923_);
  buf(_23924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  buf(_37287_[0], _23925_);
  buf(_23926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  buf(_37287_[1], _23927_);
  buf(_23928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  buf(_37287_[2], _23929_);
  buf(_23930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  buf(_37287_[3], _23931_);
  buf(_23932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  buf(_37287_[4], _23933_);
  buf(_23934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  buf(_37287_[5], _23935_);
  buf(_23936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  buf(_37287_[6], _23937_);
  buf(_23938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  buf(_37286_[0], _23939_);
  buf(_23940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  buf(_37286_[1], _23941_);
  buf(_23942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  buf(_37286_[2], _23943_);
  buf(_23944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  buf(_37286_[3], _23945_);
  buf(_23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  buf(_37286_[4], _23948_);
  buf(_23949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  buf(_37286_[5], _23950_);
  buf(_23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  buf(_37286_[6], _23952_);
  buf(_23953_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  buf(_37285_[0], _23954_);
  buf(_23955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  buf(_37285_[1], _23956_);
  buf(_23957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  buf(_37285_[2], _23958_);
  buf(_23959_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  buf(_37285_[3], _23960_);
  buf(_23961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  buf(_37285_[4], _23962_);
  buf(_23963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  buf(_37285_[5], _23964_);
  buf(_23965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  buf(_37285_[6], _23966_);
  buf(_23967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  buf(_37284_[0], _23968_);
  buf(_23969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  buf(_37284_[1], _23970_);
  buf(_23971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  buf(_37284_[2], _23972_);
  buf(_23973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  buf(_37284_[3], _23974_);
  buf(_23975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  buf(_37284_[4], _23976_);
  buf(_23977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  buf(_37284_[5], _23978_);
  buf(_23979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  buf(_37284_[6], _23980_);
  buf(_23981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  buf(_37283_[0], _23982_);
  buf(_23983_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  buf(_37283_[1], _23984_);
  buf(_23985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  buf(_37283_[2], _23986_);
  buf(_23988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  buf(_37283_[3], _23989_);
  buf(_23990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  buf(_37283_[4], _23991_);
  buf(_23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  buf(_37283_[5], _23993_);
  buf(_23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  buf(_37283_[6], _23995_);
  buf(_23996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  buf(_37282_[0], _23997_);
  buf(_23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  buf(_37282_[1], _23999_);
  buf(_24000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  buf(_37282_[2], _24001_);
  buf(_24002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  buf(_37282_[3], _24003_);
  buf(_24004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  buf(_37282_[4], _24005_);
  buf(_24006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  buf(_37282_[5], _24007_);
  buf(_24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  buf(_37282_[6], _24009_);
  buf(_24010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  buf(_37281_[0], _24011_);
  buf(_24012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  buf(_37281_[1], _24013_);
  buf(_24014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  buf(_37281_[2], _24015_);
  buf(_24016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  buf(_37281_[3], _24017_);
  buf(_24018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  buf(_37281_[4], _24019_);
  buf(_24020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  buf(_37281_[5], _24021_);
  buf(_24022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  buf(_37281_[6], _24023_);
  buf(_24024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  buf(_37280_[0], _24025_);
  buf(_24026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  buf(_37280_[1], _24027_);
  buf(_24029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  buf(_37280_[2], _24030_);
  buf(_24031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  buf(_37280_[3], _24032_);
  buf(_24033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  buf(_37280_[4], _24034_);
  buf(_24035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  buf(_37280_[5], _24036_);
  buf(_24037_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  buf(_37280_[6], _24038_);
  buf(_24039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  buf(_37279_[0], _24040_);
  buf(_24041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  buf(_37279_[1], _24042_);
  buf(_24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  buf(_37279_[2], _24044_);
  buf(_24045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  buf(_37279_[3], _24046_);
  buf(_24047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  buf(_37279_[4], _24048_);
  buf(_24049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  buf(_37279_[5], _24050_);
  buf(_24051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  buf(_37279_[6], _24052_);
  buf(_24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  buf(_37278_[0], _24054_);
  buf(_24055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  buf(_37278_[1], _24056_);
  buf(_24057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  buf(_37278_[2], _24058_);
  buf(_24059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  buf(_37278_[3], _24060_);
  buf(_24061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  buf(_37278_[4], _24062_);
  buf(_24063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  buf(_37278_[5], _24064_);
  buf(_24065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  buf(_37278_[6], _24066_);
  buf(_24067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  buf(_37277_[0], _24068_);
  buf(_24070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  buf(_37277_[1], _24071_);
  buf(_24072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  buf(_37277_[2], _24073_);
  buf(_24074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  buf(_37277_[3], _24075_);
  buf(_24076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  buf(_37277_[4], _24077_);
  buf(_24078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  buf(_37277_[5], _24079_);
  buf(_24080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  buf(_37277_[6], _24081_);
  buf(_24082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  buf(_37276_[0], _24083_);
  buf(_24084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  buf(_37276_[1], _24085_);
  buf(_24086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  buf(_37276_[2], _24087_);
  buf(_24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  buf(_37276_[3], _24089_);
  buf(_24090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  buf(_37276_[4], _24091_);
  buf(_24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  buf(_37276_[5], _24093_);
  buf(_24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  buf(_37276_[6], _24095_);
  buf(_24096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  buf(_37275_[0], _24097_);
  buf(_24098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  buf(_37275_[1], _24099_);
  buf(_24100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  buf(_37275_[2], _24101_);
  buf(_24102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  buf(_37275_[3], _24103_);
  buf(_24104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  buf(_37275_[4], _24105_);
  buf(_24106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  buf(_37275_[5], _24107_);
  buf(_24108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  buf(_37275_[6], _24109_);
  buf(_24112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  buf(_37274_[0], _24113_);
  buf(_24114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  buf(_37274_[1], _24115_);
  buf(_24116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  buf(_37274_[2], _24117_);
  buf(_24118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  buf(_37274_[3], _24119_);
  buf(_24120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  buf(_37274_[4], _24121_);
  buf(_24122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  buf(_37274_[5], _24123_);
  buf(_24124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  buf(_37274_[6], _24125_);
  buf(_24126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  buf(_37273_[0], _24127_);
  buf(_24128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  buf(_37273_[1], _24129_);
  buf(_24130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  buf(_37273_[2], _24131_);
  buf(_24132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  buf(_37273_[3], _24133_);
  buf(_24134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  buf(_37273_[4], _24135_);
  buf(_24136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  buf(_37273_[5], _24137_);
  buf(_24138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  buf(_37273_[6], _24139_);
  buf(_24140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  buf(_37272_[0], _24141_);
  buf(_24142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  buf(_37272_[1], _24143_);
  buf(_24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  buf(_37272_[2], _24145_);
  buf(_24146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  buf(_37272_[3], _24147_);
  buf(_24148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  buf(_37272_[4], _24149_);
  buf(_24150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  buf(_37272_[5], _24151_);
  buf(_24153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  buf(_37272_[6], _24154_);
  buf(_24155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  buf(_37271_[0], _24156_);
  buf(_24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  buf(_37271_[1], _24158_);
  buf(_24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  buf(_37271_[2], _24160_);
  buf(_24161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  buf(_37271_[3], _24162_);
  buf(_24163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  buf(_37271_[4], _24164_);
  buf(_24165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  buf(_37271_[5], _24166_);
  buf(_24167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  buf(_37271_[6], _24168_);
  buf(_24169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  buf(_37270_[0], _24170_);
  buf(_24171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  buf(_37270_[1], _24172_);
  buf(_24173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  buf(_37270_[2], _24174_);
  buf(_24175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  buf(_37270_[3], _24176_);
  buf(_24177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  buf(_37270_[4], _24178_);
  buf(_24179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  buf(_37270_[5], _24180_);
  buf(_24181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  buf(_37270_[6], _24182_);
  buf(_24183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  buf(_37269_[0], _24184_);
  buf(_24185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  buf(_37269_[1], _24186_);
  buf(_24187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  buf(_37269_[2], _24188_);
  buf(_24189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  buf(_37269_[3], _24190_);
  buf(_24191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  buf(_37269_[4], _24192_);
  buf(_24194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  buf(_37269_[5], _24195_);
  buf(_24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  buf(_37269_[6], _24197_);
  buf(_24198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  buf(_37268_[0], _24199_);
  buf(_24200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  buf(_37268_[1], _24201_);
  buf(_24202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  buf(_37268_[2], _24203_);
  buf(_24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  buf(_37268_[3], _24205_);
  buf(_24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  buf(_37268_[4], _24207_);
  buf(_24208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  buf(_37268_[5], _24209_);
  buf(_24210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  buf(_37268_[6], _24211_);
  buf(_24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  buf(_37267_[0], _24213_);
  buf(_24214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  buf(_37267_[1], _24215_);
  buf(_24216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  buf(_37267_[2], _24217_);
  buf(_24218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  buf(_37267_[3], _24219_);
  buf(_24220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  buf(_37267_[4], _24221_);
  buf(_24222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  buf(_37267_[5], _24223_);
  buf(_24224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  buf(_37267_[6], _24225_);
  buf(_24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  buf(_37266_[0], _24227_);
  buf(_24228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  buf(_37266_[1], _24229_);
  buf(_24230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  buf(_37266_[2], _24231_);
  buf(_24232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  buf(_37266_[3], _24233_);
  buf(_24235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  buf(_37266_[4], _24236_);
  buf(_24237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  buf(_37266_[5], _24238_);
  buf(_24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  buf(_37266_[6], _24240_);
  buf(_24241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  buf(_37265_[0], _24242_);
  buf(_24243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  buf(_37265_[1], _24244_);
  buf(_24245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  buf(_37265_[2], _24246_);
  buf(_24247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  buf(_37265_[3], _24248_);
  buf(_24249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  buf(_37265_[4], _24250_);
  buf(_24251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  buf(_37265_[5], _24252_);
  buf(_24253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  buf(_37265_[6], _24254_);
  buf(_24255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  buf(_37264_[0], _24256_);
  buf(_24257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  buf(_37264_[1], _24258_);
  buf(_24259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  buf(_37264_[2], _24260_);
  buf(_24261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  buf(_37264_[3], _24262_);
  buf(_24263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  buf(_37264_[4], _24264_);
  buf(_24265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  buf(_37264_[5], _24266_);
  buf(_24267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  buf(_37264_[6], _24268_);
  buf(_24269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  buf(_37263_[0], _24270_);
  buf(_24271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  buf(_37263_[1], _24272_);
  buf(_24273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  buf(_37263_[2], _24274_);
  buf(_24276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  buf(_37263_[3], _24277_);
  buf(_24278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  buf(_37263_[4], _24279_);
  buf(_24280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  buf(_37263_[5], _24281_);
  buf(_24282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  buf(_37263_[6], _24283_);
  buf(_24284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  buf(_37262_[0], _24285_);
  buf(_24286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  buf(_37262_[1], _24287_);
  buf(_24288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  buf(_37262_[2], _24289_);
  buf(_24290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  buf(_37262_[3], _24291_);
  buf(_24292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  buf(_37262_[4], _24293_);
  buf(_24294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  buf(_37262_[5], _24295_);
  buf(_24296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  buf(_37262_[6], _24297_);
  buf(_24298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  buf(_37261_[0], _24299_);
  buf(_24300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  buf(_37261_[1], _24301_);
  buf(_24302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  buf(_37261_[2], _24303_);
  buf(_24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  buf(_37261_[3], _24305_);
  buf(_24306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  buf(_37261_[4], _24307_);
  buf(_24308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  buf(_37261_[5], _24309_);
  buf(_24310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  buf(_37261_[6], _24311_);
  buf(_24312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  buf(_37260_[0], _24313_);
  buf(_24314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  buf(_37260_[1], _24315_);
  buf(_24317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  buf(_37260_[2], _24318_);
  buf(_24319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  buf(_37260_[3], _24320_);
  buf(_24321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  buf(_37260_[4], _24322_);
  buf(_24323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  buf(_37260_[5], _24324_);
  buf(_24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  buf(_37260_[6], _24326_);
  buf(_24327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  buf(_37259_[0], _24328_);
  buf(_24329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  buf(_37259_[1], _24330_);
  buf(_24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  buf(_37259_[2], _24332_);
  buf(_24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  buf(_37259_[3], _24334_);
  buf(_24335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  buf(_37259_[4], _24336_);
  buf(_24337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  buf(_37259_[5], _24338_);
  buf(_24339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  buf(_37259_[6], _24340_);
  buf(_24341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  buf(_37258_[0], _24342_);
  buf(_24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  buf(_37258_[1], _24344_);
  buf(_24345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  buf(_37258_[2], _24346_);
  buf(_24347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  buf(_37258_[3], _24348_);
  buf(_24349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  buf(_37258_[4], _24350_);
  buf(_24351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  buf(_37258_[5], _24352_);
  buf(_24353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  buf(_37258_[6], _24354_);
  buf(_24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  buf(_37257_[0], _24356_);
  buf(_24358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  buf(_37257_[1], _24359_);
  buf(_24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  buf(_37257_[2], _24361_);
  buf(_24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  buf(_37257_[3], _24363_);
  buf(_24364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  buf(_37257_[4], _24365_);
  buf(_24366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  buf(_37257_[5], _24367_);
  buf(_24368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  buf(_37257_[6], _24369_);
  buf(_24370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  buf(_37256_[0], _24371_);
  buf(_24372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  buf(_37256_[1], _24373_);
  buf(_24374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  buf(_37256_[2], _24375_);
  buf(_24376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  buf(_37256_[3], _24377_);
  buf(_24378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  buf(_37256_[4], _24379_);
  buf(_24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  buf(_37256_[5], _24381_);
  buf(_24382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  buf(_37256_[6], _24383_);
  buf(_24384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  buf(_37255_[0], _24385_);
  buf(_24386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  buf(_37255_[1], _24387_);
  buf(_24388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  buf(_37255_[2], _24389_);
  buf(_24390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  buf(_37255_[3], _24391_);
  buf(_24392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  buf(_37255_[4], _24393_);
  buf(_24394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  buf(_37255_[5], _24395_);
  buf(_24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  buf(_37255_[6], _24397_);
  buf(_24399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  buf(_37254_[0], _24400_);
  buf(_24401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  buf(_37254_[1], _24402_);
  buf(_24403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  buf(_37254_[2], _24404_);
  buf(_24405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  buf(_37254_[3], _24406_);
  buf(_24407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  buf(_37254_[4], _24408_);
  buf(_24409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  buf(_37254_[5], _24410_);
  buf(_24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  buf(_37254_[6], _24412_);
  buf(_24413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  buf(_37253_[0], _24414_);
  buf(_24415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  buf(_37253_[1], _24416_);
  buf(_24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  buf(_37253_[2], _24418_);
  buf(_24419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  buf(_37253_[3], _24420_);
  buf(_24421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  buf(_37253_[4], _24422_);
  buf(_24423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  buf(_37253_[5], _24424_);
  buf(_24425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  buf(_37253_[6], _24426_);
  buf(_24427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  buf(_37252_[0], _24428_);
  buf(_24429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  buf(_37252_[1], _24430_);
  buf(_24431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  buf(_37252_[2], _24432_);
  buf(_24433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  buf(_37252_[3], _24434_);
  buf(_24435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  buf(_37252_[4], _24436_);
  buf(_24437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  buf(_37252_[5], _24438_);
  buf(_24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  buf(_37252_[6], _24441_);
  buf(_24442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  buf(_37251_[0], _24443_);
  buf(_24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  buf(_37251_[1], _24445_);
  buf(_24446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  buf(_37251_[2], _24447_);
  buf(_24448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  buf(_37251_[3], _24449_);
  buf(_24450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  buf(_37251_[4], _24451_);
  buf(_24452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  buf(_37251_[5], _24453_);
  buf(_24454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  buf(_37251_[6], _24455_);
  buf(_24456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  buf(_37250_[0], _24457_);
  buf(_24458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  buf(_37250_[1], _24459_);
  buf(_24460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  buf(_37250_[2], _24461_);
  buf(_24462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  buf(_37250_[3], _24463_);
  buf(_24464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  buf(_37250_[4], _24465_);
  buf(_24466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  buf(_37250_[5], _24467_);
  buf(_24468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  buf(_37250_[6], _24469_);
  buf(_24470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  buf(_37249_[0], _24471_);
  buf(_24472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  buf(_37249_[1], _24473_);
  buf(_24474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  buf(_37249_[2], _24475_);
  buf(_24476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  buf(_37249_[3], _24477_);
  buf(_24478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  buf(_37249_[4], _24479_);
  buf(_24481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  buf(_37249_[5], _24482_);
  buf(_24483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  buf(_37249_[6], _24484_);
  buf(_24485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  buf(_37248_[0], _24486_);
  buf(_24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  buf(_37248_[1], _24488_);
  buf(_24489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  buf(_37248_[2], _24490_);
  buf(_24491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  buf(_37248_[3], _24492_);
  buf(_24493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  buf(_37248_[4], _24494_);
  buf(_24495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  buf(_37248_[5], _24496_);
  buf(_24497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  buf(_37248_[6], _24498_);
  buf(_24499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  buf(_37247_[0], _24500_);
  buf(_24501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  buf(_37247_[1], _24502_);
  buf(_24503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  buf(_37247_[2], _24504_);
  buf(_24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  buf(_37247_[3], _24506_);
  buf(_24507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  buf(_37247_[4], _24508_);
  buf(_24509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  buf(_37247_[5], _24510_);
  buf(_24511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  buf(_37247_[6], _24512_);
  buf(_24513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  buf(_37246_[0], _24514_);
  buf(_24515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  buf(_37246_[1], _24516_);
  buf(_24517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  buf(_37246_[2], _24518_);
  buf(_24519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  buf(_37246_[3], _24520_);
  buf(_24523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  buf(_37246_[4], _24524_);
  buf(_24525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  buf(_37246_[5], _24526_);
  buf(_24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  buf(_37246_[6], _24528_);
  buf(_24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  buf(_37245_[0], _24530_);
  buf(_24531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  buf(_37245_[1], _24532_);
  buf(_24533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  buf(_37245_[2], _24534_);
  buf(_24535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  buf(_37245_[3], _24536_);
  buf(_24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  buf(_37245_[4], _24538_);
  buf(_24539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  buf(_37245_[5], _24540_);
  buf(_24541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  buf(_37245_[6], _24542_);
  buf(_24543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  buf(_37244_[0], _24544_);
  buf(_24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  buf(_37244_[1], _24546_);
  buf(_24547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  buf(_37244_[2], _24548_);
  buf(_24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  buf(_37244_[3], _24550_);
  buf(_24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  buf(_37244_[4], _24552_);
  buf(_24553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  buf(_37244_[5], _24554_);
  buf(_24555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  buf(_37244_[6], _24556_);
  buf(_24557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  buf(_37243_[0], _24558_);
  buf(_24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  buf(_37243_[1], _24560_);
  buf(_24561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  buf(_37243_[2], _24562_);
  buf(_24564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  buf(_37243_[3], _24565_);
  buf(_24566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  buf(_37243_[4], _24567_);
  buf(_24568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  buf(_37243_[5], _24569_);
  buf(_24570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  buf(_37243_[6], _24571_);
  buf(_24572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  buf(_37242_[0], _24573_);
  buf(_24574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  buf(_37242_[1], _24575_);
  buf(_24576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  buf(_37242_[2], _24577_);
  buf(_24578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  buf(_37242_[3], _24579_);
  buf(_24580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  buf(_37242_[4], _24581_);
  buf(_24582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  buf(_37242_[5], _24583_);
  buf(_24584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  buf(_37242_[6], _24585_);
  buf(_24586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  buf(_37241_[0], _24587_);
  buf(_24588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  buf(_37241_[1], _24589_);
  buf(_24590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  buf(_37241_[2], _24591_);
  buf(_24592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  buf(_37241_[3], _24593_);
  buf(_24594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  buf(_37241_[4], _24595_);
  buf(_24596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  buf(_37241_[5], _24597_);
  buf(_24598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  buf(_37241_[6], _24599_);
  buf(_24600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  buf(_37240_[0], _24601_);
  buf(_24602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  buf(_37240_[1], _24603_);
  buf(_24605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  buf(_37240_[2], _24606_);
  buf(_24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  buf(_37240_[3], _24608_);
  buf(_24609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  buf(_37240_[4], _24610_);
  buf(_24611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  buf(_37240_[5], _24612_);
  buf(_24613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  buf(_37240_[6], _24614_);
  buf(_24615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  buf(_37239_[0], _24616_);
  buf(_24617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  buf(_37239_[1], _24618_);
  buf(_24619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  buf(_37239_[2], _24620_);
  buf(_24621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  buf(_37239_[3], _24622_);
  buf(_24623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  buf(_37239_[4], _24624_);
  buf(_24625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  buf(_37239_[5], _24626_);
  buf(_24627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  buf(_37239_[6], _24628_);
  buf(_24629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  buf(_37238_[0], _24630_);
  buf(_24631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  buf(_37238_[1], _24632_);
  buf(_24633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  buf(_37238_[2], _24634_);
  buf(_24635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  buf(_37238_[3], _24636_);
  buf(_24637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  buf(_37238_[4], _24638_);
  buf(_24639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  buf(_37238_[5], _24640_);
  buf(_24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  buf(_37238_[6], _24642_);
  buf(_24643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  buf(_37237_[0], _24644_);
  buf(_24646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  buf(_37237_[1], _24647_);
  buf(_24648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  buf(_37237_[2], _24649_);
  buf(_24650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  buf(_37237_[3], _24651_);
  buf(_24652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  buf(_37237_[4], _24653_);
  buf(_24654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  buf(_37237_[5], _24655_);
  buf(_24656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  buf(_37237_[6], _24657_);
  buf(_24658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  buf(_37236_[0], _24659_);
  buf(_24660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  buf(_37236_[1], _24661_);
  buf(_24662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  buf(_37236_[2], _24663_);
  buf(_24664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  buf(_37236_[3], _24665_);
  buf(_24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  buf(_37236_[4], _24667_);
  buf(_24668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  buf(_37236_[5], _24669_);
  buf(_24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  buf(_37236_[6], _24671_);
  buf(_24672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  buf(_37235_[0], _24673_);
  buf(_24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  buf(_37235_[1], _24675_);
  buf(_24676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  buf(_37235_[2], _24677_);
  buf(_24678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  buf(_37235_[3], _24679_);
  buf(_24680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  buf(_37235_[4], _24681_);
  buf(_24682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  buf(_37235_[5], _24683_);
  buf(_24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  buf(_37235_[6], _24685_);
  buf(_24687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  buf(_37234_[0], _24688_);
  buf(_24689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  buf(_37234_[1], _24690_);
  buf(_24691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  buf(_37234_[2], _24692_);
  buf(_24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  buf(_37234_[3], _24694_);
  buf(_24695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  buf(_37234_[4], _24696_);
  buf(_24697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  buf(_37234_[5], _24698_);
  buf(_24699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  buf(_37234_[6], _24700_);
  buf(_24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  buf(_37233_[0], _24702_);
  buf(_24703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  buf(_37233_[1], _24704_);
  buf(_24705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  buf(_37233_[2], _24706_);
  buf(_24707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  buf(_37233_[3], _24708_);
  buf(_24709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  buf(_37233_[4], _24710_);
  buf(_24711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  buf(_37233_[5], _24712_);
  buf(_24713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  buf(_37233_[6], _24714_);
  buf(_24715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  buf(_37232_[0], _24716_);
  buf(_24717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  buf(_37232_[1], _24718_);
  buf(_24719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  buf(_37232_[2], _24720_);
  buf(_24721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  buf(_37232_[3], _24722_);
  buf(_24723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  buf(_37232_[4], _24724_);
  buf(_24725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  buf(_37232_[5], _24726_);
  buf(_24728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  buf(_37232_[6], _24729_);
  buf(_24730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  buf(_37231_[0], _24731_);
  buf(_24732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  buf(_37231_[1], _24733_);
  buf(_24734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  buf(_37231_[2], _24735_);
  buf(_24736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  buf(_37231_[3], _24737_);
  buf(_24738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  buf(_37231_[4], _24739_);
  buf(_24740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  buf(_37231_[5], _24741_);
  buf(_24742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  buf(_37231_[6], _24743_);
  buf(_24744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  buf(_37230_[0], _24745_);
  buf(_24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  buf(_37230_[1], _24747_);
  buf(_24748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  buf(_37230_[2], _24749_);
  buf(_24750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  buf(_37230_[3], _24751_);
  buf(_24752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  buf(_37230_[4], _24753_);
  buf(_24754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  buf(_37230_[5], _24755_);
  buf(_24756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  buf(_37230_[6], _24757_);
  buf(_24758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  buf(_37229_[0], _24759_);
  buf(_24760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  buf(_37229_[1], _24761_);
  buf(_24762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  buf(_37229_[2], _24763_);
  buf(_24764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  buf(_37229_[3], _24765_);
  buf(_24766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  buf(_37229_[4], _24767_);
  buf(_24769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  buf(_37229_[5], _24770_);
  buf(_24771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  buf(_37229_[6], _24772_);
  buf(_24773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  buf(_37228_[0], _24774_);
  buf(_24775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  buf(_37228_[1], _24776_);
  buf(_24777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  buf(_37228_[2], _24778_);
  buf(_24779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  buf(_37228_[3], _24780_);
  buf(_24781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  buf(_37228_[4], _24782_);
  buf(_24783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  buf(_37228_[5], _24784_);
  buf(_24785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  buf(_37228_[6], _24786_);
  buf(_24787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  buf(_37227_[0], _24788_);
  buf(_24789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  buf(_37227_[1], _24790_);
  buf(_24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  buf(_37227_[2], _24792_);
  buf(_24793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  buf(_37227_[3], _24794_);
  buf(_24795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  buf(_37227_[4], _24796_);
  buf(_24797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  buf(_37227_[5], _24798_);
  buf(_24799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  buf(_37227_[6], _24800_);
  buf(_24801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  buf(_37225_[0], _24802_);
  buf(_24803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  buf(_37225_[1], _24804_);
  buf(_24805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  buf(_37225_[2], _24806_);
  buf(_24807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  buf(_37225_[3], _24808_);
  buf(_24810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  buf(_37225_[4], _24811_);
  buf(_24812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  buf(_37225_[5], _24813_);
  buf(_24814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  buf(_37225_[6], _24815_);
  buf(_24816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  buf(_37224_[0], _24817_);
  buf(_24818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  buf(_37224_[1], _24819_);
  buf(_24820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  buf(_37224_[2], _24821_);
  buf(_24822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  buf(_37224_[3], _24823_);
  buf(_24824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  buf(_37224_[4], _24825_);
  buf(_24826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  buf(_37224_[5], _24827_);
  buf(_24828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  buf(_37224_[6], _24829_);
  buf(_24830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  buf(_37223_[0], _24831_);
  buf(_24832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  buf(_37223_[1], _24833_);
  buf(_24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  buf(_37223_[2], _24835_);
  buf(_24836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  buf(_37223_[3], _24837_);
  buf(_24838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  buf(_37223_[4], _24839_);
  buf(_24840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  buf(_37223_[5], _24841_);
  buf(_24842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  buf(_37223_[6], _24843_);
  buf(_24844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  buf(_37222_[0], _24845_);
  buf(_24846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  buf(_37222_[1], _24847_);
  buf(_24848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  buf(_37222_[2], _24849_);
  buf(_24851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  buf(_37222_[3], _24852_);
  buf(_24853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  buf(_37222_[4], _24854_);
  buf(_24855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  buf(_37222_[5], _24856_);
  buf(_24857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  buf(_37222_[6], _24858_);
  buf(_24859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  buf(_37221_[0], _24860_);
  buf(_24861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  buf(_37221_[1], _24862_);
  buf(_24863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  buf(_37221_[2], _24864_);
  buf(_24865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  buf(_37221_[3], _24866_);
  buf(_24867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  buf(_37221_[4], _24868_);
  buf(_24869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  buf(_37221_[5], _24870_);
  buf(_24871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  buf(_37221_[6], _24872_);
  buf(_24873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  buf(_37220_[0], _24874_);
  buf(_24875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  buf(_37220_[1], _24876_);
  buf(_24877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  buf(_37220_[2], _24878_);
  buf(_24879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  buf(_37220_[3], _24880_);
  buf(_24881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  buf(_37220_[4], _24882_);
  buf(_24883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  buf(_37220_[5], _24884_);
  buf(_24885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  buf(_37220_[6], _24886_);
  buf(_24887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  buf(_37219_[0], _24888_);
  buf(_24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  buf(_37219_[1], _24890_);
  buf(_24892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  buf(_37219_[2], _24893_);
  buf(_24894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  buf(_37219_[3], _24895_);
  buf(_24896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  buf(_37219_[4], _24897_);
  buf(_24898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  buf(_37219_[5], _24899_);
  buf(_24900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  buf(_37219_[6], _24901_);
  buf(_24902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  buf(_37355_[0], _24903_);
  buf(_24904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  buf(_37355_[1], _24905_);
  buf(_24906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  buf(_37355_[2], _24907_);
  buf(_24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  buf(_37355_[3], _24909_);
  buf(_24910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  buf(_37355_[4], _24911_);
  buf(_24912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  buf(_37355_[5], _24913_);
  buf(_24914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  buf(_37355_[6], _24915_);
  buf(_24916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  buf(_37354_[0], _24917_);
  buf(_24918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  buf(_37354_[1], _24919_);
  buf(_24920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  buf(_37354_[2], _24921_);
  buf(_24922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  buf(_37354_[3], _24923_);
  buf(_24924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  buf(_37354_[4], _24925_);
  buf(_24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  buf(_37354_[5], _24927_);
  buf(_24928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  buf(_37354_[6], _24929_);
  buf(_24930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  buf(_37353_[0], _24931_);
  buf(_24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  buf(_37353_[1], _24935_);
  buf(_24936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  buf(_37353_[2], _24937_);
  buf(_24938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  buf(_37353_[3], _24939_);
  buf(_24940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  buf(_37353_[4], _24941_);
  buf(_24942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  buf(_37353_[5], _24943_);
  buf(_24944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  buf(_37353_[6], _24945_);
  buf(_24946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  buf(_37352_[0], _24947_);
  buf(_24948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  buf(_37352_[1], _24949_);
  buf(_24950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  buf(_37352_[2], _24951_);
  buf(_24952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  buf(_37352_[3], _24953_);
  buf(_24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  buf(_37352_[4], _24955_);
  buf(_24956_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  buf(_37352_[5], _24957_);
  buf(_24958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  buf(_37352_[6], _24959_);
  buf(_24960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  buf(_37351_[0], _24961_);
  buf(_24962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  buf(_37351_[1], _24963_);
  buf(_24964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  buf(_37351_[2], _24965_);
  buf(_24966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  buf(_37351_[3], _24967_);
  buf(_24968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  buf(_37351_[4], _24969_);
  buf(_24970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  buf(_37351_[5], _24971_);
  buf(_24972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  buf(_37351_[6], _24973_);
  buf(_24975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  buf(_37350_[0], _24976_);
  buf(_24977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  buf(_37350_[1], _24978_);
  buf(_24979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  buf(_37350_[2], _24980_);
  buf(_24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  buf(_37350_[3], _24982_);
  buf(_24983_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  buf(_37350_[4], _24984_);
  buf(_24985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  buf(_37350_[5], _24986_);
  buf(_24987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  buf(_37350_[6], _24988_);
  buf(_24989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  buf(_37349_[0], _24990_);
  buf(_24991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  buf(_37349_[1], _24992_);
  buf(_24993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  buf(_37349_[2], _24994_);
  buf(_24995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  buf(_37349_[3], _24996_);
  buf(_24997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  buf(_37349_[4], _24998_);
  buf(_24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  buf(_37349_[5], _25000_);
  buf(_25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  buf(_37349_[6], _25002_);
  buf(_25003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  buf(_37348_[0], _25004_);
  buf(_25005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  buf(_37348_[1], _25006_);
  buf(_25007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  buf(_37348_[2], _25008_);
  buf(_25009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  buf(_37348_[3], _25010_);
  buf(_25011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  buf(_37348_[4], _25012_);
  buf(_25013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  buf(_37348_[5], _25014_);
  buf(_25016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  buf(_37348_[6], _25017_);
  buf(_25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  buf(_37347_[0], _25019_);
  buf(_25020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  buf(_37347_[1], _25021_);
  buf(_25022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  buf(_37347_[2], _25023_);
  buf(_25024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  buf(_37347_[3], _25025_);
  buf(_25026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  buf(_37347_[4], _25027_);
  buf(_25028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  buf(_37347_[5], _25029_);
  buf(_25030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  buf(_37347_[6], _25031_);
  buf(_25032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  buf(_37346_[0], _25033_);
  buf(_25034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  buf(_37346_[1], _25035_);
  buf(_25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  buf(_37346_[2], _25037_);
  buf(_25038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  buf(_37346_[3], _25039_);
  buf(_25040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  buf(_37346_[4], _25041_);
  buf(_25042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  buf(_37346_[5], _25043_);
  buf(_25044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  buf(_37346_[6], _25045_);
  buf(_25046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  buf(_37345_[0], _25047_);
  buf(_25048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  buf(_37345_[1], _25049_);
  buf(_25050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  buf(_37345_[2], _25051_);
  buf(_25052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  buf(_37345_[3], _25053_);
  buf(_25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  buf(_37345_[4], _25055_);
  buf(_25057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  buf(_37345_[5], _25058_);
  buf(_25059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  buf(_37345_[6], _25060_);
  buf(_25061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  buf(_37344_[0], _25062_);
  buf(_25063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  buf(_37344_[1], _25064_);
  buf(_25065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  buf(_37344_[2], _25066_);
  buf(_25067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  buf(_37344_[3], _25068_);
  buf(_25069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  buf(_37344_[4], _25070_);
  buf(_25071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  buf(_37344_[5], _25072_);
  buf(_25073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  buf(_37344_[6], _25074_);
  buf(_25075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  buf(_37343_[0], _25076_);
  buf(_25077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  buf(_37343_[1], _25078_);
  buf(_25079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  buf(_37343_[2], _25080_);
  buf(_25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  buf(_37343_[3], _25082_);
  buf(_25083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  buf(_37343_[4], _25084_);
  buf(_25085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  buf(_37343_[5], _25086_);
  buf(_25087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  buf(_37343_[6], _25088_);
  buf(_25089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  buf(_37342_[0], _25090_);
  buf(_25091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  buf(_37342_[1], _25092_);
  buf(_25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  buf(_37342_[2], _25094_);
  buf(_25095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  buf(_37342_[3], _25096_);
  buf(_25098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  buf(_37342_[4], _25099_);
  buf(_25100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  buf(_37342_[5], _25101_);
  buf(_25102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  buf(_37342_[6], _25103_);
  buf(_25104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  buf(_37337_[0], _25105_);
  buf(_25106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  buf(_37337_[1], _25107_);
  buf(_25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  buf(_37337_[2], _25109_);
  buf(_25110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  buf(_37337_[3], _25111_);
  buf(_25112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  buf(_37337_[4], _25113_);
  buf(_25114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  buf(_37337_[5], _25115_);
  buf(_25116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  buf(_37337_[6], _25117_);
  buf(_25118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  buf(_37336_[0], _25119_);
  buf(_25120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  buf(_37336_[1], _25121_);
  buf(_25122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  buf(_37336_[2], _25123_);
  buf(_25124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  buf(_37336_[3], _25125_);
  buf(_25126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  buf(_37336_[4], _25127_);
  buf(_25128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  buf(_37336_[5], _25129_);
  buf(_25130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  buf(_37336_[6], _25131_);
  buf(_25132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  buf(_37335_[0], _25133_);
  buf(_25134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  buf(_37335_[1], _25135_);
  buf(_25136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  buf(_37335_[2], _25137_);
  buf(_25139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  buf(_37335_[3], _25140_);
  buf(_25141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  buf(_37335_[4], _25142_);
  buf(_25143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  buf(_37335_[5], _25144_);
  buf(_25145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  buf(_37335_[6], _25146_);
  buf(_25147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  buf(_37334_[0], _25148_);
  buf(_25149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  buf(_37334_[1], _25150_);
  buf(_25151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  buf(_37334_[2], _25152_);
  buf(_25153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  buf(_37334_[3], _25154_);
  buf(_25155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  buf(_37334_[4], _25156_);
  buf(_25157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  buf(_37334_[5], _25158_);
  buf(_25159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  buf(_37334_[6], _25160_);
  buf(_25161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  buf(_37333_[0], _25162_);
  buf(_25163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  buf(_37333_[1], _25164_);
  buf(_25165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  buf(_37333_[2], _25166_);
  buf(_25167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  buf(_37333_[3], _25168_);
  buf(_25169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  buf(_37333_[4], _25170_);
  buf(_25171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  buf(_37333_[5], _25172_);
  buf(_25173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  buf(_37333_[6], _25174_);
  buf(_25175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  buf(_37332_[0], _25176_);
  buf(_25177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  buf(_37332_[1], _25178_);
  buf(_25180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  buf(_37332_[2], _25181_);
  buf(_25182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  buf(_37332_[3], _25183_);
  buf(_25184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  buf(_37332_[4], _25185_);
  buf(_25186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  buf(_37332_[5], _25187_);
  buf(_25188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  buf(_37332_[6], _25189_);
  buf(_25190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  buf(_37215_[0], _25191_);
  buf(_25192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  buf(_37215_[1], _25193_);
  buf(_25194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  buf(_37215_[2], _25195_);
  buf(_25196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  buf(_37215_[3], _25197_);
  buf(_25198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  buf(_37215_[4], _25199_);
  buf(_25200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  buf(_37215_[5], _25201_);
  buf(_25202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  buf(_37215_[6], _25203_);
  buf(_25204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  buf(_37214_[0], _25205_);
  buf(_25206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  buf(_37214_[1], _25207_);
  buf(_25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  buf(_37214_[2], _25209_);
  buf(_25210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  buf(_37214_[3], _25211_);
  buf(_25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  buf(_37214_[4], _25213_);
  buf(_25214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  buf(_37214_[5], _25215_);
  buf(_25216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  buf(_37214_[6], _25217_);
  buf(_25218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  buf(_37213_[0], _25219_);
  buf(_25221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  buf(_37213_[1], _25222_);
  buf(_25223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  buf(_37213_[2], _25224_);
  buf(_25225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  buf(_37213_[3], _25226_);
  buf(_25227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  buf(_37213_[4], _25228_);
  buf(_25229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  buf(_37213_[5], _25230_);
  buf(_25231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  buf(_37213_[6], _25232_);
  buf(_25233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  buf(_37212_[0], _25234_);
  buf(_25235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  buf(_37212_[1], _25236_);
  buf(_25237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  buf(_37212_[2], _25238_);
  buf(_25239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  buf(_37212_[3], _25240_);
  buf(_25241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  buf(_37212_[4], _25242_);
  buf(_25243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  buf(_37212_[5], _25244_);
  buf(_25245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  buf(_37212_[6], _25246_);
  buf(_25247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  buf(_37211_[0], _25248_);
  buf(_25249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  buf(_37211_[1], _25250_);
  buf(_25251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  buf(_37211_[2], _25252_);
  buf(_25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  buf(_37211_[3], _25254_);
  buf(_25255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  buf(_37211_[4], _25256_);
  buf(_25257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  buf(_37211_[5], _25258_);
  buf(_25259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  buf(_37211_[6], _25260_);
  buf(_25262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  buf(_37210_[0], _25263_);
  buf(_25264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  buf(_37210_[1], _25265_);
  buf(_25266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  buf(_37210_[2], _25267_);
  buf(_25268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  buf(_37210_[3], _25269_);
  buf(_25270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  buf(_37210_[4], _25271_);
  buf(_25272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  buf(_37210_[5], _25273_);
  buf(_25274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  buf(_37210_[6], _25275_);
  buf(_25276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  buf(_37209_[0], _25277_);
  buf(_25278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  buf(_37209_[1], _25279_);
  buf(_25280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  buf(_37209_[2], _25281_);
  buf(_25282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  buf(_37209_[3], _25283_);
  buf(_25284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  buf(_37209_[4], _25285_);
  buf(_25286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  buf(_37209_[5], _25287_);
  buf(_25288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  buf(_37209_[6], _25289_);
  buf(_25290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  buf(_37208_[0], _25291_);
  buf(_25292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  buf(_37208_[1], _25293_);
  buf(_25294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  buf(_37208_[2], _25295_);
  buf(_25296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  buf(_37208_[3], _25297_);
  buf(_25298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  buf(_37208_[4], _25299_);
  buf(_25300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  buf(_37208_[5], _25301_);
  buf(_25303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  buf(_37208_[6], _25304_);
  buf(_25305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  buf(_37207_[0], _25306_);
  buf(_25307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  buf(_37207_[1], _25308_);
  buf(_25309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  buf(_37207_[2], _25310_);
  buf(_25311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  buf(_37207_[3], _25312_);
  buf(_25313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  buf(_37207_[4], _25314_);
  buf(_25315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  buf(_37207_[5], _25316_);
  buf(_25317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  buf(_37207_[6], _25318_);
  buf(_25319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  buf(_37205_[0], _25320_);
  buf(_25321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  buf(_37205_[1], _25322_);
  buf(_25323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  buf(_37205_[2], _25324_);
  buf(_25325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  buf(_37205_[3], _25326_);
  buf(_25327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  buf(_37205_[4], _25328_);
  buf(_25329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  buf(_37205_[5], _25330_);
  buf(_25331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  buf(_37205_[6], _25332_);
  buf(_25333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  buf(_37204_[0], _25334_);
  buf(_25335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  buf(_37204_[1], _25336_);
  buf(_25337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  buf(_37204_[2], _25338_);
  buf(_25339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  buf(_37204_[3], _25340_);
  buf(_25341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  buf(_37204_[4], _25342_);
  buf(_25345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  buf(_37204_[5], _25346_);
  buf(_25347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  buf(_37204_[6], _25348_);
  buf(_25349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  buf(_37203_[0], _25350_);
  buf(_25351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  buf(_37203_[1], _25352_);
  buf(_25353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  buf(_37203_[2], _25354_);
  buf(_25355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  buf(_37203_[3], _25356_);
  buf(_25357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  buf(_37203_[4], _25358_);
  buf(_25359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  buf(_37203_[5], _25360_);
  buf(_25361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  buf(_37203_[6], _25362_);
  buf(_25363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  buf(_37202_[0], _25364_);
  buf(_25365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  buf(_37202_[1], _25366_);
  buf(_25367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  buf(_37202_[2], _25368_);
  buf(_25369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  buf(_37202_[3], _25370_);
  buf(_25371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  buf(_37202_[4], _25372_);
  buf(_25373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  buf(_37202_[5], _25374_);
  buf(_25375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  buf(_37202_[6], _25376_);
  buf(_25377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  buf(_37201_[0], _25378_);
  buf(_25379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  buf(_37201_[1], _25380_);
  buf(_25381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  buf(_37201_[2], _25382_);
  buf(_25383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  buf(_37201_[3], _25384_);
  buf(_25386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  buf(_37201_[4], _25387_);
  buf(_25388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  buf(_37201_[5], _25389_);
  buf(_25390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  buf(_37201_[6], _25391_);
  buf(_25392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  buf(_37200_[0], _25393_);
  buf(_25394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  buf(_37200_[1], _25395_);
  buf(_25396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  buf(_37200_[2], _25397_);
  buf(_25398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  buf(_37200_[3], _25399_);
  buf(_25400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  buf(_37200_[4], _25401_);
  buf(_25402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  buf(_37200_[5], _25403_);
  buf(_25404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  buf(_37200_[6], _25405_);
  buf(_25406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  buf(_37199_[0], _25407_);
  buf(_25408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  buf(_37199_[1], _25409_);
  buf(_25410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  buf(_37199_[2], _25411_);
  buf(_25412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  buf(_37199_[3], _25413_);
  buf(_25414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  buf(_37199_[4], _25415_);
  buf(_25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  buf(_37199_[5], _25417_);
  buf(_25418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  buf(_37199_[6], _25419_);
  buf(_25420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  buf(_37198_[0], _25421_);
  buf(_25422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  buf(_37198_[1], _25423_);
  buf(_25424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  buf(_37198_[2], _25425_);
  buf(_25427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  buf(_37198_[3], _25428_);
  buf(_25429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  buf(_37198_[4], _25430_);
  buf(_25431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  buf(_37198_[5], _25432_);
  buf(_25433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  buf(_37198_[6], _25434_);
  buf(_25435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  buf(_37197_[0], _25436_);
  buf(_25437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  buf(_37197_[1], _25438_);
  buf(_25439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  buf(_37197_[2], _25440_);
  buf(_25441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  buf(_37197_[3], _25442_);
  buf(_25443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  buf(_37197_[4], _25444_);
  buf(_25445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  buf(_37197_[5], _25446_);
  buf(_25447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  buf(_37197_[6], _25448_);
  buf(_25449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  buf(_37196_[0], _25450_);
  buf(_25451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  buf(_37196_[1], _25452_);
  buf(_25453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  buf(_37196_[2], _25454_);
  buf(_25455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  buf(_37196_[3], _25456_);
  buf(_25457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  buf(_37196_[4], _25458_);
  buf(_25459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  buf(_37196_[5], _25460_);
  buf(_25461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  buf(_37196_[6], _25462_);
  buf(_25463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  buf(_37194_[0], _25464_);
  buf(_25465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  buf(_37194_[1], _25466_);
  buf(_25468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  buf(_37194_[2], _25469_);
  buf(_25470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  buf(_37194_[3], _25471_);
  buf(_25472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  buf(_37194_[4], _25473_);
  buf(_25474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  buf(_37194_[5], _25475_);
  buf(_25476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  buf(_37194_[6], _25477_);
  buf(_25478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  buf(_37193_[0], _25479_);
  buf(_25480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  buf(_37193_[1], _25481_);
  buf(_25482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  buf(_37193_[2], _25483_);
  buf(_25484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  buf(_37193_[3], _25485_);
  buf(_25486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  buf(_37193_[4], _25487_);
  buf(_25488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  buf(_37193_[5], _25489_);
  buf(_25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  buf(_37193_[6], _25491_);
  buf(_25492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  buf(_37192_[0], _25493_);
  buf(_25494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  buf(_37192_[1], _25495_);
  buf(_25496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  buf(_37192_[2], _25497_);
  buf(_25498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  buf(_37192_[3], _25499_);
  buf(_25500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  buf(_37192_[4], _25501_);
  buf(_25502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  buf(_37192_[5], _25503_);
  buf(_25504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  buf(_37192_[6], _25505_);
  buf(_25506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  buf(_37191_[0], _25507_);
  buf(_25509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  buf(_37191_[1], _25510_);
  buf(_25511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  buf(_37191_[2], _25512_);
  buf(_25513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  buf(_37191_[3], _25514_);
  buf(_25515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  buf(_37191_[4], _25516_);
  buf(_25517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  buf(_37191_[5], _25518_);
  buf(_25519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  buf(_37191_[6], _25520_);
  buf(_25521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  buf(_37190_[0], _25522_);
  buf(_25523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  buf(_37190_[1], _25524_);
  buf(_25525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  buf(_37190_[2], _25526_);
  buf(_25527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  buf(_37190_[3], _25528_);
  buf(_25529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  buf(_37190_[4], _25530_);
  buf(_25531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  buf(_37190_[5], _25532_);
  buf(_25533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  buf(_37190_[6], _25534_);
  buf(_25535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  buf(_37189_[0], _25536_);
  buf(_25537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  buf(_37189_[1], _25538_);
  buf(_25539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  buf(_37189_[2], _25540_);
  buf(_25541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  buf(_37189_[3], _25542_);
  buf(_25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  buf(_37189_[4], _25544_);
  buf(_25545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  buf(_37189_[5], _25546_);
  buf(_25547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  buf(_37189_[6], _25548_);
  buf(_25550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  buf(_37188_[0], _25551_);
  buf(_25552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  buf(_37188_[1], _25553_);
  buf(_25554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  buf(_37188_[2], _25555_);
  buf(_25556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  buf(_37188_[3], _25557_);
  buf(_25558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  buf(_37188_[4], _25559_);
  buf(_25560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  buf(_37188_[5], _25561_);
  buf(_25562_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  buf(_37188_[6], _25563_);
  buf(_25564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  buf(_37187_[0], _25565_);
  buf(_25566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  buf(_37187_[1], _25567_);
  buf(_25568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  buf(_37187_[2], _25569_);
  buf(_25570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  buf(_37187_[3], _25571_);
  buf(_25572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  buf(_37187_[4], _25573_);
  buf(_25574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  buf(_37187_[5], _25575_);
  buf(_25576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  buf(_37187_[6], _25577_);
  buf(_25578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  buf(_37186_[0], _25579_);
  buf(_25580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  buf(_37186_[1], _25581_);
  buf(_25582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  buf(_37186_[2], _25583_);
  buf(_25584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  buf(_37186_[3], _25585_);
  buf(_25586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  buf(_37186_[4], _25587_);
  buf(_25589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  buf(_37186_[5], _25591_);
  buf(_25594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  buf(_37186_[6], _25596_);
  buf(_25598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  buf(_37185_[0], _25600_);
  buf(_25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  buf(_37185_[1], _25604_);
  buf(_25606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  buf(_37185_[2], _25608_);
  buf(_25610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  buf(_37185_[3], _25612_);
  buf(_25614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  buf(_37185_[4], _25616_);
  buf(_25618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  buf(_37185_[5], _25620_);
  buf(_25622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  buf(_37185_[6], _25624_);
  buf(_25626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  buf(_37183_[0], _25628_);
  buf(_25630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  buf(_37183_[1], _25632_);
  buf(_25634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  buf(_37183_[2], _25636_);
  buf(_25638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  buf(_37183_[3], _25640_);
  buf(_25642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  buf(_37183_[4], _25644_);
  buf(_25646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  buf(_37183_[5], _25648_);
  buf(_25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  buf(_37183_[6], _25652_);
  buf(_25654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  buf(_37182_[0], _25656_);
  buf(_25658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  buf(_37182_[1], _25660_);
  buf(_25662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  buf(_37182_[2], _25664_);
  buf(_25666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  buf(_37182_[3], _25668_);
  buf(_25670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  buf(_37182_[4], _25672_);
  buf(_25675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  buf(_37182_[5], _25677_);
  buf(_25679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  buf(_37182_[6], _25681_);
  buf(_25683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  buf(_37181_[0], _25685_);
  buf(_25687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  buf(_37181_[1], _25689_);
  buf(_25691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  buf(_37181_[2], _25693_);
  buf(_25695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  buf(_37181_[3], _25697_);
  buf(_25699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  buf(_37181_[4], _25701_);
  buf(_25703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  buf(_37181_[5], _25705_);
  buf(_25707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  buf(_37181_[6], _25709_);
  buf(_25711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  buf(_37180_[0], _25713_);
  buf(_25715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  buf(_37180_[1], _25717_);
  buf(_25719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  buf(_37180_[2], _25721_);
  buf(_25723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  buf(_37180_[3], _25725_);
  buf(_25727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  buf(_37180_[4], _25729_);
  buf(_25731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  buf(_37180_[5], _25733_);
  buf(_25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  buf(_37180_[6], _25737_);
  buf(_25739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  buf(_37179_[0], _25741_);
  buf(_25743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  buf(_37179_[1], _25745_);
  buf(_25747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  buf(_37179_[2], _25749_);
  buf(_25751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  buf(_37179_[3], _25753_);
  buf(_25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  buf(_37179_[4], _25758_);
  buf(_25760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  buf(_37179_[5], _25762_);
  buf(_25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  buf(_37179_[6], _25766_);
  buf(_25768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  buf(_37178_[0], _25770_);
  buf(_25772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  buf(_37178_[1], _25774_);
  buf(_25776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  buf(_37178_[2], _25778_);
  buf(_25780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  buf(_37178_[3], _25782_);
  buf(_25784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  buf(_37178_[4], _25786_);
  buf(_25788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  buf(_37178_[5], _25790_);
  buf(_25792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  buf(_37178_[6], _25794_);
  buf(_25796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  buf(_37177_[0], _25798_);
  buf(_25800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  buf(_37177_[1], _25802_);
  buf(_25804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  buf(_37177_[2], _25806_);
  buf(_25808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  buf(_37177_[3], _25810_);
  buf(_25812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  buf(_37177_[4], _25814_);
  buf(_25816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  buf(_37177_[5], _25818_);
  buf(_25820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  buf(_37177_[6], _25822_);
  buf(_25824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  buf(_37176_[0], _25826_);
  buf(_25828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  buf(_37176_[1], _25830_);
  buf(_25832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  buf(_37176_[2], _25834_);
  buf(_25837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  buf(_37176_[3], _25839_);
  buf(_25841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  buf(_37176_[4], _25843_);
  buf(_25845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  buf(_37176_[5], _25847_);
  buf(_25849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  buf(_37176_[6], _25851_);
  buf(_25853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  buf(_37175_[0], _25855_);
  buf(_25857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  buf(_37175_[1], _25859_);
  buf(_25861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  buf(_37175_[2], _25863_);
  buf(_25865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  buf(_37175_[3], _25867_);
  buf(_25869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  buf(_37175_[4], _25871_);
  buf(_25873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  buf(_37175_[5], _25875_);
  buf(_25877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  buf(_37175_[6], _25879_);
  buf(_25881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  buf(_37174_[0], _25883_);
  buf(_25885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  buf(_37174_[1], _25887_);
  buf(_25889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  buf(_37174_[2], _25891_);
  buf(_25893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  buf(_37174_[3], _25895_);
  buf(_25897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  buf(_37174_[4], _25899_);
  buf(_25901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  buf(_37174_[5], _25903_);
  buf(_25905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  buf(_37174_[6], _25907_);
  buf(_25909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  buf(_37172_[0], _25911_);
  buf(_25913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  buf(_37172_[1], _25915_);
  buf(_25919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  buf(_37172_[2], _25921_);
  buf(_25923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  buf(_37172_[3], _25925_);
  buf(_25927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  buf(_37172_[4], _25929_);
  buf(_25931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  buf(_37172_[5], _25933_);
  buf(_25935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  buf(_37172_[6], _25937_);
  buf(_25939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  buf(_37171_[0], _25941_);
  buf(_25943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  buf(_37171_[1], _25945_);
  buf(_25947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  buf(_37171_[2], _25949_);
  buf(_25951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  buf(_37171_[3], _25953_);
  buf(_25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  buf(_37171_[4], _25957_);
  buf(_25959_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  buf(_37171_[5], _25961_);
  buf(_25963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  buf(_37171_[6], _25965_);
  buf(_25967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  buf(_37170_[0], _25969_);
  buf(_25971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  buf(_37170_[1], _25973_);
  buf(_25975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  buf(_37170_[2], _25977_);
  buf(_25979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  buf(_37170_[3], _25981_);
  buf(_25983_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  buf(_37170_[4], _25985_);
  buf(_25987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  buf(_37170_[5], _25989_);
  buf(_25991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  buf(_37170_[6], _25993_);
  buf(_25995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  buf(_37169_[0], _25997_);
  buf(_26000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  buf(_37169_[1], _26002_);
  buf(_26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  buf(_37169_[2], _26006_);
  buf(_26008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  buf(_37169_[3], _26010_);
  buf(_26012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  buf(_37169_[4], _26014_);
  buf(_26016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  buf(_37169_[5], _26018_);
  buf(_26020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  buf(_37169_[6], _26022_);
  buf(_26024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  buf(_37168_[0], _26026_);
  buf(_26028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  buf(_37168_[1], _26030_);
  buf(_26032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  buf(_37168_[2], _26034_);
  buf(_26036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  buf(_37168_[3], _26038_);
  buf(_26040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  buf(_37168_[4], _26042_);
  buf(_26044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  buf(_37168_[5], _26046_);
  buf(_26048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  buf(_37168_[6], _26050_);
  buf(_26052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  buf(_37167_[0], _26054_);
  buf(_26056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  buf(_37167_[1], _26058_);
  buf(_26060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  buf(_37167_[2], _26062_);
  buf(_26064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  buf(_37167_[3], _26066_);
  buf(_26068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  buf(_37167_[4], _26070_);
  buf(_26072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  buf(_37167_[5], _26074_);
  buf(_26076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  buf(_37167_[6], _26078_);
  buf(_26081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  buf(_37166_[0], _26083_);
  buf(_26085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  buf(_37166_[1], _26087_);
  buf(_26089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  buf(_37166_[2], _26091_);
  buf(_26093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  buf(_37166_[3], _26095_);
  buf(_26097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  buf(_37166_[4], _26099_);
  buf(_26101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  buf(_37166_[5], _26103_);
  buf(_26105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  buf(_37166_[6], _26107_);
  buf(_26109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  buf(_37165_[0], _26111_);
  buf(_26113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  buf(_37165_[1], _26115_);
  buf(_26117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  buf(_37165_[2], _26119_);
  buf(_26121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  buf(_37165_[3], _26123_);
  buf(_26125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  buf(_37165_[4], _26127_);
  buf(_26129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  buf(_37165_[5], _26131_);
  buf(_26133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  buf(_37165_[6], _26135_);
  buf(_26137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  buf(_37164_[0], _26139_);
  buf(_26141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  buf(_37164_[1], _26143_);
  buf(_26145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  buf(_37164_[2], _26147_);
  buf(_26149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  buf(_37164_[3], _26151_);
  buf(_26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  buf(_37164_[4], _26155_);
  buf(_26157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  buf(_37164_[5], _26159_);
  buf(_26162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  buf(_37164_[6], _26164_);
  buf(_26166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  buf(_37163_[0], _26168_);
  buf(_26170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  buf(_37163_[1], _26172_);
  buf(_26174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  buf(_37163_[2], _26176_);
  buf(_26178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  buf(_37163_[3], _26180_);
  buf(_26182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  buf(_37163_[4], _26184_);
  buf(_26186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  buf(_37163_[5], _26188_);
  buf(_26190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  buf(_37163_[6], _26192_);
  buf(_26194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  buf(_37329_[0], _26196_);
  buf(_26198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  buf(_37329_[1], _26200_);
  buf(_26202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  buf(_37329_[2], _26204_);
  buf(_26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  buf(_37329_[3], _26208_);
  buf(_26210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  buf(_37329_[4], _26212_);
  buf(_26214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  buf(_37329_[5], _26216_);
  buf(_26218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  buf(_37329_[6], _26220_);
  buf(_26222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  buf(_37328_[0], _26224_);
  buf(_26226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  buf(_37328_[1], _26228_);
  buf(_26230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  buf(_37328_[2], _26232_);
  buf(_26234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  buf(_37328_[3], _26236_);
  buf(_26238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  buf(_37328_[4], _26240_);
  buf(_26243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  buf(_37328_[5], _26245_);
  buf(_26247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  buf(_37328_[6], _26249_);
  buf(_26251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  buf(_37327_[0], _26253_);
  buf(_26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  buf(_37327_[1], _26257_);
  buf(_26259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  buf(_37327_[2], _26261_);
  buf(_26263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  buf(_37327_[3], _26265_);
  buf(_26267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  buf(_37327_[4], _26269_);
  buf(_26271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  buf(_37327_[5], _26273_);
  buf(_26275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  buf(_37327_[6], _26277_);
  buf(_26279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  buf(_37326_[0], _26281_);
  buf(_26283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  buf(_37326_[1], _26285_);
  buf(_26287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  buf(_37326_[2], _26289_);
  buf(_26291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  buf(_37326_[3], _26293_);
  buf(_26295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  buf(_37326_[4], _26297_);
  buf(_26299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  buf(_37326_[5], _26301_);
  buf(_26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  buf(_37326_[6], _26305_);
  buf(_26307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  buf(_37325_[0], _26309_);
  buf(_26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  buf(_37325_[1], _26313_);
  buf(_26315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  buf(_37325_[2], _26317_);
  buf(_26319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  buf(_37325_[3], _26321_);
  buf(_26324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  buf(_37325_[4], _26326_);
  buf(_26328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  buf(_37325_[5], _26330_);
  buf(_26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  buf(_37325_[6], _26334_);
  buf(_26336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  buf(_37324_[0], _26338_);
  buf(_26340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  buf(_37324_[1], _26342_);
  buf(_26344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  buf(_37324_[2], _26346_);
  buf(_26348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  buf(_37324_[3], _26350_);
  buf(_26352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  buf(_37324_[4], _26354_);
  buf(_26356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  buf(_37324_[5], _26358_);
  buf(_26360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  buf(_37324_[6], _26362_);
  buf(_26364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  buf(_37323_[0], _26366_);
  buf(_26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  buf(_37323_[1], _26370_);
  buf(_26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  buf(_37323_[2], _26374_);
  buf(_26376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  buf(_37323_[3], _26378_);
  buf(_26380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  buf(_37323_[4], _26382_);
  buf(_26384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  buf(_37323_[5], _26386_);
  buf(_26388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  buf(_37323_[6], _26390_);
  buf(_26392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  buf(_37322_[0], _26394_);
  buf(_26396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  buf(_37322_[1], _26398_);
  buf(_26400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  buf(_37322_[2], _26402_);
  buf(_26405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  buf(_37322_[3], _26407_);
  buf(_26409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  buf(_37322_[4], _26411_);
  buf(_26413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  buf(_37322_[5], _26415_);
  buf(_26417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  buf(_37322_[6], _26419_);
  buf(_26421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  buf(_37321_[0], _26423_);
  buf(_26425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  buf(_37321_[1], _26427_);
  buf(_26429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  buf(_37321_[2], _26431_);
  buf(_26433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  buf(_37321_[3], _26435_);
  buf(_26437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  buf(_37321_[4], _26439_);
  buf(_26441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  buf(_37321_[5], _26443_);
  buf(_26445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  buf(_37321_[6], _26447_);
  buf(_26449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  buf(_37320_[0], _26451_);
  buf(_26453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  buf(_37320_[1], _26455_);
  buf(_26457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  buf(_37320_[2], _26459_);
  buf(_26461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  buf(_37320_[3], _26463_);
  buf(_26465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  buf(_37320_[4], _26467_);
  buf(_26469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  buf(_37320_[5], _26471_);
  buf(_26473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  buf(_37320_[6], _26475_);
  buf(_26477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  buf(_37319_[0], _26479_);
  buf(_26481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  buf(_37319_[1], _26483_);
  buf(_26486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  buf(_37319_[2], _26488_);
  buf(_26490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  buf(_37319_[3], _26492_);
  buf(_26494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  buf(_37319_[4], _26496_);
  buf(_26498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  buf(_37319_[5], _26500_);
  buf(_26502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  buf(_37319_[6], _26504_);
  buf(_26506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  buf(_37318_[0], _26508_);
  buf(_26510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  buf(_37318_[1], _26512_);
  buf(_26514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  buf(_37318_[2], _26516_);
  buf(_26518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  buf(_37318_[3], _26520_);
  buf(_26522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  buf(_37318_[4], _26524_);
  buf(_26526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  buf(_37318_[5], _26528_);
  buf(_26530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  buf(_37318_[6], _26532_);
  buf(_26534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  buf(_37317_[0], _26536_);
  buf(_26538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  buf(_37317_[1], _26540_);
  buf(_26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  buf(_37317_[2], _26544_);
  buf(_26546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  buf(_37317_[3], _26548_);
  buf(_26550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  buf(_37317_[4], _26552_);
  buf(_26554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  buf(_37317_[5], _26556_);
  buf(_26558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  buf(_37317_[6], _26560_);
  buf(_26562_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  buf(_37316_[0], _26564_);
  buf(_26567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  buf(_37316_[1], _26569_);
  buf(_26571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  buf(_37316_[2], _26573_);
  buf(_26575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  buf(_37316_[3], _26577_);
  buf(_26579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  buf(_37316_[4], _26581_);
  buf(_26583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  buf(_37316_[5], _26585_);
  buf(_26587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  buf(_37316_[6], _26589_);
  buf(_26591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  buf(_37315_[0], _26593_);
  buf(_26595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  buf(_37315_[1], _26597_);
  buf(_26599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  buf(_37315_[2], _26601_);
  buf(_26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  buf(_37315_[3], _26605_);
  buf(_26607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  buf(_37315_[4], _26609_);
  buf(_26611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  buf(_37315_[5], _26613_);
  buf(_26615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  buf(_37315_[6], _26617_);
  buf(_26619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  buf(_37314_[0], _26621_);
  buf(_26623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  buf(_37314_[1], _26625_);
  buf(_26627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  buf(_37314_[2], _26629_);
  buf(_26631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  buf(_37314_[3], _26633_);
  buf(_26635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  buf(_37314_[4], _26637_);
  buf(_26639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  buf(_37314_[5], _26641_);
  buf(_26643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  buf(_37314_[6], _26645_);
  buf(_26648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  buf(_37313_[0], _26650_);
  buf(_26652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  buf(_37313_[1], _26654_);
  buf(_26656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  buf(_37313_[2], _26658_);
  buf(_26660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  buf(_37313_[3], _26662_);
  buf(_26664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  buf(_37313_[4], _26666_);
  buf(_26668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  buf(_37313_[5], _26670_);
  buf(_26672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  buf(_37313_[6], _26674_);
  buf(_26676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  buf(_37312_[0], _26678_);
  buf(_26680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  buf(_37312_[1], _26682_);
  buf(_26684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  buf(_37312_[2], _26686_);
  buf(_26688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  buf(_37312_[3], _26690_);
  buf(_26692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  buf(_37312_[4], _26694_);
  buf(_26696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  buf(_37312_[5], _26698_);
  buf(_26700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  buf(_37312_[6], _26702_);
  buf(_26704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  buf(_37311_[0], _26706_);
  buf(_26708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  buf(_37311_[1], _26710_);
  buf(_26712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  buf(_37311_[2], _26714_);
  buf(_26716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  buf(_37311_[3], _26718_);
  buf(_26720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  buf(_37311_[4], _26722_);
  buf(_26724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  buf(_37311_[5], _26726_);
  buf(_26730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  buf(_37311_[6], _26732_);
  buf(_26734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  buf(_37310_[0], _26736_);
  buf(_26738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  buf(_37310_[1], _26740_);
  buf(_26742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  buf(_37310_[2], _26744_);
  buf(_26746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  buf(_37310_[3], _26748_);
  buf(_26750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  buf(_37310_[4], _26752_);
  buf(_26754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  buf(_37310_[5], _26756_);
  buf(_26758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  buf(_37310_[6], _26760_);
  buf(_26762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  buf(_37309_[0], _26764_);
  buf(_26766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  buf(_37309_[1], _26768_);
  buf(_26770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  buf(_37309_[2], _26772_);
  buf(_26774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  buf(_37309_[3], _26776_);
  buf(_26778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  buf(_37309_[4], _26780_);
  buf(_26782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  buf(_37309_[5], _26784_);
  buf(_26786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  buf(_37309_[6], _26788_);
  buf(_26790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  buf(_37308_[0], _26792_);
  buf(_26794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  buf(_37308_[1], _26796_);
  buf(_26798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  buf(_37308_[2], _26800_);
  buf(_26802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  buf(_37308_[3], _26804_);
  buf(_26806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  buf(_37308_[4], _26808_);
  buf(_26811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  buf(_37308_[5], _26813_);
  buf(_26815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  buf(_37308_[6], _26817_);
  buf(_26819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  buf(_37307_[0], _26821_);
  buf(_26823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  buf(_37307_[1], _26825_);
  buf(_26827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  buf(_37307_[2], _26829_);
  buf(_26831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  buf(_37307_[3], _26833_);
  buf(_26835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  buf(_37307_[4], _26837_);
  buf(_26839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  buf(_37307_[5], _26841_);
  buf(_26843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  buf(_37307_[6], _26845_);
  buf(_26847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  buf(_37306_[0], _26849_);
  buf(_26851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  buf(_37306_[1], _26853_);
  buf(_26855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  buf(_37306_[2], _26857_);
  buf(_26859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  buf(_37306_[3], _26861_);
  buf(_26863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  buf(_37306_[4], _26865_);
  buf(_26867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  buf(_37306_[5], _26869_);
  buf(_26871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  buf(_37306_[6], _26873_);
  buf(_26875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  buf(_37305_[0], _26877_);
  buf(_26879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  buf(_37305_[1], _26881_);
  buf(_26883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  buf(_37305_[2], _26885_);
  buf(_26887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  buf(_37305_[3], _26889_);
  buf(_26892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  buf(_37305_[4], _26894_);
  buf(_26896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  buf(_37305_[5], _26898_);
  buf(_26900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  buf(_37305_[6], _26902_);
  buf(_26904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  buf(_37416_[0], _26906_);
  buf(_26908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  buf(_37416_[1], _26910_);
  buf(_26912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  buf(_37416_[2], _26914_);
  buf(_26916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  buf(_37416_[3], _26918_);
  buf(_26920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  buf(_37416_[4], _26922_);
  buf(_26924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  buf(_37416_[5], _26926_);
  buf(_26928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  buf(_37416_[6], _26930_);
  buf(_26932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  buf(_37415_[0], _26934_);
  buf(_26936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  buf(_37415_[1], _26938_);
  buf(_26940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  buf(_37415_[2], _26942_);
  buf(_26944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  buf(_37415_[3], _26946_);
  buf(_26948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  buf(_37415_[4], _26950_);
  buf(_26952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  buf(_37415_[5], _26954_);
  buf(_26956_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  buf(_37415_[6], _26958_);
  buf(_26960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  buf(_37414_[0], _26962_);
  buf(_26964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  buf(_37414_[1], _26966_);
  buf(_26968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  buf(_37414_[2], _26970_);
  buf(_26973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  buf(_37414_[3], _26975_);
  buf(_26977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  buf(_37414_[4], _26979_);
  buf(_26981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  buf(_37414_[5], _26983_);
  buf(_26985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  buf(_37414_[6], _26987_);
  buf(_26989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  buf(_37304_[0], _26991_);
  buf(_26993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  buf(_37304_[1], _26995_);
  buf(_26997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  buf(_37304_[2], _26999_);
  buf(_27001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  buf(_37304_[3], _27003_);
  buf(_27005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  buf(_37304_[4], _27007_);
  buf(_27009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  buf(_37304_[5], _27011_);
  buf(_27013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  buf(_37304_[6], _27015_);
  buf(_27017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  buf(_37303_[0], _27019_);
  buf(_27021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  buf(_37303_[1], _27023_);
  buf(_27025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  buf(_37303_[2], _27027_);
  buf(_27029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  buf(_37303_[3], _27031_);
  buf(_27033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  buf(_37303_[4], _27035_);
  buf(_27037_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  buf(_37303_[5], _27039_);
  buf(_27041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  buf(_37303_[6], _27043_);
  buf(_27045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  buf(_37412_[0], _27047_);
  buf(_27049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  buf(_37412_[1], _27051_);
  buf(_27054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  buf(_37412_[2], _27056_);
  buf(_27058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  buf(_37412_[3], _27060_);
  buf(_27062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  buf(_37412_[4], _27064_);
  buf(_27066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  buf(_37412_[5], _27068_);
  buf(_27070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  buf(_37412_[6], _27072_);
  buf(_27074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  buf(_37411_[0], _27076_);
  buf(_27078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  buf(_37411_[1], _27080_);
  buf(_27082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  buf(_37411_[2], _27084_);
  buf(_27086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  buf(_37411_[3], _27088_);
  buf(_27090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  buf(_37411_[4], _27092_);
  buf(_27094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  buf(_37411_[5], _27096_);
  buf(_27098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  buf(_37411_[6], _27100_);
  buf(_27102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  buf(_37410_[0], _27104_);
  buf(_27106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  buf(_37410_[1], _27108_);
  buf(_27110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  buf(_37410_[2], _27112_);
  buf(_27114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  buf(_37410_[3], _27116_);
  buf(_27118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  buf(_37410_[4], _27120_);
  buf(_27122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  buf(_37410_[5], _27124_);
  buf(_27126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  buf(_37410_[6], _27128_);
  buf(_27130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  buf(_37409_[0], _27132_);
  buf(_27135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  buf(_37409_[1], _27137_);
  buf(_27139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  buf(_37409_[2], _27141_);
  buf(_27143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  buf(_37409_[3], _27145_);
  buf(_27147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  buf(_37409_[4], _27149_);
  buf(_27151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  buf(_37409_[5], _27153_);
  buf(_27155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  buf(_37409_[6], _27157_);
  buf(_27159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  buf(_37408_[0], _27161_);
  buf(_27163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  buf(_37408_[1], _27165_);
  buf(_27167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  buf(_37408_[2], _27169_);
  buf(_27171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  buf(_37408_[3], _27173_);
  buf(_27175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  buf(_37408_[4], _27177_);
  buf(_27179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  buf(_37408_[5], _27181_);
  buf(_27183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  buf(_37408_[6], _27185_);
  buf(_27187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  buf(_37407_[0], _27189_);
  buf(_27191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  buf(_37407_[1], _27193_);
  buf(_27195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  buf(_37407_[2], _27197_);
  buf(_27199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  buf(_37407_[3], _27201_);
  buf(_27203_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  buf(_37407_[4], _27205_);
  buf(_27207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  buf(_37407_[5], _27209_);
  buf(_27211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  buf(_37407_[6], _27213_);
  buf(_27216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  buf(_37406_[0], _27218_);
  buf(_27220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  buf(_37406_[1], _27222_);
  buf(_27224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  buf(_37406_[2], _27226_);
  buf(_27228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  buf(_37406_[3], _27230_);
  buf(_27232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  buf(_37406_[4], _27234_);
  buf(_27236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  buf(_37406_[5], _27238_);
  buf(_27240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  buf(_37406_[6], _27242_);
  buf(_27244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  buf(_37405_[0], _27246_);
  buf(_27248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  buf(_37405_[1], _27250_);
  buf(_27252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  buf(_37405_[2], _27254_);
  buf(_27256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  buf(_37405_[3], _27258_);
  buf(_27260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  buf(_37405_[4], _27262_);
  buf(_27264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  buf(_37405_[5], _27266_);
  buf(_27268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  buf(_37405_[6], _27270_);
  buf(_27272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  buf(_37404_[0], _27274_);
  buf(_27276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  buf(_37404_[1], _27278_);
  buf(_27280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  buf(_37404_[2], _27282_);
  buf(_27284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  buf(_37404_[3], _27286_);
  buf(_27288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  buf(_37404_[4], _27290_);
  buf(_27292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  buf(_37404_[5], _27294_);
  buf(_27297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  buf(_37404_[6], _27299_);
  buf(_27301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  buf(_37403_[0], _27303_);
  buf(_27305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  buf(_37403_[1], _27307_);
  buf(_27309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  buf(_37403_[2], _27311_);
  buf(_27313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  buf(_37403_[3], _27315_);
  buf(_27317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  buf(_37403_[4], _27319_);
  buf(_27321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  buf(_37403_[5], _27323_);
  buf(_27325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  buf(_37403_[6], _27327_);
  buf(_27329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  buf(_37401_[0], _27331_);
  buf(_27333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  buf(_37401_[1], _27335_);
  buf(_27337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  buf(_37401_[2], _27339_);
  buf(_27341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  buf(_37401_[3], _27343_);
  buf(_27345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  buf(_37401_[4], _27347_);
  buf(_27349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  buf(_37401_[5], _27351_);
  buf(_27353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  buf(_37401_[6], _27355_);
  buf(_27357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  buf(_37400_[0], _27359_);
  buf(_27361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  buf(_37400_[1], _27363_);
  buf(_27365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  buf(_37400_[2], _27367_);
  buf(_27369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  buf(_37400_[3], _27371_);
  buf(_27373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  buf(_37400_[4], _27375_);
  buf(_27378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  buf(_37400_[5], _27380_);
  buf(_27382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  buf(_37400_[6], _27384_);
  buf(_27386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  buf(_37399_[0], _27388_);
  buf(_27390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  buf(_37399_[1], _27392_);
  buf(_27394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  buf(_37399_[2], _27396_);
  buf(_27398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  buf(_37399_[3], _27400_);
  buf(_27402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  buf(_37399_[4], _27404_);
  buf(_27406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  buf(_37399_[5], _27408_);
  buf(_27410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  buf(_37399_[6], _27412_);
  buf(_27414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  buf(_37398_[0], _27416_);
  buf(_27418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  buf(_37398_[1], _27420_);
  buf(_27422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  buf(_37398_[2], _27424_);
  buf(_27426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  buf(_37398_[3], _27428_);
  buf(_27430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  buf(_37398_[4], _27432_);
  buf(_27434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  buf(_37398_[5], _27436_);
  buf(_27438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  buf(_37398_[6], _27440_);
  buf(_27442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  buf(_37397_[0], _27444_);
  buf(_27446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  buf(_37397_[1], _27448_);
  buf(_27450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  buf(_37397_[2], _27452_);
  buf(_27454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  buf(_37397_[3], _27456_);
  buf(_27459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  buf(_37397_[4], _27461_);
  buf(_27463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  buf(_37397_[5], _27465_);
  buf(_27467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  buf(_37397_[6], _27469_);
  buf(_27471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  buf(_37396_[0], _27473_);
  buf(_27475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  buf(_37396_[1], _27477_);
  buf(_27479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  buf(_37396_[2], _27481_);
  buf(_27483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  buf(_37396_[3], _27485_);
  buf(_27487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  buf(_37396_[4], _27489_);
  buf(_27491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  buf(_37396_[5], _27493_);
  buf(_27495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  buf(_37396_[6], _27497_);
  buf(_27499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  buf(_37392_[0], _27501_);
  buf(_27503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  buf(_37392_[1], _27505_);
  buf(_27507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  buf(_37392_[2], _27509_);
  buf(_27511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  buf(_37392_[3], _27513_);
  buf(_27515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  buf(_37392_[4], _27517_);
  buf(_27519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  buf(_37392_[5], _27521_);
  buf(_27523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  buf(_37392_[6], _27525_);
  buf(_27527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  buf(_37390_[0], _27529_);
  buf(_27531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  buf(_37390_[1], _27533_);
  buf(_27535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  buf(_37390_[2], _27537_);
  buf(_27541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  buf(_37390_[3], _27543_);
  buf(_27545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  buf(_37390_[4], _27547_);
  buf(_27549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  buf(_37390_[5], _27551_);
  buf(_27553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  buf(_37390_[6], _27555_);
  buf(_27557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  buf(_37389_[0], _27559_);
  buf(_27561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  buf(_37389_[1], _27563_);
  buf(_27565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  buf(_37389_[2], _27567_);
  buf(_27569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  buf(_37389_[3], _27571_);
  buf(_27573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  buf(_37389_[4], _27575_);
  buf(_27577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  buf(_37389_[5], _27579_);
  buf(_27581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  buf(_37389_[6], _27583_);
  buf(_27585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  buf(_37388_[0], _27587_);
  buf(_27589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  buf(_37388_[1], _27591_);
  buf(_27593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  buf(_37388_[2], _27595_);
  buf(_27597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  buf(_37388_[3], _27599_);
  buf(_27601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  buf(_37388_[4], _27603_);
  buf(_27605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  buf(_37388_[5], _27607_);
  buf(_27609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  buf(_37388_[6], _27611_);
  buf(_27613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  buf(_37387_[0], _27615_);
  buf(_27617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  buf(_37387_[1], _27619_);
  buf(_27622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  buf(_37387_[2], _27624_);
  buf(_27626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  buf(_37387_[3], _27628_);
  buf(_27630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  buf(_37387_[4], _27632_);
  buf(_27634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  buf(_37387_[5], _27636_);
  buf(_27638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  buf(_37387_[6], _27640_);
  buf(_27642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  buf(_37386_[0], _27644_);
  buf(_27646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  buf(_37386_[1], _27648_);
  buf(_27650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  buf(_37386_[2], _27652_);
  buf(_27654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  buf(_37386_[3], _27656_);
  buf(_27658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  buf(_37386_[4], _27660_);
  buf(_27662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  buf(_37386_[5], _27664_);
  buf(_27666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  buf(_37386_[6], _27668_);
  buf(_27670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  buf(_37384_[0], _27672_);
  buf(_27674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  buf(_37384_[1], _27676_);
  buf(_27678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  buf(_37384_[2], _27680_);
  buf(_27682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  buf(_37384_[3], _27684_);
  buf(_27686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  buf(_37384_[4], _27688_);
  buf(_27690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  buf(_37384_[5], _27692_);
  buf(_27694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  buf(_37384_[6], _27696_);
  buf(_27698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  buf(_37383_[0], _27700_);
  buf(_27703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  buf(_37383_[1], _27705_);
  buf(_27707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  buf(_37383_[2], _27709_);
  buf(_27711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  buf(_37383_[3], _27713_);
  buf(_27715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  buf(_37383_[4], _27717_);
  buf(_27719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  buf(_37383_[5], _27721_);
  buf(_27723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  buf(_37383_[6], _27725_);
  buf(_27727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  buf(_37382_[0], _27729_);
  buf(_27731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  buf(_37382_[1], _27733_);
  buf(_27735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  buf(_37382_[2], _27737_);
  buf(_27739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  buf(_37382_[3], _27741_);
  buf(_27743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  buf(_37382_[4], _27745_);
  buf(_27747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  buf(_37382_[5], _27749_);
  buf(_27751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  buf(_37382_[6], _27753_);
  buf(_27755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  buf(_37381_[0], _27757_);
  buf(_27759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  buf(_37381_[1], _27761_);
  buf(_27763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  buf(_37381_[2], _27765_);
  buf(_27767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  buf(_37381_[3], _27769_);
  buf(_27771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  buf(_37381_[4], _27773_);
  buf(_27775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  buf(_37381_[5], _27777_);
  buf(_27779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  buf(_37381_[6], _27781_);
  buf(_27784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  buf(_37379_[0], _27786_);
  buf(_27788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  buf(_37379_[1], _27790_);
  buf(_27792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  buf(_37379_[2], _27794_);
  buf(_27796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  buf(_37379_[3], _27798_);
  buf(_27800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  buf(_37379_[4], _27802_);
  buf(_27804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  buf(_37379_[5], _27806_);
  buf(_27808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  buf(_37379_[6], _27810_);
  buf(_27812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  buf(_37378_[0], _27814_);
  buf(_27816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  buf(_37378_[1], _27818_);
  buf(_27820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  buf(_37378_[2], _27822_);
  buf(_27824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  buf(_37378_[3], _27826_);
  buf(_27828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  buf(_37378_[4], _27830_);
  buf(_27832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  buf(_37378_[5], _27834_);
  buf(_27836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  buf(_37378_[6], _27838_);
  buf(_27840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  buf(_37377_[0], _27842_);
  buf(_27844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  buf(_37377_[1], _27846_);
  buf(_27848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  buf(_37377_[2], _27850_);
  buf(_27852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  buf(_37377_[3], _27854_);
  buf(_27856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  buf(_37377_[4], _27858_);
  buf(_27860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  buf(_37377_[5], _27862_);
  buf(_27865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  buf(_37377_[6], _27867_);
  buf(_27869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  buf(_37376_[0], _27871_);
  buf(_27873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  buf(_37376_[1], _27875_);
  buf(_27877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  buf(_37376_[2], _27879_);
  buf(_27881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  buf(_37376_[3], _27883_);
  buf(_27885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  buf(_37376_[4], _27887_);
  buf(_27889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  buf(_37376_[5], _27891_);
  buf(_27893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  buf(_37376_[6], _27895_);
  buf(_27897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  buf(_37374_[0], _27899_);
  buf(_27901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  buf(_37374_[1], _27903_);
  buf(_27905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  buf(_37374_[2], _27907_);
  buf(_27909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  buf(_37374_[3], _27911_);
  buf(_27913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  buf(_37374_[4], _27915_);
  buf(_27917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  buf(_37374_[5], _27919_);
  buf(_27921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  buf(_37374_[6], _27923_);
  buf(_27925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  buf(_37372_[0], _27927_);
  buf(_27929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  buf(_37372_[1], _27931_);
  buf(_27933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  buf(_37372_[2], _27935_);
  buf(_27937_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  buf(_37372_[3], _27939_);
  buf(_27941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  buf(_37372_[4], _27943_);
  buf(_27946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  buf(_37372_[5], _27948_);
  buf(_27950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  buf(_37372_[6], _27952_);
  buf(_27954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  buf(_37370_[0], _27956_);
  buf(_27958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  buf(_37370_[1], _27960_);
  buf(_27962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  buf(_37370_[2], _27964_);
  buf(_27966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  buf(_37370_[3], _27968_);
  buf(_27970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  buf(_37370_[4], _27972_);
  buf(_27974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  buf(_37370_[5], _27976_);
  buf(_27978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  buf(_37370_[6], _27980_);
  buf(_27982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  buf(_37368_[0], _27984_);
  buf(_27986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  buf(_37368_[1], _27988_);
  buf(_27990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  buf(_37368_[2], _27992_);
  buf(_27994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  buf(_37368_[3], _27996_);
  buf(_27998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  buf(_37368_[4], _28000_);
  buf(_28002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  buf(_37368_[5], _28004_);
  buf(_28006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  buf(_37368_[6], _28008_);
  buf(_28010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  buf(_37367_[0], _28012_);
  buf(_28014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  buf(_37367_[1], _28016_);
  buf(_28018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  buf(_37367_[2], _28020_);
  buf(_28022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  buf(_37367_[3], _28024_);
  buf(_28027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  buf(_37367_[4], _28029_);
  buf(_28031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  buf(_37367_[5], _28033_);
  buf(_28035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  buf(_37367_[6], _28037_);
  buf(_28039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  buf(_37366_[0], _28041_);
  buf(_28043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  buf(_37366_[1], _28045_);
  buf(_28047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  buf(_37366_[2], _28049_);
  buf(_28051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  buf(_37366_[3], _28053_);
  buf(_28055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  buf(_37366_[4], _28057_);
  buf(_28059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  buf(_37366_[5], _28061_);
  buf(_28063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  buf(_37366_[6], _28065_);
  buf(_28067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  buf(_37173_[0], _28069_);
  buf(_28071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  buf(_37173_[1], _28073_);
  buf(_28075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  buf(_37173_[2], _28077_);
  buf(_28079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  buf(_37173_[3], _28081_);
  buf(_28083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  buf(_37173_[4], _28085_);
  buf(_28087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  buf(_37173_[5], _28089_);
  buf(_28091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  buf(_37173_[6], _28093_);
  buf(_28095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  buf(_37330_[0], _28097_);
  buf(_28099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  buf(_37330_[1], _28101_);
  buf(_28103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  buf(_37330_[2], _28105_);
  buf(_28108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  buf(_37330_[3], _28110_);
  buf(_28112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  buf(_37330_[4], _28114_);
  buf(_28116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  buf(_37330_[5], _28118_);
  buf(_28120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  buf(_37330_[6], _28122_);
  buf(_28124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  buf(_37418_[0], _28126_);
  buf(_28128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  buf(_37418_[1], _28130_);
  buf(_28132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  buf(_37418_[2], _28134_);
  buf(_28136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  buf(_37418_[3], _28138_);
  buf(_28140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  buf(_37418_[4], _28142_);
  buf(_28144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  buf(_37418_[5], _28146_);
  buf(_28148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  buf(_37418_[6], _28150_);
  buf(_28152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  buf(_37417_[0], _28154_);
  buf(_28156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  buf(_37417_[1], _28158_);
  buf(_28160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  buf(_37417_[2], _28162_);
  buf(_28164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  buf(_37417_[3], _28166_);
  buf(_28168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  buf(_37417_[4], _28170_);
  buf(_28172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  buf(_37417_[5], _28174_);
  buf(_28176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  buf(_37417_[6], _28178_);
  buf(_28180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  buf(_37413_[0], _28182_);
  buf(_28184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  buf(_37413_[1], _28186_);
  buf(_28189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  buf(_37413_[2], _28191_);
  buf(_28193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  buf(_37413_[3], _28195_);
  buf(_28197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  buf(_37413_[4], _28199_);
  buf(_28201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  buf(_37413_[5], _28203_);
  buf(_28205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  buf(_37413_[6], _28207_);
  buf(_28209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  buf(_37362_[0], _28211_);
  buf(_28213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  buf(_37362_[1], _28215_);
  buf(_28217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  buf(_37362_[2], _28219_);
  buf(_28221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  buf(_37362_[3], _28223_);
  buf(_28225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  buf(_37362_[4], _28227_);
  buf(_28229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  buf(_37362_[5], _28231_);
  buf(_28233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  buf(_37362_[6], _28235_);
  buf(_28237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  buf(_37402_[0], _28239_);
  buf(_28241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  buf(_37402_[1], _28243_);
  buf(_28245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  buf(_37402_[2], _28247_);
  buf(_28249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  buf(_37402_[3], _28251_);
  buf(_28253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  buf(_37402_[4], _28255_);
  buf(_28257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  buf(_37402_[5], _28259_);
  buf(_28261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  buf(_37402_[6], _28263_);
  buf(_28265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  buf(_37391_[0], _28267_);
  buf(_28270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  buf(_37391_[1], _28272_);
  buf(_28274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  buf(_37391_[2], _28276_);
  buf(_28278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  buf(_37391_[3], _28280_);
  buf(_28282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  buf(_37391_[4], _28284_);
  buf(_28286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  buf(_37391_[5], _28288_);
  buf(_28290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  buf(_37391_[6], _28292_);
  buf(_28294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  buf(_37380_[0], _28296_);
  buf(_28298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  buf(_37380_[1], _28300_);
  buf(_28302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  buf(_37380_[2], _28304_);
  buf(_28306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  buf(_37380_[3], _28308_);
  buf(_28310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  buf(_37380_[4], _28312_);
  buf(_28314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  buf(_37380_[5], _28316_);
  buf(_28318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  buf(_37380_[6], _28320_);
  buf(_28322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  buf(_37363_[0], _28324_);
  buf(_28326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  buf(_37363_[1], _28328_);
  buf(_28330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  buf(_37363_[2], _28332_);
  buf(_28334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  buf(_37363_[3], _28336_);
  buf(_28338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  buf(_37363_[4], _28340_);
  buf(_28342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  buf(_37363_[5], _28344_);
  buf(_28346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  buf(_37363_[6], _28348_);
  buf(_28352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  buf(_37369_[0], _28354_);
  buf(_28356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  buf(_37369_[1], _28358_);
  buf(_28360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  buf(_37369_[2], _28362_);
  buf(_28364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  buf(_37369_[3], _28366_);
  buf(_28368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  buf(_37369_[4], _28370_);
  buf(_28372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  buf(_37369_[5], _28374_);
  buf(_28376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  buf(_37369_[6], _28378_);
  buf(_28380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  buf(_37358_[0], _28382_);
  buf(_28384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  buf(_37358_[1], _28386_);
  buf(_28388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  buf(_37358_[2], _28390_);
  buf(_28392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  buf(_37358_[3], _28394_);
  buf(_28396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  buf(_37358_[4], _28398_);
  buf(_28400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  buf(_37358_[5], _28402_);
  buf(_28404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  buf(_37358_[6], _28406_);
  buf(_28408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  buf(_37331_[0], _28410_);
  buf(_28412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  buf(_37331_[1], _28414_);
  buf(_28416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  buf(_37331_[2], _28418_);
  buf(_28420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  buf(_37331_[3], _28422_);
  buf(_28424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  buf(_37331_[4], _28426_);
  buf(_28428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  buf(_37331_[5], _28430_);
  buf(_28433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  buf(_37331_[6], _28435_);
  buf(_28437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  buf(_37361_[5], _28439_);
  buf(_28441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  buf(_37361_[4], _28443_);
  buf(_28445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  buf(_37361_[3], _28447_);
  buf(_28449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  buf(_37361_[6], _28451_);
  buf(_28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  buf(_37361_[2], _28455_);
  buf(_28457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  buf(_37361_[1], _28459_);
  buf(_29296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  buf(_30277_, p1_in[7]);
  buf(_30279_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(_30283_, p2_in[7]);
  buf(_30285_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(_30288_, p3_in[7]);
  buf(_30290_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(_30297_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(_30301_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(_30308_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(_30313_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(_30321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(_30325_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(_30331_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(_30339_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(_30346_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(_30358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(_30374_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(_30379_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(_30392_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(_30396_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(_30402_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(_30409_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(_30424_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(_30428_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(_30440_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(_30451_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(_30456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(_30459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(_30466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(_30471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(_30478_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(_30483_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(_30490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(_30497_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(_30512_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(_30517_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(_30531_, p0_in[0]);
  buf(_30534_, p0_in[1]);
  buf(_30537_, p0_in[2]);
  buf(_30540_, p0_in[3]);
  buf(_30543_, p0_in[4]);
  buf(_30546_, p0_in[5]);
  buf(_30549_, p0_in[6]);
  buf(_30552_, p1_in[0]);
  buf(_30555_, p1_in[1]);
  buf(_30558_, p1_in[2]);
  buf(_30561_, p1_in[3]);
  buf(_30564_, p1_in[4]);
  buf(_30567_, p1_in[5]);
  buf(_30570_, p1_in[6]);
  buf(_30573_, p2_in[0]);
  buf(_30576_, p2_in[1]);
  buf(_30579_, p2_in[2]);
  buf(_30582_, p2_in[3]);
  buf(_30585_, p2_in[4]);
  buf(_30588_, p2_in[5]);
  buf(_30591_, p2_in[6]);
  buf(_30594_, p3_in[0]);
  buf(_30597_, p3_in[1]);
  buf(_30601_, p3_in[2]);
  buf(_30604_, p3_in[3]);
  buf(_30607_, p3_in[4]);
  buf(_30610_, p3_in[5]);
  buf(_30613_, p3_in[6]);
  buf(_30655_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(_30666_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(_30670_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(_30677_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(_30685_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(_30689_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(_30691_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(_30702_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(_30705_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(_30736_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(_30743_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(_30761_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(_30765_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(_30769_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(_30773_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(_30777_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(_30780_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(_30783_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(_30794_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(_30797_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(_30800_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(_30803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(_30806_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(_30809_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(_30812_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(_30822_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  buf(_30855_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  buf(_30857_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  buf(_30868_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  buf(_30870_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  buf(_30873_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  buf(_30875_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  buf(_30878_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  buf(_30951_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  buf(_30961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(_30964_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(_30971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  buf(_30975_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(_30978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(_30981_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(_30984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(_30990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  buf(_30995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  buf(_30997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  buf(_30999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(_31018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(_31022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(_31029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(_31031_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(_31037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(_31064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(_31066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(_31078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(_31082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(_31135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(_31144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(_31150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(_31158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(_31176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(_31178_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(_31202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(_31204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(_31208_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(_31210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(_31216_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(_31232_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(_31243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(_31246_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(_31251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(_31254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(_31268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(_31271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(_31275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(_31277_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(_31285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(_31290_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(_00018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(_00022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(_00155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(_00158_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(_00162_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(_00201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  buf(_00204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(_00207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(_00224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(_00230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(_00236_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(_00246_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(_00250_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(_00256_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(_00264_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  buf(_00270_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(_00277_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  buf(_00289_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(_00291_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff );
  buf(_00315_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(_00318_, \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(_00327_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(_00340_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  buf(_00343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(_00345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  buf(_00347_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  buf(_00350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(_00374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  buf(_00382_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(_00390_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(_00402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(_00408_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  buf(_00417_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  buf(_00435_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(_00453_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(_00464_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(_00473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  buf(_00495_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(_00508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(_00512_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(_00517_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(_00546_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(_00549_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(_00551_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(_00554_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(_00556_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(_00559_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(_00561_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(_00565_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  buf(_00627_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  buf(_00641_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  buf(_00762_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(_00765_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  buf(_00776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  buf(_00784_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(_00791_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  buf(_00801_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(_00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  buf(_00806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  buf(_00810_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  buf(_00813_, rxd_i);
  buf(_00814_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  buf(_00818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(_00824_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  buf(_00831_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  buf(_00834_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(_00839_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(_00841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(_00847_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  buf(_00848_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  buf(_00859_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  buf(_00869_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  buf(_00877_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  buf(_00878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(_00888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(_00894_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  buf(_00900_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  buf(_00904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  buf(_00916_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(_00920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(_00929_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(_00941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(_00947_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  buf(_00953_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  buf(_00961_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  buf(_00963_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  buf(_00971_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  buf(_00973_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  buf(_00978_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  buf(_00981_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  buf(_00983_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  buf(_00985_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  buf(_00988_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  buf(_00990_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  buf(_00992_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  buf(_00995_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  buf(_00996_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  buf(_01000_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  buf(_01013_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  buf(_01015_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(_01016_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  buf(_01018_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(_01020_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  buf(_01022_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(_01023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  buf(_01025_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(_01027_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  buf(_01029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(_01030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  buf(_01032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(_01034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  buf(_01036_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(_01039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  buf(_01042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  buf(_01185_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(_01187_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(_01189_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(_01191_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(_01193_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(_01195_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(_01197_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(_01224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(_01226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans );
  buf(_01229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(_01234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event );
  buf(_01238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(_01249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(_01252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(_01259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  buf(_01263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(_01265_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(_01268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(_01284_, t2_i);
  buf(_01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  buf(_01291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(_01295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(_01299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  buf(_01303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(_01307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(_01345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(_01369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(_01374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(_01383_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(_01389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(_01405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(_01409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(_01412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(_01415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(_01421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(_01423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(_01432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(_01441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(_01444_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(_01447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(_01450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(_01453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(_01456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(_01459_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(_01469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(_01473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(_01476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(_01479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(_01482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(_01485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(_01488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(_01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(_01589_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(_01597_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(_01606_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(_01609_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(_01617_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(_01620_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(_01627_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(_01678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(_01703_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(_01710_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(_01714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(_01718_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(_01722_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(_01728_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(_01740_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(_01866_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  buf(_01880_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  buf(_01904_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  buf(_01977_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  buf(_01981_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  buf(_01983_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  buf(_01985_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  buf(_01988_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  buf(_01991_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  buf(_01993_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  buf(_01995_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  buf(_01998_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  buf(_02000_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  buf(_02002_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  buf(_02005_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  buf(_02008_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  buf(_02091_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  buf(_02093_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  buf(_02096_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  buf(_02212_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  buf(_02214_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  buf(_02216_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  buf(_02218_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  buf(_02220_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  buf(_02222_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  buf(_02224_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  buf(_02586_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(_02809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(_03047_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(_03049_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(_03074_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(_03076_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(_03078_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(_03080_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(_03082_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(_03083_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(_03085_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(_03089_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(_03090_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(_03113_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(_03116_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(_03119_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(_03122_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(_03128_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(_03131_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(_03135_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  buf(_03138_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  buf(_03167_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(_03169_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(_03172_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(_03174_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(_03177_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(_03181_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(_03183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(_03185_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(_03188_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(_03194_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(_03268_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  buf(_03270_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  buf(_03272_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  buf(_03274_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  buf(_03276_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  buf(_03278_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  buf(_03280_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  buf(_03282_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(_03284_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(_03285_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(_03287_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(_03291_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(_03293_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(_03295_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(_03297_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(_03299_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(_03301_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(_03308_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(_03313_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(_03330_, \oc8051_top_1.oc8051_decoder1.state [1]);
  buf(_03332_, \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(_03341_, \oc8051_top_1.oc8051_decoder1.op [7]);
  buf(_03355_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(_03358_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  buf(_03360_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  buf(_03362_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2]);
  buf(_03364_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  buf(_03366_, \oc8051_top_1.oc8051_decoder1.wr );
  buf(_03783_, \oc8051_top_1.oc8051_decoder1.state [0]);
  buf(_03785_, \oc8051_top_1.oc8051_decoder1.op [0]);
  buf(_03788_, \oc8051_top_1.oc8051_decoder1.op [1]);
  buf(_03791_, \oc8051_top_1.oc8051_decoder1.op [2]);
  buf(_03793_, \oc8051_top_1.oc8051_decoder1.op [3]);
  buf(_03796_, \oc8051_top_1.oc8051_decoder1.op [4]);
  buf(_03799_, \oc8051_top_1.oc8051_decoder1.op [5]);
  buf(_03802_, \oc8051_top_1.oc8051_decoder1.op [6]);
  buf(_03809_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  buf(_03811_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  buf(_03813_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  buf(_03815_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  buf(_03817_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0]);
  buf(_03819_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1]);
  buf(_03821_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  buf(_03823_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  buf(_04340_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  buf(_04342_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  buf(_04344_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  buf(_04349_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  buf(_04358_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(_04361_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  buf(_04368_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(_04371_, \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(_04376_, \oc8051_top_1.oc8051_rom1.ea_int );
  buf(_04386_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(_04388_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  buf(_04390_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  buf(_04412_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  buf(_04414_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  buf(_04417_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  buf(_04442_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  buf(_04449_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  buf(_04458_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  buf(_04466_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(_35657_[15], _04469_);
  buf(_04471_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(_35658_[15], _04473_);
  buf(_04510_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  buf(_04514_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  buf(_04617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  buf(_04636_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  buf(_04637_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  buf(_04658_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  buf(_04660_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  buf(_04666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(_37361_[0], _04678_);
  buf(_04680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(_04682_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  buf(_04684_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(_04686_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  buf(_04689_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  buf(_04693_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  buf(_04696_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(_04717_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(_04720_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(_04724_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(_04728_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(_04731_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(_04736_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(_04740_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(_04744_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(_04748_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(_04751_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(_04754_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(_04757_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(_04761_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(_04764_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(_04768_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(_04772_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(_04774_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(_04778_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(_04782_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(_04786_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(_04790_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(_04794_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(_04798_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(_04801_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(_04811_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  buf(_04814_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  buf(_04817_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  buf(_04820_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  buf(_04861_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  buf(_04868_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  buf(_04877_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  buf(_04879_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  buf(_04889_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(_04893_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(_04897_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(_04901_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(_04905_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(_04908_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(_04912_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(_04945_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  buf(_04950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  buf(_04956_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  buf(_04960_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  buf(_05028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(_05031_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(_05034_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(_05036_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(_05040_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(_05043_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(_05046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(_05048_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(_05051_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(_05054_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(_05057_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(_05060_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(_05063_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(_05066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(_05069_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(_35657_[0], _05072_);
  buf(_35657_[1], _05074_);
  buf(_35657_[2], _05076_);
  buf(_35657_[3], _05078_);
  buf(_35657_[4], _05079_);
  buf(_35657_[5], _05081_);
  buf(_35657_[6], _05083_);
  buf(_35657_[7], _05085_);
  buf(_35657_[8], _05087_);
  buf(_35657_[9], _05089_);
  buf(_35657_[10], _05091_);
  buf(_35657_[11], _05093_);
  buf(_35657_[12], _05095_);
  buf(_35657_[13], _05097_);
  buf(_35657_[14], _05099_);
  buf(_05101_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(_05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(_05107_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(_05110_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(_05112_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(_05115_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(_05118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(_05121_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(_05124_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(_05127_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(_05130_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(_05133_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(_05136_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(_05139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(_05142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(_35658_[0], _05145_);
  buf(_35658_[1], _05147_);
  buf(_35658_[2], _05149_);
  buf(_35658_[3], _05151_);
  buf(_35658_[4], _05153_);
  buf(_35658_[5], _05155_);
  buf(_35658_[6], _05157_);
  buf(_35658_[7], _05159_);
  buf(_35658_[8], _05161_);
  buf(_35658_[9], _05163_);
  buf(_35658_[10], _05165_);
  buf(_35658_[11], _05167_);
  buf(_35658_[12], _05170_);
  buf(_35658_[13], _05172_);
  buf(_35658_[14], _05174_);
  buf(_05339_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  buf(_05341_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  buf(_05342_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  buf(_05344_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  buf(_05346_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  buf(_05348_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  buf(_05350_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  buf(_05355_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  buf(_05359_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  buf(_05362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  buf(_05367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  buf(_05375_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  buf(_05379_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  buf(_05382_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  buf(_05388_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  buf(_05390_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  buf(_05392_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  buf(_05394_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  buf(_05398_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  buf(_05403_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  buf(_05405_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  buf(_05407_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  buf(_05409_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  buf(_05413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  buf(_05415_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  buf(_05420_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  buf(_05422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  buf(_05427_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  buf(_05429_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  buf(_05433_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  buf(_05439_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  buf(_05443_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  buf(_05446_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  buf(_05448_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  buf(_05450_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  buf(_05452_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  buf(_05453_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  buf(_05455_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  buf(_05457_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  buf(_05459_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  buf(_05461_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  buf(_05464_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  buf(_05468_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  buf(_05472_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  buf(_05478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  buf(_05491_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  buf(_05493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  buf(_05497_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  buf(_05608_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  buf(_05614_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  buf(_05618_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  buf(_05623_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  buf(_05627_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  buf(_05631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  buf(_05636_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  buf(_05897_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  buf(_05900_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  buf(_05915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  buf(_05918_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  buf(_05921_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  buf(_05924_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  buf(_05927_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  buf(_05931_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  buf(_05935_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  buf(_05937_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  buf(_05942_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  buf(_05946_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  buf(_05949_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  buf(_05954_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  buf(_05957_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  buf(_05959_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  buf(_05963_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  buf(_05964_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  buf(_05967_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  buf(_06040_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  buf(_06042_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  buf(_06043_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  buf(_06045_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  buf(_06047_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  buf(_06049_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  buf(_06051_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  buf(_06059_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  buf(_06061_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  buf(_06063_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  buf(_06065_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  buf(_06067_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  buf(_06072_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  buf(_06091_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(_06094_, \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(_06101_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  buf(_06114_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(_06117_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(_06119_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(_06122_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(_06125_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(_06128_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(_06131_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(_06133_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  buf(_06135_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  buf(_06165_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0]);
  buf(_06167_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1]);
  buf(_06169_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2]);
  buf(_06170_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3]);
  buf(_06172_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4]);
  buf(_06174_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5]);
  buf(_06176_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6]);
  buf(_06243_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  buf(_06264_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  buf(_06269_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  buf(_06359_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  buf(_06376_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(_06380_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  buf(_06384_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(_06388_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(_06392_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(_06398_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  buf(_06402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  buf(_06406_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  buf(_06411_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  buf(_06415_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  buf(_06422_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  buf(_06426_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  buf(_06438_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  buf(_06441_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  buf(_06444_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  buf(_06476_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  buf(_06479_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  buf(_06482_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  buf(_06489_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  buf(_06492_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  buf(_06495_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  buf(_06503_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(_06506_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(_06509_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(_06512_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(_06516_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(_06519_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(_06522_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(_06525_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(_06528_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(_06531_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(_06534_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(_06537_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(_06540_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(_06543_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(_06546_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(_06549_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(_06552_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(_06555_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(_06558_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(_06561_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(_06564_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(_06567_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(_06570_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(_06573_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(_06577_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(_06580_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(_06583_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(_06586_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(_06589_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  buf(_06592_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  buf(_06595_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  buf(_06598_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  buf(_06601_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  buf(_06604_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  buf(_06607_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  buf(_06610_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  buf(_06613_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  buf(_06616_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  buf(_06619_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  buf(_06622_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  buf(_06625_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  buf(_06628_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  buf(_06713_, p0_in[7]);
  buf(_06938_, \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  buf(_06940_, \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  buf(_06971_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  buf(_07283_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  buf(_07539_, word_in[7]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07543_);
  buf(_07546_, \oc8051_symbolic_cxrom1.regvalid [11]);
  buf(_07549_, word_in[15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07552_);
  buf(_07558_, word_in[23]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07561_);
  buf(_07569_, word_in[31]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [31], _07572_);
  buf(_07605_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  buf(_07607_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  buf(_07638_, \oc8051_symbolic_cxrom1.regvalid [8]);
  buf(_33904_[7], _07650_);
  buf(_07658_, \oc8051_symbolic_cxrom1.regvalid [0]);
  buf(_33955_, _07676_);
  buf(_07679_, \oc8051_symbolic_cxrom1.regvalid [1]);
  buf(_33505_[13], _07683_);
  buf(_07690_, \oc8051_symbolic_cxrom1.regvalid [14]);
  buf(_33505_[1], _07704_);
  buf(_07708_, \oc8051_symbolic_cxrom1.regvalid [2]);
  buf(_33505_[11], _07718_);
  buf(_33505_[8], _07724_);
  buf(_07726_, \oc8051_symbolic_cxrom1.regvalid [12]);
  buf(_07731_, \oc8051_symbolic_cxrom1.regvalid [9]);
  buf(_33505_[2], _07740_);
  buf(_07743_, \oc8051_symbolic_cxrom1.regvalid [3]);
  buf(_33505_[3], _07777_);
  buf(_07780_, \oc8051_symbolic_cxrom1.regvalid [4]);
  buf(_33505_[15], _07787_);
  buf(_33505_[4], _07814_);
  buf(_07817_, \oc8051_symbolic_cxrom1.regvalid [5]);
  buf(_33505_[9], _07832_);
  buf(_07835_, \oc8051_symbolic_cxrom1.regvalid [10]);
  buf(_33505_[5], _07860_);
  buf(_07863_, \oc8051_symbolic_cxrom1.regvalid [6]);
  buf(_33505_[12], _07873_);
  buf(_33505_[7], _07878_);
  buf(_07880_, \oc8051_symbolic_cxrom1.regvalid [13]);
  buf(_33505_[14], _07897_);
  buf(_07902_, \oc8051_symbolic_cxrom1.regvalid [15]);
  buf(_33505_[6], _07911_);
  buf(_07915_, \oc8051_symbolic_cxrom1.regvalid [7]);
  buf(_33505_[10], _07929_);
  buf(_08006_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  buf(_08008_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  buf(_08010_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  buf(_08012_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  buf(_08014_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  buf(_08016_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  buf(_08018_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  buf(_08020_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  buf(_08022_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  buf(_08025_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  buf(_08027_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  buf(_08029_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  buf(_08031_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  buf(_08033_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  buf(_08035_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  buf(_08037_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  buf(_33880_[7], _08109_);
  buf(_33908_[7], _08135_);
  buf(_33912_[7], _08161_);
  buf(_33916_[7], _08178_);
  buf(_33920_[7], _08204_);
  buf(_33924_[7], _08217_);
  buf(_33928_[7], _08230_);
  buf(_33932_[7], _08244_);
  buf(_33936_[7], _08269_);
  buf(_33940_[7], _08282_);
  buf(_33884_[7], _08297_);
  buf(_33888_[7], _08310_);
  buf(_33892_[7], _08327_);
  buf(_33896_[7], _08341_);
  buf(_33900_[7], _08354_);
  buf(_33904_[0], _08367_);
  buf(_33904_[1], _08371_);
  buf(_33904_[2], _08375_);
  buf(_33904_[3], _08380_);
  buf(_33904_[4], _08384_);
  buf(_33904_[5], _08388_);
  buf(_33904_[6], _08392_);
  buf(_08395_, word_in[0]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [0], _08398_);
  buf(_08400_, word_in[1]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [1], _08403_);
  buf(_08405_, word_in[2]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [2], _08408_);
  buf(_08410_, word_in[3]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [3], _08412_);
  buf(_08414_, word_in[4]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [4], _08416_);
  buf(_08418_, word_in[5]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [5], _08420_);
  buf(_08422_, word_in[6]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [6], _08424_);
  buf(_08426_, word_in[8]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [8], _08429_);
  buf(_08431_, word_in[9]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [9], _08434_);
  buf(_08436_, word_in[10]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [10], _08439_);
  buf(_08441_, word_in[11]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [11], _08445_);
  buf(_08447_, word_in[12]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [12], _08450_);
  buf(_08452_, word_in[13]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [13], _08455_);
  buf(_08457_, word_in[14]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [14], _08460_);
  buf(_08469_, word_in[16]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [16], _08472_);
  buf(_08474_, word_in[17]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [17], _08477_);
  buf(_08479_, word_in[18]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [18], _08482_);
  buf(_08484_, word_in[19]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [19], _08487_);
  buf(_08489_, word_in[20]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [20], _08492_);
  buf(_08494_, word_in[21]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [21], _08497_);
  buf(_08499_, word_in[22]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [22], _08502_);
  buf(_08504_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  buf(_08506_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  buf(_08510_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  buf(_08512_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  buf(_08515_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  buf(_08517_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  buf(_08520_, word_in[24]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [24], _08523_);
  buf(_08525_, word_in[25]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [25], _08528_);
  buf(_08530_, word_in[26]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [26], _08533_);
  buf(_08535_, word_in[27]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [27], _08538_);
  buf(_08540_, word_in[28]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [28], _08543_);
  buf(_08545_, word_in[29]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [29], _08548_);
  buf(_08550_, word_in[30]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [30], _08553_);
  buf(_08556_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  buf(_08558_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  buf(_08565_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  buf(_08567_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  buf(_08570_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  buf(_08573_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  buf(_08576_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  buf(_08578_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  buf(_08696_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  buf(_08699_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  buf(_08702_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  buf(_08704_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  buf(_08707_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  buf(_08709_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  buf(_08711_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  buf(_08713_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  buf(_08729_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  buf(_08731_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  buf(_08734_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  buf(_08736_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  buf(_08809_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  buf(_08811_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  buf(_08814_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  buf(_08816_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  buf(_08818_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  buf(_08820_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  buf(_08825_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  buf(_08827_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  buf(_08830_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  buf(_08832_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  buf(_08835_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  buf(_08837_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  buf(_08847_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  buf(_08849_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  buf(_08852_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  buf(_08854_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  buf(_08859_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  buf(_08861_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  buf(_08864_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  buf(_08866_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  buf(_08876_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  buf(_08878_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  buf(_08895_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  buf(_08898_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  buf(_08900_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  buf(_08902_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  buf(_08905_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  buf(_08907_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  buf(_08911_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  buf(_08913_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  buf(_08916_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  buf(_08918_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  buf(_08921_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  buf(_08923_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  buf(_08926_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  buf(_08928_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  buf(_08932_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  buf(_08934_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  buf(_08936_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  buf(_08938_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  buf(_08942_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  buf(_08944_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  buf(_08950_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  buf(_08952_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  buf(_08969_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  buf(_08971_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  buf(_08980_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  buf(_08982_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  buf(_08986_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  buf(_08988_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  buf(_08993_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  buf(_08995_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  buf(_08998_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  buf(_09000_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  buf(_09003_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  buf(_09005_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  buf(_09010_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  buf(_09012_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  buf(_09016_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  buf(_09018_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  buf(_09021_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  buf(_09023_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  buf(_09032_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  buf(_09034_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  buf(_09037_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  buf(_09039_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  buf(_09043_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  buf(_09045_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  buf(_09048_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  buf(_09050_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  buf(_09054_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  buf(_09056_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  buf(_09058_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  buf(_09060_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  buf(_33900_[0], _09144_);
  buf(_33900_[1], _09147_);
  buf(_33900_[2], _09150_);
  buf(_33900_[3], _09153_);
  buf(_33900_[4], _09156_);
  buf(_33900_[5], _09160_);
  buf(_33900_[6], _09163_);
  buf(_33896_[0], _09180_);
  buf(_33896_[1], _09183_);
  buf(_33896_[2], _09186_);
  buf(_33896_[3], _09189_);
  buf(_33896_[4], _09192_);
  buf(_33896_[5], _09195_);
  buf(_33896_[6], _09198_);
  buf(_33892_[0], _09216_);
  buf(_33892_[1], _09219_);
  buf(_33892_[2], _09222_);
  buf(_33892_[3], _09225_);
  buf(_33892_[4], _09228_);
  buf(_33892_[5], _09231_);
  buf(_33892_[6], _09234_);
  buf(_33888_[0], _09251_);
  buf(_33888_[1], _09254_);
  buf(_33888_[2], _09257_);
  buf(_33888_[3], _09261_);
  buf(_33888_[4], _09264_);
  buf(_33888_[5], _09267_);
  buf(_33888_[6], _09270_);
  buf(_33884_[0], _09287_);
  buf(_33884_[1], _09290_);
  buf(_33884_[2], _09293_);
  buf(_33884_[3], _09296_);
  buf(_33884_[4], _09299_);
  buf(_33884_[5], _09302_);
  buf(_33884_[6], _09305_);
  buf(_33940_[0], _09324_);
  buf(_33940_[1], _09327_);
  buf(_33940_[2], _09330_);
  buf(_33940_[3], _09333_);
  buf(_33940_[4], _09336_);
  buf(_33940_[5], _09339_);
  buf(_33940_[6], _09342_);
  buf(_33936_[0], _09359_);
  buf(_33936_[1], _09363_);
  buf(_33936_[2], _09366_);
  buf(_33936_[3], _09369_);
  buf(_33936_[4], _09372_);
  buf(_33936_[5], _09375_);
  buf(_33936_[6], _09378_);
  buf(_33932_[0], _09395_);
  buf(_33932_[1], _09398_);
  buf(_33932_[2], _09401_);
  buf(_33932_[3], _09404_);
  buf(_33932_[4], _09407_);
  buf(_33932_[5], _09410_);
  buf(_33932_[6], _09413_);
  buf(_33928_[0], _09431_);
  buf(_33928_[1], _09434_);
  buf(_33928_[2], _09437_);
  buf(_33928_[3], _09440_);
  buf(_33928_[4], _09443_);
  buf(_33928_[5], _09446_);
  buf(_33928_[6], _09449_);
  buf(_33924_[0], _09467_);
  buf(_33924_[1], _09470_);
  buf(_33924_[2], _09473_);
  buf(_33924_[3], _09476_);
  buf(_33924_[4], _09479_);
  buf(_33924_[5], _09482_);
  buf(_33924_[6], _09485_);
  buf(_33920_[0], _09502_);
  buf(_33920_[1], _09505_);
  buf(_33920_[2], _09508_);
  buf(_33920_[3], _09511_);
  buf(_33920_[4], _09514_);
  buf(_33920_[5], _09518_);
  buf(_33920_[6], _09521_);
  buf(_33916_[0], _09538_);
  buf(_33916_[1], _09541_);
  buf(_33916_[2], _09544_);
  buf(_33916_[3], _09547_);
  buf(_33916_[4], _09550_);
  buf(_33916_[5], _09553_);
  buf(_33916_[6], _09556_);
  buf(_33912_[0], _09574_);
  buf(_33912_[1], _09577_);
  buf(_33912_[2], _09580_);
  buf(_33912_[3], _09583_);
  buf(_33912_[4], _09586_);
  buf(_33912_[5], _09589_);
  buf(_33912_[6], _09592_);
  buf(_33908_[0], _09609_);
  buf(_33908_[1], _09612_);
  buf(_33908_[2], _09615_);
  buf(_33908_[3], _09619_);
  buf(_33908_[4], _09622_);
  buf(_33908_[5], _09625_);
  buf(_33908_[6], _09628_);
  buf(_09644_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  buf(_09646_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  buf(_09648_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  buf(_09649_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  buf(_09651_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  buf(_33880_[0], _09654_);
  buf(_33880_[1], _09657_);
  buf(_33880_[2], _09660_);
  buf(_33880_[3], _09663_);
  buf(_33880_[4], _09666_);
  buf(_33880_[5], _09669_);
  buf(_33880_[6], _09673_);
  buf(_09696_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  buf(_09698_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  buf(_09700_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  buf(_09702_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  buf(_09704_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  buf(_10219_, first_instr);
  buf(property_invalid, _10258_);
  buf(_00000_, _10272_);
endmodule
