
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jc, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_05542_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_05543_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_05544_, _05543_, _05542_);
  not (_05545_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_05546_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_05547_, _05546_, _05545_);
  not (_05548_, _05547_);
  nor (_05549_, _05548_, _05544_);
  nor (_05550_, _05549_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_05551_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not (_05552_, rst);
  not (_05553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_05554_, _05550_, _05553_);
  and (_05555_, _05554_, _05552_);
  and (_00395_, _05555_, _05551_);
  not (_05556_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_05557_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _05556_);
  and (_05558_, _05557_, _05552_);
  not (_05559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_05560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor (_05561_, _05560_, _05559_);
  and (_05562_, _05561_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_05563_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_05564_, _05563_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not (_05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_05566_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _05565_);
  and (_05567_, _05566_, _05564_);
  and (_05568_, _05567_, _05562_);
  and (_05569_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not (_05570_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_05571_, _05560_, _05570_);
  and (_05572_, _05571_, _05569_);
  not (_05573_, _05560_);
  and (_05574_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_05575_, _05574_, _05573_);
  nor (_05576_, _05575_, _05572_);
  nor (_05577_, _05576_, _05562_);
  or (_05579_, _05577_, _05568_);
  and (_05580_, _05560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_05582_, _05580_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_05583_, _05582_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_05584_, _05583_, _05579_);
  and (_05585_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_05586_, _05582_, _05568_);
  or (_05587_, _05586_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_05588_, _05587_, _05585_);
  and (_05589_, _05588_, _05584_);
  or (_01099_, _05589_, _05558_);
  nor (_05590_, rst, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_05591_, _05590_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_05592_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  not (_05593_, _05562_);
  nor (_05594_, _05567_, _05593_);
  and (_05595_, _05594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor (_05596_, _05562_, _05572_);
  or (_05597_, _05596_, _05595_);
  and (_05598_, _05597_, _05592_);
  not (_05599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_05600_, _05586_, _05599_);
  or (_05601_, _05600_, _05598_);
  nand (_05602_, _05582_, _05599_);
  and (_05603_, _05602_, _05585_);
  and (_05604_, _05603_, _05601_);
  or (_03276_, _05604_, _05591_);
  not (_05605_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_05606_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_05607_, _05606_, _05605_);
  and (_05608_, _05607_, _05547_);
  not (_05609_, _05608_);
  not (_05611_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_05612_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_05613_, _05612_, _05542_);
  or (_05614_, _05613_, _05611_);
  not (_05615_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_05616_, _05543_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or (_05617_, _05616_, _05615_);
  and (_05618_, _05617_, _05614_);
  and (_05619_, _05612_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_05620_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_05621_, _05620_, _05618_);
  not (_05622_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_05623_, _05622_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_05624_, _05623_, _05542_);
  not (_05625_, _05624_);
  nand (_05626_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_05627_, _05612_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_05628_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nand (_05629_, _05628_, _05626_);
  nor (_05630_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_05631_, _05630_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  not (_05632_, _05631_);
  and (_05633_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_05634_, _05633_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_05635_, _05634_, _05629_);
  or (_05636_, _05635_, _05621_);
  or (_05637_, _05636_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05638_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_05639_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _05638_);
  not (_05640_, _05639_);
  and (_05641_, _05640_, _05637_);
  or (_05642_, _05641_, _05609_);
  not (_05643_, _05607_);
  nor (_05644_, _05547_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_05645_, _05644_, _05643_);
  nand (_05646_, _05645_, _05642_);
  nand (_05647_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_05648_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_05649_, _05648_, _05647_);
  not (_05650_, _05616_);
  nand (_05651_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not (_05652_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_05653_, _05631_, _05652_);
  and (_05654_, _05653_, _05651_);
  nand (_05655_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_05656_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_05657_, _05613_, _05656_);
  and (_05658_, _05657_, _05655_);
  and (_05659_, _05658_, _05654_);
  and (_05660_, _05659_, _05649_);
  or (_05661_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_05662_, _05661_, _05660_);
  and (_05663_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05664_, _05663_);
  and (_05665_, _05664_, _05662_);
  nand (_05666_, _05665_, _05608_);
  nor (_05667_, _05547_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_05668_, _05667_, _05643_);
  and (_05669_, _05668_, _05666_);
  and (_05670_, _05669_, _05646_);
  not (_05671_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_05673_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nand (_05674_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_05675_, _05674_, _05673_);
  nand (_05676_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  not (_05677_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_05678_, _05613_, _05677_);
  and (_05679_, _05678_, _05676_);
  nand (_05680_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_05681_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_05682_, _05681_, _05680_);
  and (_05683_, _05682_, _05679_);
  nand (_05684_, _05683_, _05675_);
  nand (_05685_, _05684_, _05671_);
  nand (_05686_, _05685_, _05638_);
  nor (_05687_, _05638_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  not (_05688_, _05687_);
  and (_05689_, _05688_, _05686_);
  or (_05690_, _05689_, _05609_);
  nor (_05691_, _05547_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_05692_, _05691_, _05643_);
  and (_05693_, _05692_, _05690_);
  nand (_05694_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  not (_05695_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_05696_, _05631_, _05695_);
  and (_05697_, _05696_, _05694_);
  nand (_05698_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not (_05699_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_05700_, _05613_, _05699_);
  and (_05701_, _05700_, _05698_);
  nand (_05702_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand (_05703_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_05704_, _05703_, _05702_);
  and (_05705_, _05704_, _05701_);
  and (_05706_, _05705_, _05697_);
  or (_05707_, _05706_, _05661_);
  and (_05708_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05709_, _05708_);
  nand (_05710_, _05709_, _05707_);
  or (_05711_, _05710_, _05609_);
  nor (_05712_, _05547_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_05713_, _05712_, _05643_);
  nand (_05714_, _05713_, _05711_);
  and (_05715_, _05714_, _05693_);
  and (_05716_, _05715_, _05670_);
  and (_05717_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_05718_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_05719_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_05720_, _05719_, _05718_);
  or (_05721_, _05720_, _05717_);
  and (_05722_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_05723_, _05722_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_05724_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not (_05725_, _05613_);
  and (_05726_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_05727_, _05726_, _05724_);
  or (_05728_, _05727_, _05723_);
  or (_05729_, _05728_, _05721_);
  or (_05730_, _05729_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_05731_, _05638_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  not (_05732_, _05731_);
  and (_05733_, _05732_, _05730_);
  or (_05734_, _05733_, _05609_);
  nor (_05735_, _05547_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_05736_, _05735_, _05643_);
  and (_05737_, _05736_, _05734_);
  not (_05738_, _05737_);
  nor (_05739_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_05740_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_05741_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_05742_, _05741_, _05740_);
  not (_05743_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_05744_, _05616_, _05743_);
  nand (_05745_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_05746_, _05745_, _05744_);
  nand (_05747_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_05748_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or (_05749_, _05613_, _05748_);
  and (_05750_, _05749_, _05747_);
  and (_05751_, _05750_, _05746_);
  nand (_05752_, _05751_, _05742_);
  nand (_05753_, _05752_, _05739_);
  and (_05754_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not (_05755_, _05754_);
  and (_05756_, _05755_, _05753_);
  nand (_05757_, _05756_, _05608_);
  nor (_05758_, _05547_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_05759_, _05758_, _05643_);
  and (_05760_, _05759_, _05757_);
  not (_05761_, _05760_);
  not (_05762_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or (_05763_, _05613_, _05762_);
  not (_05765_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_05766_, _05624_, _05765_);
  and (_05767_, _05766_, _05763_);
  not (_05768_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_05769_, _05616_, _05768_);
  not (_05770_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_05771_, _05631_, _05770_);
  and (_05772_, _05771_, _05769_);
  and (_05773_, _05772_, _05767_);
  nand (_05774_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_05775_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_05776_, _05775_, _05774_);
  and (_05777_, _05776_, _05773_);
  or (_05778_, _05777_, _05661_);
  and (_05779_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05780_, _05779_);
  nand (_05781_, _05780_, _05778_);
  or (_05782_, _05781_, _05609_);
  nor (_05783_, _05547_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_05784_, _05783_, _05643_);
  nand (_05785_, _05784_, _05782_);
  not (_05786_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_05787_, _05613_, _05786_);
  not (_05788_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_05789_, _05624_, _05788_);
  and (_05790_, _05789_, _05787_);
  not (_05791_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_05792_, _05616_, _05791_);
  nand (_05793_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_05794_, _05793_, _05792_);
  and (_05795_, _05794_, _05790_);
  nand (_05796_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_05797_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_05798_, _05797_, _05796_);
  and (_05799_, _05798_, _05795_);
  or (_05800_, _05799_, _05661_);
  and (_05801_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05802_, _05801_);
  nand (_05803_, _05802_, _05800_);
  or (_05804_, _05803_, _05609_);
  nor (_05805_, _05547_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_05806_, _05805_, _05643_);
  nand (_05807_, _05806_, _05804_);
  and (_05808_, _05807_, _05785_);
  and (_05809_, _05808_, _05761_);
  and (_05810_, _05809_, _05738_);
  and (_05811_, _05810_, _05716_);
  and (_05812_, _05784_, _05782_);
  nor (_05813_, _05807_, _05760_);
  and (_05814_, _05813_, _05812_);
  and (_05815_, _05737_, _05716_);
  and (_05816_, _05815_, _05814_);
  or (_05817_, _05816_, _05811_);
  not (_05818_, _05669_);
  not (_05819_, _05646_);
  not (_05820_, _05714_);
  nor (_05821_, _05820_, _05693_);
  and (_05822_, _05821_, _05819_);
  and (_05823_, _05822_, _05818_);
  and (_05824_, _05809_, _05737_);
  and (_05825_, _05824_, _05823_);
  and (_05826_, _05807_, _05812_);
  and (_05827_, _05826_, _05760_);
  and (_05828_, _05827_, _05737_);
  and (_05829_, _05828_, _05823_);
  and (_05830_, _05814_, _05738_);
  and (_05831_, _05830_, _05823_);
  nor (_05832_, _05831_, _05829_);
  not (_05833_, _05832_);
  or (_05834_, _05833_, _05825_);
  or (_05835_, _05834_, _05817_);
  not (_05836_, _05807_);
  and (_05837_, _05836_, _05760_);
  and (_05838_, _05837_, _05815_);
  and (_05839_, _05826_, _05761_);
  and (_05840_, _05839_, _05737_);
  and (_05841_, _05840_, _05823_);
  and (_05842_, _05815_, _05809_);
  or (_05843_, _05842_, _05841_);
  or (_05844_, _05843_, _05838_);
  and (_05845_, _05830_, _05716_);
  and (_05846_, _05814_, _05737_);
  and (_05847_, _05846_, _05823_);
  or (_05848_, _05847_, _05845_);
  and (_05849_, _05818_, _05646_);
  and (_05850_, _05849_, _05821_);
  and (_05851_, _05850_, _05814_);
  nor (_05852_, _05807_, _05812_);
  and (_05853_, _05852_, _05760_);
  and (_05854_, _05853_, _05738_);
  and (_05855_, _05854_, _05822_);
  nor (_05856_, _05855_, _05851_);
  and (_05857_, _05839_, _05738_);
  and (_05858_, _05857_, _05716_);
  and (_05859_, _05852_, _05761_);
  and (_05860_, _05859_, _05738_);
  and (_05861_, _05860_, _05822_);
  nor (_05862_, _05861_, _05858_);
  nand (_05864_, _05862_, _05856_);
  or (_05865_, _05864_, _05848_);
  or (_05867_, _05865_, _05844_);
  or (_05868_, _05867_, _05835_);
  and (_05869_, _05821_, _05670_);
  and (_05870_, _05869_, _05737_);
  and (_05872_, _05857_, _05820_);
  or (_05873_, _05872_, _05870_);
  nor (_05874_, _05737_, _05646_);
  and (_05875_, _05874_, _05715_);
  and (_05876_, _05875_, _05839_);
  and (_05877_, _05859_, _05737_);
  and (_05878_, _05877_, _05822_);
  or (_05879_, _05878_, _05876_);
  or (_05880_, _05879_, _05873_);
  or (_05881_, _05880_, _05868_);
  and (_05882_, _05881_, _05547_);
  and (_05883_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_05884_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_05885_, \oc8051_top_1.oc8051_decoder1.state [1], _05545_);
  and (_05886_, _05885_, _05884_);
  and (_05887_, _05850_, _05824_);
  and (_05888_, _05887_, _05886_);
  or (_05889_, _05870_, _05825_);
  and (_05890_, _05889_, _05886_);
  not (_05891_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_05892_, \oc8051_top_1.oc8051_decoder1.state [0], _05545_);
  and (_05893_, _05892_, _05891_);
  and (_05894_, _05849_, _05715_);
  and (_05895_, _05827_, _05738_);
  and (_05896_, _05895_, _05894_);
  and (_05897_, _05894_, _05857_);
  nor (_05898_, _05897_, _05896_);
  not (_05900_, _05898_);
  and (_05901_, _05900_, _05893_);
  or (_05902_, _05901_, _05890_);
  or (_05903_, _05902_, _05888_);
  or (_05904_, _05903_, _05883_);
  or (_05905_, _05904_, _05882_);
  and (_04490_, _05905_, _05552_);
  or (_05906_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not (_05907_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_05908_, _05550_, _05907_);
  and (_05909_, _05908_, _05552_);
  and (_05764_, _05909_, _05906_);
  not (_05910_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_05911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor (_05912_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_05913_, _05912_, _05911_);
  or (_05914_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor (_05915_, _05914_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_05916_, _05915_, _05913_);
  and (_05917_, _05916_, _05910_);
  and (_05918_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_05919_, _05918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_07307_, _05919_, _05552_);
  or (_05920_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not (_05921_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_05922_, _05550_, _05921_);
  and (_05923_, _05922_, _05552_);
  and (_08287_, _05923_, _05920_);
  and (_05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_05925_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_05926_, _05925_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_05927_, _05926_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_05928_, _05927_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_05930_, _05928_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_05931_, _05930_);
  not (_05933_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05934_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05545_);
  and (_05935_, _05934_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_05936_, _05935_, _05933_);
  not (_05937_, _05936_);
  nor (_05938_, _05928_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_05939_, _05938_, _05937_);
  and (_05940_, _05939_, _05931_);
  not (_05941_, _05940_);
  not (_05942_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_05943_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05545_);
  and (_05944_, _05943_, _05942_);
  and (_05945_, _05944_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05946_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  not (_05947_, _05946_);
  and (_05948_, _05944_, _05933_);
  and (_05949_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  not (_05950_, _05949_);
  nor (_05951_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_05952_, _05951_, _05934_);
  and (_05953_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_05954_, _05935_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor (_05955_, _05954_, _05953_);
  and (_05956_, _05955_, _05950_);
  and (_05957_, _05956_, _05947_);
  and (_05958_, _05957_, _05941_);
  not (_05959_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_05960_, _05930_, _05959_);
  and (_05961_, _05930_, _05959_);
  nor (_05962_, _05961_, _05960_);
  nor (_05963_, _05962_, _05937_);
  not (_05964_, _05963_);
  and (_05965_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_05966_, _05945_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and (_05967_, _05948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or (_05968_, _05967_, _05966_);
  or (_05969_, _05968_, _05954_);
  nor (_05970_, _05969_, _05965_);
  and (_05971_, _05970_, _05964_);
  and (_05972_, _05971_, _05958_);
  not (_05973_, _05927_);
  nor (_05974_, _05926_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_05975_, _05974_, _05937_);
  and (_05976_, _05975_, _05973_);
  not (_05977_, _05976_);
  and (_05978_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  not (_05979_, _05978_);
  and (_05980_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_05981_, _05980_, _05954_);
  and (_05982_, _05981_, _05979_);
  and (_05983_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_05984_, _05951_, _05942_);
  or (_05985_, _05984_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_05986_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_05987_, _05986_, _05983_);
  and (_05988_, _05987_, _05982_);
  and (_05989_, _05988_, _05977_);
  not (_05990_, _05928_);
  nor (_05991_, _05927_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_05992_, _05991_, _05937_);
  and (_05993_, _05992_, _05990_);
  not (_05994_, _05993_);
  and (_05995_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_05996_, _05945_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_05997_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  or (_05998_, _05997_, _05996_);
  or (_05999_, _05998_, _05954_);
  nor (_06000_, _05999_, _05995_);
  and (_06001_, _06000_, _05994_);
  and (_06002_, _06001_, _05989_);
  and (_06003_, _06002_, _05972_);
  and (_06004_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_06006_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  nor (_06008_, _06006_, _06004_);
  not (_06009_, _05926_);
  nor (_06010_, _05925_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_06011_, _06010_, _05937_);
  and (_06012_, _06011_, _06009_);
  and (_06014_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and (_06015_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_06016_, _06015_, _06014_);
  not (_06018_, _06016_);
  nor (_06019_, _06018_, _06012_);
  and (_06020_, _06019_, _06008_);
  and (_06021_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  and (_06022_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_06023_, _06022_, _06021_);
  and (_06024_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  not (_06025_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_06026_, _05936_, _06025_);
  and (_06027_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  or (_06028_, _06027_, _06026_);
  nor (_06029_, _06028_, _06024_);
  and (_06030_, _06029_, _06023_);
  not (_06031_, _06030_);
  nor (_06032_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_06033_, _06032_, _05924_);
  and (_06034_, _06033_, _05936_);
  and (_06035_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_06037_, _06035_, _06034_);
  and (_06038_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_06039_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_06040_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_06041_, _06040_, _06039_);
  nor (_06042_, _06041_, _06038_);
  and (_06043_, _06042_, _06037_);
  nor (_06044_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_06045_, _06044_, _05925_);
  and (_06046_, _06045_, _05936_);
  and (_06047_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_06048_, _06047_, _06046_);
  and (_06049_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_06050_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_06051_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_06052_, _06051_, _06050_);
  nor (_06053_, _06052_, _06049_);
  and (_06054_, _06053_, _06048_);
  and (_06055_, _06054_, _06043_);
  and (_06056_, _06055_, _06031_);
  and (_06057_, _06056_, _06020_);
  and (_06058_, _06057_, _06003_);
  and (_06059_, _06043_, _06030_);
  and (_06060_, _06059_, _06054_);
  and (_06061_, _06060_, _06020_);
  and (_06062_, _06061_, _06003_);
  or (_06063_, _06062_, _06058_);
  not (_06064_, _06020_);
  and (_06065_, _06060_, _06064_);
  not (_06066_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_06067_, \oc8051_top_1.oc8051_decoder1.wr , _05545_);
  and (_06068_, _06067_, _06066_);
  and (_06069_, _06055_, _06003_);
  nand (_06070_, _06069_, _06068_);
  or (_06071_, _06070_, _06065_);
  or (_06072_, _06071_, _06063_);
  and (_06073_, _06072_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  not (_06074_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  not (_06075_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_06076_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _06075_);
  or (_06077_, _06076_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_06078_, _06077_, _06074_);
  not (_06079_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  not (_06080_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_06081_, _06080_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_06082_, _06081_, _06075_);
  or (_06083_, _06082_, _06079_);
  and (_06084_, _06083_, _06078_);
  not (_06085_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_06086_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_06087_, _06086_, _06080_);
  or (_06088_, _06087_, _06085_);
  or (_06089_, _06076_, _06080_);
  not (_06090_, _06089_);
  nand (_06091_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_06092_, _06091_, _06088_);
  and (_06093_, _06092_, _06084_);
  nor (_06094_, _06086_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_06095_, _06094_);
  not (_06096_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_06097_, _06096_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_06098_, _06097_, ABINPUT[6]);
  nand (_06099_, _06096_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_06100_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_06101_, _06100_, _06098_);
  or (_06102_, _06101_, _06095_);
  not (_06103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_06104_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_06105_, _06104_, _06080_);
  or (_06106_, _06105_, _06103_);
  and (_06107_, _06104_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06108_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_06109_, _06108_, _06106_);
  and (_06110_, _06109_, _06102_);
  nand (_06111_, _06110_, _06093_);
  and (_06112_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05545_);
  and (_06113_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05545_);
  nor (_06114_, _06113_, _06112_);
  and (_06115_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _05545_);
  and (_06116_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _05545_);
  nor (_06117_, _06116_, _06115_);
  and (_06118_, _06117_, _06114_);
  not (_06119_, _06118_);
  and (_06120_, _06115_, _06114_);
  not (_06121_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not (_06122_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_06123_, _06113_, _06122_);
  and (_06124_, _06123_, _06121_);
  nor (_06125_, _06124_, _06120_);
  and (_06126_, _06125_, _06119_);
  and (_06127_, _06112_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06128_, _06127_, _06121_);
  not (_06129_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06130_, _06112_, _06129_);
  and (_06131_, _06130_, _06116_);
  nor (_06132_, _06131_, _06128_);
  and (_06133_, _06132_, _06126_);
  not (_06134_, _06133_);
  and (_06135_, _06134_, _06111_);
  and (_06136_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_06137_, _06136_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor (_06138_, _06097_, ABINPUT[0]);
  nor (_06139_, _06099_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_06140_, _06139_, _06138_);
  nor (_06141_, _06140_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_06142_, _06141_, _06137_);
  not (_06143_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  or (_06144_, _06077_, _06143_);
  not (_06145_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  or (_06146_, _06082_, _06145_);
  and (_06147_, _06146_, _06144_);
  not (_06148_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_06149_, _06087_, _06148_);
  nand (_06150_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_06151_, _06150_, _06149_);
  and (_06152_, _06151_, _06147_);
  or (_06153_, _06097_, ABINPUT[5]);
  or (_06154_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_06155_, _06154_, _06153_);
  or (_06156_, _06155_, _06095_);
  not (_06157_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_06158_, _06105_, _06157_);
  nand (_06159_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_06160_, _06159_, _06158_);
  and (_06161_, _06160_, _06156_);
  nand (_06162_, _06161_, _06152_);
  nor (_06163_, _06162_, _06142_);
  not (_06164_, _06162_);
  not (_06165_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  or (_06166_, _06077_, _06165_);
  not (_06167_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  or (_06168_, _06082_, _06167_);
  and (_06169_, _06168_, _06166_);
  not (_06170_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_06171_, _06087_, _06170_);
  nand (_06172_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_06173_, _06172_, _06171_);
  and (_06174_, _06173_, _06169_);
  or (_06175_, _06097_, ABINPUT[4]);
  or (_06176_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_06177_, _06176_, _06175_);
  or (_06178_, _06177_, _06095_);
  not (_06179_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_06180_, _06105_, _06179_);
  nand (_06181_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_06182_, _06181_, _06180_);
  and (_06183_, _06182_, _06178_);
  nand (_06184_, _06183_, _06174_);
  not (_06185_, _06184_);
  not (_06186_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  nor (_06187_, _06077_, _06186_);
  not (_06188_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  nor (_06189_, _06082_, _06188_);
  nor (_06190_, _06189_, _06187_);
  and (_06191_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_06192_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_06193_, _06087_, _06192_);
  nor (_06194_, _06193_, _06191_);
  and (_06195_, _06194_, _06190_);
  or (_06196_, _06097_, ABINPUT[1]);
  or (_06197_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_06198_, _06197_, _06196_);
  and (_06199_, _06198_, _06094_);
  and (_06200_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not (_06201_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_06202_, _06105_, _06201_);
  nor (_06203_, _06202_, _06200_);
  not (_06204_, _06203_);
  nor (_06205_, _06204_, _06199_);
  and (_06206_, _06205_, _06195_);
  not (_06207_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  or (_06208_, _06082_, _06207_);
  not (_06209_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  or (_06210_, _06077_, _06209_);
  and (_06211_, _06210_, _06208_);
  nand (_06212_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not (_06213_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_06214_, _06105_, _06213_);
  and (_06215_, _06214_, _06212_);
  and (_06216_, _06215_, _06211_);
  not (_06217_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_06218_, _06089_, _06217_);
  not (_06219_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_06220_, _06087_, _06219_);
  and (_06221_, _06220_, _06218_);
  or (_06222_, _06097_, ABINPUT[3]);
  or (_06223_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_06224_, _06223_, _06222_);
  or (_06225_, _06224_, _06095_);
  and (_06226_, _06225_, _06221_);
  nand (_06227_, _06226_, _06216_);
  not (_06228_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  or (_06229_, _06077_, _06228_);
  not (_06230_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  or (_06231_, _06082_, _06230_);
  and (_06232_, _06231_, _06229_);
  not (_06233_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_06234_, _06089_, _06233_);
  not (_06235_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_06236_, _06087_, _06235_);
  and (_06237_, _06236_, _06234_);
  and (_06238_, _06237_, _06232_);
  or (_06239_, _06097_, ABINPUT[2]);
  or (_06240_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_06241_, _06240_, _06239_);
  or (_06242_, _06241_, _06095_);
  not (_06243_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_06244_, _06105_, _06243_);
  nand (_06245_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_06246_, _06245_, _06244_);
  and (_06247_, _06246_, _06242_);
  nand (_06248_, _06247_, _06238_);
  nor (_06249_, _06248_, _06227_);
  and (_06250_, _06249_, _06206_);
  and (_06251_, _06250_, _06185_);
  and (_06252_, _06251_, _06164_);
  not (_06253_, _06142_);
  not (_06254_, _06248_);
  nor (_06255_, _06206_, _06254_);
  and (_06256_, _06255_, _06227_);
  and (_06257_, _06256_, _06184_);
  and (_06258_, _06257_, _06253_);
  nor (_06259_, _06258_, _06252_);
  nor (_06260_, _06259_, _06163_);
  and (_06261_, _06260_, _06111_);
  nor (_06262_, _06260_, _06111_);
  not (_06263_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06265_, _06116_, _06263_);
  and (_06266_, _06127_, _06265_);
  not (_06267_, _06266_);
  or (_06268_, _06267_, _06262_);
  nor (_06269_, _06268_, _06261_);
  nor (_06270_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not (_06271_, _06270_);
  or (_06272_, _06271_, _06101_);
  nand (_06273_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06274_, _06273_, _06074_);
  not (_06275_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_06276_, _06275_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06277_, _06276_, _06103_);
  and (_06278_, _06277_, _06274_);
  nand (_06279_, _06278_, _06272_);
  nor (_06280_, _06279_, _06111_);
  and (_06281_, _06115_, _06121_);
  and (_06282_, _06130_, _06281_);
  not (_06283_, _06282_);
  nor (_06284_, _06283_, _06280_);
  not (_06285_, _06284_);
  and (_06286_, _06279_, _06111_);
  and (_06287_, _06116_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06288_, _06287_, _06123_);
  and (_06289_, _06288_, _06286_);
  and (_06290_, _06265_, _06123_);
  not (_06291_, _06290_);
  nor (_06292_, _06291_, _06111_);
  nor (_06293_, _06292_, _06289_);
  nand (_06294_, _06293_, _06285_);
  and (_06295_, _06127_, _06287_);
  and (_06296_, _06279_, _06142_);
  and (_06297_, _06253_, _06111_);
  or (_06298_, _06297_, _06296_);
  and (_06299_, _06298_, _06295_);
  and (_06300_, _06130_, _06117_);
  nor (_06301_, _06286_, _06280_);
  and (_06302_, _06301_, _06300_);
  or (_06303_, _06302_, _06299_);
  or (_06304_, _06303_, _06294_);
  or (_06305_, _06304_, _06269_);
  nor (_06306_, _06305_, _06135_);
  not (_06307_, _06306_);
  and (_06308_, _06056_, _06064_);
  and (_06309_, _06308_, _06003_);
  and (_06310_, _06309_, _06068_);
  and (_06311_, _06310_, _06307_);
  or (_06312_, _06311_, _06073_);
  and (_10361_, _06312_, _05552_);
  not (_06313_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_06314_, _06123_, _06117_);
  and (_06315_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_06316_, _06315_, _06313_);
  and (_06317_, _06315_, _06313_);
  or (_06318_, _06317_, _06316_);
  and (_10695_, _06318_, _05552_);
  not (_06319_, _05586_);
  nor (_06320_, _06319_, _05577_);
  nor (_06321_, _06320_, _05556_);
  or (_06322_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_06323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _05556_);
  or (_06324_, _06323_, _05586_);
  and (_06325_, _06324_, _05552_);
  and (_11021_, _06325_, _06322_);
  nor (_06326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_11823_, _06326_, rst);
  nor (_06327_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_06328_, _06327_);
  and (_06329_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  not (_06330_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_06331_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _06330_);
  not (_06332_, _06331_);
  or (_06333_, _06271_, _06177_);
  or (_06334_, _06273_, _06165_);
  or (_06335_, _06276_, _06179_);
  and (_06336_, _06335_, _06334_);
  and (_06337_, _06336_, _06333_);
  or (_06339_, _06337_, _06332_);
  and (_06340_, _06278_, _06272_);
  not (_06341_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_06342_, _06341_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_06343_, _06342_);
  or (_06344_, _06343_, _06340_);
  and (_06345_, _06344_, _06339_);
  or (_06346_, _06342_, _06331_);
  or (_06347_, _06271_, _06241_);
  or (_06348_, _06273_, _06228_);
  or (_06349_, _06276_, _06243_);
  and (_06350_, _06349_, _06348_);
  and (_06351_, _06350_, _06347_);
  or (_06352_, _06351_, _06346_);
  and (_06353_, _06352_, _06328_);
  and (_06354_, _06353_, _06345_);
  or (_06355_, _06097_, ABINPUT[8]);
  or (_06356_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_06357_, _06356_, _06355_);
  or (_06358_, _06357_, _06271_);
  not (_06359_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or (_06360_, _06273_, _06359_);
  not (_06361_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_06362_, _06276_, _06361_);
  and (_06363_, _06362_, _06360_);
  and (_06364_, _06363_, _06358_);
  and (_06365_, _06364_, _06327_);
  nor (_06366_, _06365_, _06354_);
  and (_06367_, _06366_, _06248_);
  not (_06368_, _06206_);
  or (_06369_, _06271_, _06224_);
  or (_06370_, _06273_, _06209_);
  or (_06371_, _06276_, _06213_);
  and (_06372_, _06371_, _06370_);
  and (_06373_, _06372_, _06369_);
  or (_06374_, _06373_, _06332_);
  or (_06375_, _06271_, _06155_);
  or (_06376_, _06273_, _06143_);
  or (_06377_, _06276_, _06157_);
  and (_06378_, _06377_, _06376_);
  and (_06379_, _06378_, _06375_);
  or (_06380_, _06379_, _06343_);
  and (_06381_, _06380_, _06374_);
  nand (_06382_, _06270_, _06198_);
  or (_06383_, _06273_, _06186_);
  or (_06384_, _06276_, _06201_);
  and (_06385_, _06384_, _06383_);
  and (_06386_, _06385_, _06382_);
  or (_06387_, _06386_, _06346_);
  and (_06388_, _06387_, _06328_);
  nand (_06389_, _06388_, _06381_);
  or (_06390_, _06097_, ABINPUT[7]);
  or (_06391_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_06392_, _06391_, _06390_);
  or (_06393_, _06392_, _06271_);
  not (_06394_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  or (_06395_, _06273_, _06394_);
  not (_06396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_06397_, _06276_, _06396_);
  and (_06398_, _06397_, _06395_);
  nand (_06399_, _06398_, _06393_);
  or (_06400_, _06399_, _06328_);
  and (_06401_, _06400_, _06389_);
  and (_06402_, _06401_, _06368_);
  and (_06403_, _06402_, _06367_);
  and (_06404_, _06401_, _06227_);
  nand (_06405_, _06404_, _06367_);
  or (_06406_, _06404_, _06367_);
  and (_06407_, _06406_, _06405_);
  and (_06408_, _06407_, _06403_);
  and (_06409_, _06401_, _06184_);
  nand (_06410_, _06400_, _06389_);
  or (_06411_, _06410_, _06254_);
  and (_06412_, _06366_, _06227_);
  and (_06413_, _06412_, _06411_);
  nand (_06414_, _06413_, _06409_);
  or (_06415_, _06413_, _06409_);
  and (_06416_, _06415_, _06414_);
  nand (_06417_, _06416_, _06408_);
  not (_06418_, _06417_);
  nand (_06419_, _06414_, _06405_);
  or (_06420_, _06365_, _06354_);
  or (_06421_, _06420_, _06185_);
  or (_06422_, _06410_, _06164_);
  or (_06423_, _06422_, _06421_);
  nand (_06424_, _06422_, _06421_);
  and (_06425_, _06424_, _06423_);
  nand (_06426_, _06425_, _06419_);
  or (_06427_, _06425_, _06419_);
  and (_06428_, _06427_, _06426_);
  and (_06429_, _06428_, _06418_);
  and (_06430_, _06425_, _06419_);
  and (_06431_, _06366_, _06162_);
  and (_06432_, _06431_, _06409_);
  not (_06433_, _06111_);
  or (_06434_, _06420_, _06433_);
  or (_06435_, _06434_, _06422_);
  and (_06436_, _06401_, _06111_);
  or (_06437_, _06436_, _06431_);
  and (_06438_, _06437_, _06435_);
  nand (_06439_, _06438_, _06432_);
  or (_06440_, _06438_, _06432_);
  and (_06441_, _06440_, _06439_);
  nand (_06442_, _06441_, _06430_);
  or (_06443_, _06441_, _06430_);
  and (_06444_, _06443_, _06442_);
  nand (_06445_, _06444_, _06429_);
  or (_06446_, _06444_, _06429_);
  and (_06447_, _06446_, _06445_);
  and (_06448_, _06447_, _06329_);
  nor (_06449_, _06447_, _06329_);
  or (_06450_, _06449_, _06448_);
  and (_06451_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_06452_, _06416_, _06408_);
  and (_06453_, _06452_, _06417_);
  nand (_06454_, _06453_, _06451_);
  and (_06455_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  not (_06456_, _06455_);
  nor (_06457_, _06407_, _06403_);
  or (_06458_, _06457_, _06408_);
  or (_06459_, _06458_, _06456_);
  or (_06461_, _06453_, _06451_);
  nand (_06462_, _06461_, _06454_);
  or (_06463_, _06462_, _06459_);
  nand (_06464_, _06463_, _06454_);
  and (_06465_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nand (_06466_, _06428_, _06418_);
  or (_06467_, _06428_, _06418_);
  and (_06469_, _06467_, _06466_);
  nand (_06470_, _06469_, _06465_);
  or (_06471_, _06469_, _06465_);
  and (_06472_, _06471_, _06470_);
  nand (_06473_, _06472_, _06464_);
  or (_06474_, _06473_, _06450_);
  not (_06475_, _06470_);
  nor (_06476_, _06475_, _06448_);
  or (_06477_, _06476_, _06449_);
  and (_06478_, _06477_, _06474_);
  and (_06479_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  not (_06480_, _06445_);
  not (_06481_, _06434_);
  not (_06482_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  or (_06483_, _06082_, _06482_);
  or (_06485_, _06077_, _06394_);
  and (_06486_, _06485_, _06483_);
  not (_06487_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_06488_, _06087_, _06487_);
  not (_06489_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_06490_, _06089_, _06489_);
  and (_06491_, _06490_, _06488_);
  and (_06492_, _06491_, _06486_);
  or (_06493_, _06392_, _06095_);
  or (_06494_, _06105_, _06396_);
  nand (_06495_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_06496_, _06495_, _06494_);
  and (_06497_, _06496_, _06493_);
  and (_06498_, _06497_, _06492_);
  or (_06499_, _06498_, _06435_);
  not (_06500_, _06498_);
  and (_06501_, _06500_, _06401_);
  not (_06502_, _06501_);
  nand (_06503_, _06502_, _06435_);
  and (_06504_, _06503_, _06499_);
  nand (_06505_, _06504_, _06481_);
  or (_06506_, _06501_, _06481_);
  nand (_06507_, _06506_, _06505_);
  and (_06508_, _06442_, _06439_);
  nand (_06509_, _06508_, _06507_);
  or (_06510_, _06508_, _06507_);
  and (_06511_, _06510_, _06509_);
  nand (_06512_, _06511_, _06480_);
  or (_06513_, _06511_, _06480_);
  and (_06514_, _06513_, _06512_);
  nand (_06515_, _06514_, _06479_);
  or (_06516_, _06514_, _06479_);
  nand (_06517_, _06516_, _06515_);
  or (_06518_, _06517_, _06478_);
  not (_06519_, _06518_);
  and (_06520_, _06517_, _06478_);
  nor (_06521_, _06520_, _06519_);
  and (_12386_, _06521_, _05552_);
  and (_06522_, _05934_, _05933_);
  not (_06523_, _06522_);
  and (_06524_, _06523_, _06068_);
  and (_06525_, _06524_, _06020_);
  and (_06526_, _06525_, _06060_);
  not (_06527_, _05989_);
  and (_06528_, _06001_, _06527_);
  nor (_06529_, _05971_, _05958_);
  and (_06530_, _06529_, _06528_);
  and (_06531_, _06530_, _06526_);
  not (_06532_, _06531_);
  and (_06533_, _06532_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_06534_, _06336_, _06333_);
  and (_06535_, _06534_, _06295_);
  and (_06536_, _06256_, _06253_);
  and (_06537_, _06250_, _06142_);
  nor (_06538_, _06537_, _06536_);
  nor (_06539_, _06538_, _06185_);
  and (_06540_, _06538_, _06185_);
  or (_06541_, _06540_, _06267_);
  nor (_06542_, _06541_, _06539_);
  nor (_06543_, _06542_, _06535_);
  nor (_06544_, _06534_, _06184_);
  nor (_06545_, _06544_, _06283_);
  not (_06546_, _06300_);
  and (_06547_, _06534_, _06184_);
  or (_06549_, _06547_, _06544_);
  nor (_06550_, _06549_, _06546_);
  or (_06551_, _06550_, _06545_);
  not (_06552_, _06551_);
  and (_06553_, _06547_, _06288_);
  nor (_06554_, _06291_, _06184_);
  nor (_06555_, _06554_, _06553_);
  and (_06556_, _06184_, _06134_);
  not (_06557_, _06556_);
  and (_06558_, _06557_, _06555_);
  and (_06559_, _06558_, _06552_);
  and (_06560_, _06559_, _06543_);
  nor (_06561_, _06560_, _06532_);
  nor (_06562_, _06561_, _06533_);
  nor (_13222_, _06562_, rst);
  or (_06563_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not (_06564_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_06565_, _05550_, _06564_);
  and (_06566_, _06565_, _05552_);
  and (_01193_, _06566_, _06563_);
  and (_06567_, _05822_, _05669_);
  and (_06568_, _06567_, _05839_);
  and (_06569_, _05837_, _05812_);
  and (_06570_, _06569_, _05738_);
  not (_06571_, _06570_);
  nor (_06572_, _05850_, _05822_);
  nor (_06573_, _06572_, _06571_);
  nor (_06574_, _06573_, _06568_);
  not (_06575_, _06574_);
  and (_06576_, _05547_, _05552_);
  nand (_01436_, _06576_, _06575_);
  or (_06577_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_06578_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _05556_);
  or (_06579_, _06578_, _05586_);
  and (_06580_, _06579_, _05552_);
  and (_01904_, _06580_, _06577_);
  and (_06581_, _06265_, _06114_);
  not (_06582_, _06581_);
  not (_06583_, _06364_);
  not (_06584_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  or (_06585_, _06082_, _06584_);
  or (_06586_, _06077_, _06359_);
  and (_06587_, _06586_, _06585_);
  not (_06588_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_06589_, _06089_, _06588_);
  not (_06590_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_06591_, _06087_, _06590_);
  and (_06593_, _06591_, _06589_);
  and (_06594_, _06593_, _06587_);
  or (_06595_, _06357_, _06095_);
  or (_06596_, _06105_, _06361_);
  nand (_06597_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_06598_, _06597_, _06596_);
  and (_06599_, _06598_, _06595_);
  and (_06600_, _06599_, _06594_);
  and (_06601_, _06600_, _06583_);
  and (_06602_, _06600_, _06364_);
  nor (_06603_, _06600_, _06364_);
  nor (_06604_, _06603_, _06602_);
  nor (_06605_, _06498_, _06399_);
  not (_06606_, _06399_);
  nor (_06608_, _06498_, _06606_);
  and (_06609_, _06498_, _06606_);
  nor (_06611_, _06609_, _06608_);
  and (_06612_, _06340_, _06111_);
  nor (_06613_, _06379_, _06162_);
  nor (_06614_, _06613_, _06301_);
  nor (_06615_, _06614_, _06612_);
  nor (_06616_, _06615_, _06611_);
  nor (_06617_, _06616_, _06605_);
  and (_06618_, _06615_, _06611_);
  nor (_06619_, _06618_, _06616_);
  not (_06620_, _06619_);
  and (_06621_, _06613_, _06301_);
  nor (_06622_, _06621_, _06614_);
  not (_06624_, _06622_);
  nand (_06625_, _06378_, _06375_);
  and (_06626_, _06625_, _06162_);
  nor (_06627_, _06625_, _06162_);
  nor (_06628_, _06627_, _06626_);
  not (_06629_, _06628_);
  not (_06630_, _06549_);
  nand (_06631_, _06372_, _06369_);
  and (_06632_, _06631_, _06227_);
  nor (_06633_, _06631_, _06227_);
  nor (_06634_, _06633_, _06632_);
  nand (_06635_, _06350_, _06347_);
  and (_06636_, _06635_, _06248_);
  nor (_06637_, _06635_, _06248_);
  nor (_06638_, _06637_, _06636_);
  nand (_06639_, _06385_, _06382_);
  and (_06640_, _06639_, _06206_);
  nor (_06641_, _06640_, _06638_);
  and (_06642_, _06351_, _06248_);
  nor (_06643_, _06642_, _06641_);
  nor (_06644_, _06643_, _06634_);
  and (_06645_, _06373_, _06227_);
  nor (_06646_, _06645_, _06644_);
  nor (_06647_, _06646_, _06630_);
  and (_06648_, _06646_, _06630_);
  nor (_06649_, _06648_, _06647_);
  and (_06650_, _06643_, _06634_);
  nor (_06651_, _06650_, _06644_);
  not (_06652_, _06651_);
  and (_06653_, _06640_, _06638_);
  nor (_06654_, _06653_, _06641_);
  not (_06655_, _06654_);
  nor (_06656_, _06386_, _06206_);
  and (_06657_, _06386_, _06206_);
  nor (_06658_, _06657_, _06656_);
  nor (_06659_, _06658_, _06253_);
  and (_06660_, _06659_, _06655_);
  and (_06661_, _06660_, _06652_);
  not (_06662_, _06661_);
  nor (_06663_, _06662_, _06649_);
  nand (_06664_, _06337_, _06184_);
  nor (_06665_, _06337_, _06184_);
  or (_06666_, _06646_, _06665_);
  and (_06667_, _06666_, _06664_);
  or (_06668_, _06667_, _06663_);
  and (_06669_, _06668_, _06629_);
  and (_06670_, _06669_, _06624_);
  and (_06671_, _06670_, _06620_);
  nor (_06672_, _06671_, _06617_);
  nor (_06673_, _06672_, _06604_);
  nor (_06674_, _06673_, _06601_);
  nor (_06675_, _06674_, _06582_);
  not (_06676_, _06675_);
  and (_06677_, _06281_, _06114_);
  not (_06678_, _06677_);
  not (_06679_, _06603_);
  not (_06680_, _06634_);
  and (_06681_, _06656_, _06638_);
  nor (_06682_, _06681_, _06636_);
  nor (_06683_, _06682_, _06680_);
  nor (_06684_, _06683_, _06632_);
  nor (_06685_, _06684_, _06630_);
  and (_06686_, _06684_, _06630_);
  nor (_06687_, _06686_, _06685_);
  and (_06688_, _06658_, _06142_);
  and (_06689_, _06688_, _06638_);
  and (_06690_, _06682_, _06680_);
  nor (_06692_, _06690_, _06683_);
  and (_06693_, _06692_, _06689_);
  not (_06694_, _06693_);
  nor (_06695_, _06694_, _06687_);
  nor (_06696_, _06684_, _06544_);
  or (_06697_, _06696_, _06547_);
  or (_06698_, _06697_, _06695_);
  and (_06699_, _06698_, _06628_);
  and (_06700_, _06699_, _06301_);
  not (_06701_, _06611_);
  and (_06702_, _06626_, _06301_);
  nor (_06703_, _06702_, _06286_);
  nor (_06704_, _06703_, _06701_);
  and (_06705_, _06703_, _06701_);
  nor (_06706_, _06705_, _06704_);
  and (_06707_, _06706_, _06700_);
  not (_06708_, _06707_);
  nor (_06709_, _06704_, _06608_);
  and (_06710_, _06709_, _06708_);
  or (_06711_, _06710_, _06602_);
  and (_06712_, _06711_, _06679_);
  nor (_06713_, _06712_, _06678_);
  nor (_06714_, _06500_, _06111_);
  not (_06715_, _06714_);
  and (_06716_, _06281_, _06123_);
  nor (_06717_, _06249_, _06185_);
  and (_06718_, _06717_, _06716_);
  and (_06719_, _06718_, _06162_);
  nor (_06720_, _06719_, _06715_);
  nor (_06721_, _06720_, _06600_);
  nor (_06722_, _06721_, _06142_);
  not (_06723_, _06722_);
  not (_06724_, _06716_);
  nor (_06725_, _06600_, _06253_);
  not (_06726_, _06725_);
  nor (_06727_, _06726_, _06720_);
  nor (_06728_, _06727_, _06724_);
  and (_06729_, _06728_, _06723_);
  not (_06730_, _06718_);
  and (_06731_, _06140_, _06137_);
  and (_06732_, _06130_, _06265_);
  and (_06733_, _06288_, _06140_);
  nor (_06734_, _06733_, _06732_);
  nor (_06735_, _06734_, _06731_);
  and (_06736_, _06127_, _06281_);
  and (_06737_, _06368_, _06736_);
  nor (_06738_, _06737_, _06735_);
  nor (_06739_, _06142_, _06140_);
  not (_06740_, _06140_);
  nor (_06741_, _06740_, _06137_);
  nor (_06742_, _06741_, _06546_);
  nor (_06743_, _06742_, _06282_);
  nor (_06744_, _06743_, _06739_);
  not (_06745_, _06744_);
  and (_06746_, _06130_, _06287_);
  not (_06747_, _06600_);
  and (_06748_, _06747_, _06746_);
  or (_06749_, _06290_, _06142_);
  and (_06750_, _06127_, _06117_);
  and (_06751_, _06740_, _06750_);
  nor (_06752_, _06751_, _06118_);
  nand (_06753_, _06752_, _06142_);
  and (_06754_, _06753_, _06749_);
  nor (_06755_, _06754_, _06748_);
  and (_06756_, _06755_, _06745_);
  and (_06757_, _06756_, _06738_);
  and (_06758_, _06757_, _06730_);
  not (_06759_, _06758_);
  nor (_06760_, _06759_, _06729_);
  not (_06761_, _06760_);
  nor (_06762_, _06761_, _06713_);
  and (_06763_, _06762_, _06676_);
  not (_06764_, _06001_);
  and (_06765_, _06764_, _05958_);
  nor (_06766_, _06527_, _05971_);
  and (_06767_, _06766_, _06020_);
  and (_06768_, _06767_, _06765_);
  not (_06769_, _06054_);
  nor (_06770_, _06043_, _06030_);
  and (_06771_, _06770_, _06769_);
  and (_06772_, _06771_, _06768_);
  nand (_06773_, _06772_, _06763_);
  and (_06774_, _06523_, _06067_);
  and (_06775_, _06774_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or (_06776_, _06772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_06777_, _06776_, _06775_);
  and (_06778_, _06777_, _06773_);
  and (_06779_, _06766_, _06765_);
  and (_06781_, _06779_, _06061_);
  not (_06782_, _06781_);
  and (_06783_, _06600_, _06253_);
  not (_06784_, _06783_);
  not (_06785_, _06295_);
  and (_06786_, _06364_, _06142_);
  nor (_06787_, _06786_, _06785_);
  and (_06788_, _06787_, _06784_);
  and (_06789_, _06714_, _06252_);
  nor (_06790_, _06789_, _06253_);
  and (_06791_, _06162_, _06111_);
  and (_06792_, _06791_, _06257_);
  and (_06793_, _06792_, _06500_);
  nor (_06794_, _06793_, _06142_);
  or (_06795_, _06794_, _06790_);
  and (_06796_, _06795_, _06600_);
  nor (_06797_, _06795_, _06600_);
  nor (_06798_, _06797_, _06796_);
  and (_06799_, _06798_, _06266_);
  nor (_06800_, _06799_, _06788_);
  nor (_06801_, _06602_, _06283_);
  and (_06802_, _06604_, _06300_);
  nor (_06803_, _06802_, _06801_);
  and (_06804_, _06603_, _06288_);
  and (_06805_, _06600_, _06290_);
  nor (_06806_, _06805_, _06804_);
  nor (_06807_, _06600_, _06133_);
  not (_06808_, _06807_);
  and (_06809_, _06808_, _06806_);
  and (_06810_, _06809_, _06803_);
  and (_06811_, _06810_, _06800_);
  nor (_06812_, _06811_, _06782_);
  and (_06813_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_06814_, _06813_, _06812_);
  and (_06815_, _06814_, _06524_);
  not (_06816_, _06774_);
  and (_06817_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_06818_, _06817_, rst);
  or (_06819_, _06818_, _06815_);
  or (_02004_, _06819_, _06778_);
  or (_06820_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_06821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _05556_);
  or (_06822_, _06821_, _05586_);
  and (_06823_, _06822_, _05552_);
  and (_02117_, _06823_, _06820_);
  or (_06824_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_06825_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _05556_);
  or (_06826_, _06825_, _05586_);
  and (_06827_, _06826_, _05552_);
  and (_02328_, _06827_, _06824_);
  and (_06828_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and (_06829_, _06747_, _06366_);
  and (_06830_, _06829_, _06502_);
  or (_06831_, _06600_, _06410_);
  or (_06832_, _06498_, _06420_);
  or (_06833_, _06832_, _06831_);
  nand (_06834_, _06832_, _06831_);
  and (_06835_, _06834_, _06833_);
  not (_06836_, _06835_);
  or (_06837_, _06836_, _06505_);
  or (_06838_, _06836_, _06499_);
  and (_06839_, _06838_, _06837_);
  not (_06840_, _06839_);
  nand (_06841_, _06840_, _06830_);
  or (_06842_, _06840_, _06830_);
  and (_06843_, _06842_, _06841_);
  nor (_06844_, _06507_, _06439_);
  nand (_06845_, _06836_, _06505_);
  nand (_06846_, _06845_, _06837_);
  nand (_06847_, _06846_, _06499_);
  and (_06848_, _06847_, _06838_);
  nand (_06849_, _06848_, _06844_);
  or (_06850_, _06848_, _06844_);
  and (_06851_, _06850_, _06849_);
  or (_06852_, _06507_, _06442_);
  nand (_06853_, _06852_, _06512_);
  nand (_06854_, _06853_, _06851_);
  nand (_06855_, _06854_, _06849_);
  nand (_06856_, _06855_, _06843_);
  and (_06857_, _06841_, _06833_);
  nand (_06858_, _06857_, _06856_);
  nand (_06859_, _06858_, _06828_);
  or (_06860_, _06858_, _06828_);
  nand (_06861_, _06860_, _06859_);
  and (_06862_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or (_06863_, _06855_, _06843_);
  and (_06864_, _06863_, _06856_);
  nand (_06865_, _06864_, _06862_);
  or (_06866_, _06865_, _06861_);
  nand (_06867_, _06866_, _06859_);
  and (_06868_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_06869_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_06870_, _06869_, _06868_);
  and (_06871_, _06870_, _06867_);
  and (_06872_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or (_06873_, _06853_, _06851_);
  and (_06874_, _06873_, _06854_);
  nand (_06875_, _06874_, _06872_);
  or (_06876_, _06874_, _06872_);
  nand (_06877_, _06876_, _06875_);
  and (_06878_, _06518_, _06515_);
  or (_06879_, _06878_, _06877_);
  and (_06880_, _06879_, _06875_);
  or (_06881_, _06864_, _06862_);
  nand (_06882_, _06881_, _06865_);
  nor (_06883_, _06882_, _06861_);
  nand (_06884_, _06870_, _06883_);
  nor (_06885_, _06884_, _06880_);
  nor (_06886_, _06885_, _06871_);
  or (_06887_, _06882_, _06880_);
  and (_06888_, _06887_, _06865_);
  or (_06889_, _06888_, _06861_);
  nand (_06890_, _06889_, _06859_);
  nand (_06891_, _06890_, _06868_);
  not (_06892_, _06869_);
  nand (_06893_, _06892_, _06891_);
  and (_06895_, _06893_, _06886_);
  and (_03645_, _06895_, _05552_);
  or (_06896_, _06885_, _06871_);
  and (_06897_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_06898_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_06899_, _06898_, _06897_);
  nand (_06901_, _06899_, _06896_);
  nand (_06902_, _06897_, _06896_);
  not (_06903_, _06898_);
  nand (_06904_, _06903_, _06902_);
  and (_06905_, _06904_, _06901_);
  and (_03742_, _06905_, _05552_);
  or (_06906_, _06897_, _06896_);
  and (_06908_, _06906_, _06902_);
  and (_04571_, _06908_, _05552_);
  and (_06910_, _06001_, _05958_);
  not (_06911_, _05971_);
  and (_06913_, _06020_, _06527_);
  and (_06915_, _06913_, _06911_);
  and (_06916_, _06915_, _06910_);
  and (_06918_, _06916_, _06771_);
  nand (_06919_, _06918_, _06763_);
  or (_06921_, _06918_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_06922_, _06921_, _06775_);
  and (_06924_, _06922_, _06919_);
  not (_06925_, _05958_);
  nor (_06926_, _05971_, _06925_);
  and (_06927_, _06926_, _06528_);
  and (_06928_, _06927_, _06061_);
  nand (_06929_, _06928_, _06811_);
  or (_06930_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_06931_, _06930_, _06524_);
  and (_06932_, _06931_, _06929_);
  and (_06933_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_06934_, _06933_, rst);
  or (_06935_, _06934_, _06932_);
  or (_05142_, _06935_, _06924_);
  or (_06936_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_06937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _05556_);
  or (_06938_, _06937_, _05586_);
  and (_06939_, _06938_, _05552_);
  and (_05539_, _06939_, _06936_);
  or (_06940_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_06941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _05556_);
  or (_06942_, _06941_, _05586_);
  and (_06943_, _06942_, _05552_);
  and (_05540_, _06943_, _06940_);
  or (_06944_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_06945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _05556_);
  or (_06946_, _06945_, _05586_);
  and (_06947_, _06946_, _05552_);
  and (_05541_, _06947_, _06944_);
  and (_06948_, _06065_, _06003_);
  and (_06949_, _06948_, _06068_);
  nand (_06950_, _06949_, _06306_);
  or (_06951_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_06952_, _06951_, _05552_);
  and (_05578_, _06952_, _06950_);
  not (_06953_, _06058_);
  nor (_06954_, _06560_, _06953_);
  not (_06955_, _06068_);
  and (_06956_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_06957_, _06956_, _06955_);
  or (_06958_, _06957_, _06954_);
  or (_06959_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_06960_, _06959_, _05552_);
  and (_05581_, _06960_, _06958_);
  not (_06962_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_06963_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05545_);
  and (_06965_, _06963_, _06962_);
  not (_06966_, _06965_);
  not (_06967_, _06524_);
  and (_06968_, _06764_, _05989_);
  and (_06969_, _06968_, _06529_);
  nand (_06970_, _06969_, _06061_);
  or (_06971_, _06970_, _06967_);
  and (_06972_, _06971_, _06966_);
  not (_06973_, _06972_);
  or (_06974_, _06639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_06975_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_06976_, _06631_, _06975_);
  and (_06977_, _06976_, _06974_);
  or (_06978_, _06977_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_06979_, _06625_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_06980_, _06399_, _06975_);
  and (_06981_, _06980_, _06979_);
  or (_06982_, _06981_, _06313_);
  nand (_06983_, _06982_, _06978_);
  and (_06984_, _06982_, _06978_);
  nor (_06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_06986_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_06987_, _06986_);
  nand (_06988_, _06985_, _06600_);
  and (_06989_, _06988_, _06987_);
  not (_06990_, _06989_);
  or (_06991_, _06990_, _06984_);
  nor (_06992_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_06993_, _06992_);
  nand (_06994_, _06985_, _06498_);
  and (_06995_, _06994_, _06993_);
  not (_06996_, _06995_);
  and (_06997_, _06635_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_06998_, _06997_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_06999_, _06534_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07000_, _06279_, _06975_);
  and (_07001_, _07000_, _06999_);
  or (_07002_, _07001_, _06313_);
  and (_07003_, _07002_, _06998_);
  or (_07004_, _07003_, _06996_);
  or (_07005_, _06989_, _06983_);
  and (_07006_, _07005_, _06991_);
  not (_07007_, _07006_);
  or (_07008_, _07007_, _07004_);
  and (_07009_, _07008_, _06991_);
  nand (_07010_, _07002_, _06998_);
  or (_07011_, _07010_, _06995_);
  and (_07012_, _07011_, _07004_);
  and (_07013_, _07012_, _07006_);
  not (_07014_, _06985_);
  or (_07015_, _07014_, _06111_);
  nor (_07016_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_07017_, _07016_);
  nand (_07018_, _07017_, _07015_);
  and (_07019_, _06639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07020_, _07019_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07021_, _06631_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07022_, _06625_, _06975_);
  and (_07023_, _07022_, _07021_);
  or (_07024_, _07023_, _06313_);
  and (_07025_, _07024_, _07020_);
  or (_07026_, _07025_, _07018_);
  or (_07027_, _06635_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07028_, _06534_, _06975_);
  and (_07029_, _07028_, _07027_);
  and (_07030_, _07029_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07031_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_07032_, _07031_);
  or (_07033_, _07014_, _06162_);
  nand (_07034_, _07033_, _07032_);
  or (_07035_, _07034_, _07030_);
  and (_07036_, _07017_, _07015_);
  nand (_07037_, _07024_, _07020_);
  or (_07038_, _07037_, _07036_);
  nand (_07039_, _07038_, _07026_);
  or (_07040_, _07039_, _07035_);
  nand (_07041_, _07040_, _07026_);
  nand (_07042_, _07041_, _07013_);
  and (_07043_, _07042_, _07009_);
  and (_07044_, _06977_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07045_, _07044_);
  nor (_07046_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_07047_, _07046_);
  or (_07048_, _07014_, _06184_);
  and (_07049_, _07048_, _07047_);
  nand (_07050_, _07049_, _07045_);
  or (_07051_, _07049_, _07045_);
  nand (_07052_, _07051_, _07050_);
  nand (_07053_, _06997_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07054_, _07014_, _06227_);
  nor (_07055_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_07056_, _07055_);
  and (_07057_, _07056_, _07054_);
  nand (_07058_, _07057_, _07053_);
  and (_07059_, _07019_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07060_, _07014_, _06248_);
  nor (_07061_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_07062_, _07061_);
  nand (_07063_, _07062_, _07060_);
  and (_07064_, _07063_, _07059_);
  or (_07065_, _07057_, _07053_);
  nand (_07066_, _07065_, _07058_);
  or (_07067_, _07066_, _07064_);
  and (_07068_, _07067_, _07058_);
  or (_07069_, _07068_, _07052_);
  nand (_07070_, _07069_, _07050_);
  nand (_07071_, _07034_, _07030_);
  and (_07072_, _07071_, _07035_);
  and (_07073_, _07038_, _07026_);
  and (_07074_, _07073_, _07072_);
  and (_07075_, _07074_, _07013_);
  nand (_07076_, _07075_, _07070_);
  nand (_07077_, _07076_, _07043_);
  nor (_07078_, _07029_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07079_, _06279_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07081_, _06364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07082_, _07081_, _07079_);
  and (_07084_, _07082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07086_, _07084_, _07078_);
  not (_07087_, _07086_);
  and (_07088_, _06364_, _06606_);
  nor (_07089_, _07088_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_07090_, _07001_, _06981_);
  not (_07091_, _07023_);
  and (_07092_, _07082_, _07091_);
  nand (_07093_, _07092_, _07090_);
  and (_07094_, _07093_, _06313_);
  nor (_07095_, _07094_, _07089_);
  and (_07096_, _07095_, _07087_);
  nand (_07097_, _07096_, _07077_);
  not (_07098_, _07012_);
  and (_07099_, _07025_, _07018_);
  not (_07100_, _07035_);
  and (_07101_, _07072_, _07070_);
  nor (_07102_, _07101_, _07100_);
  or (_07103_, _07102_, _07099_);
  and (_07104_, _07103_, _07026_);
  nor (_07105_, _07104_, _07098_);
  and (_07106_, _07104_, _07098_);
  nor (_07108_, _07106_, _07105_);
  nor (_07110_, _07108_, _07097_);
  and (_07111_, _07097_, _06996_);
  nor (_07112_, _07111_, _07110_);
  and (_07114_, _07112_, _06983_);
  nor (_07115_, _07112_, _06983_);
  nor (_07116_, _07115_, _07114_);
  and (_07117_, _07096_, _07077_);
  nand (_07118_, _07039_, _07102_);
  or (_07119_, _07039_, _07102_);
  nand (_07120_, _07119_, _07118_);
  nand (_07121_, _07120_, _07117_);
  and (_07122_, _07097_, _07018_);
  not (_07123_, _07122_);
  and (_07124_, _07123_, _07121_);
  and (_07125_, _07124_, _07010_);
  nor (_07126_, _07072_, _07070_);
  or (_07127_, _07126_, _07101_);
  and (_07128_, _07127_, _07117_);
  and (_07129_, _07097_, _07034_);
  nor (_07130_, _07129_, _07128_);
  and (_07131_, _07130_, _07037_);
  not (_07132_, _07131_);
  nor (_07133_, _07124_, _07010_);
  or (_07134_, _07133_, _07125_);
  nor (_07135_, _07134_, _07132_);
  nor (_07136_, _07135_, _07125_);
  not (_07137_, _07030_);
  and (_07138_, _07068_, _07052_);
  not (_07140_, _07138_);
  and (_07141_, _07140_, _07069_);
  or (_07142_, _07141_, _07097_);
  or (_07143_, _07117_, _07049_);
  and (_07144_, _07143_, _07142_);
  nor (_07145_, _07144_, _07137_);
  not (_07146_, _07145_);
  not (_07147_, _07059_);
  or (_07148_, _07097_, _07147_);
  nand (_07149_, _07148_, _07063_);
  or (_07150_, _07148_, _07063_);
  and (_07151_, _07150_, _07149_);
  nand (_07152_, _07151_, _07053_);
  or (_07153_, _07151_, _07053_);
  and (_07154_, _07153_, _07152_);
  and (_07155_, _06985_, _06206_);
  nor (_07156_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_07157_, _07156_, _07155_);
  nor (_07158_, _07157_, _07147_);
  not (_07159_, _07158_);
  nand (_07160_, _07159_, _07154_);
  and (_07161_, _07160_, _07152_);
  or (_07162_, _07117_, _07057_);
  and (_07163_, _07066_, _07064_);
  not (_07164_, _07163_);
  and (_07165_, _07164_, _07067_);
  or (_07166_, _07165_, _07097_);
  and (_07167_, _07166_, _07162_);
  nand (_07168_, _07167_, _07045_);
  or (_07169_, _07167_, _07045_);
  nand (_07170_, _07169_, _07168_);
  or (_07171_, _07170_, _07161_);
  and (_07172_, _07144_, _07137_);
  not (_07173_, _07172_);
  and (_07174_, _07173_, _07168_);
  nand (_07175_, _07174_, _07171_);
  and (_07176_, _07175_, _07146_);
  nor (_07177_, _07130_, _07037_);
  nor (_07178_, _07177_, _07131_);
  not (_07179_, _07178_);
  nor (_07181_, _07134_, _07179_);
  nand (_07182_, _07181_, _07176_);
  nand (_07183_, _07182_, _07136_);
  nand (_07184_, _07183_, _07116_);
  not (_07185_, _07114_);
  and (_07186_, _07097_, _06989_);
  not (_07187_, _07105_);
  and (_07188_, _07187_, _07004_);
  nand (_07189_, _07188_, _07006_);
  or (_07190_, _07188_, _07006_);
  nand (_07191_, _07190_, _07189_);
  and (_07192_, _07191_, _07117_);
  nor (_07193_, _07192_, _07186_);
  or (_07194_, _07193_, _07086_);
  and (_07195_, _07194_, _07185_);
  nand (_07196_, _07195_, _07184_);
  and (_07197_, _07193_, _07086_);
  not (_07198_, _07197_);
  and (_07199_, _07198_, _07095_);
  and (_07200_, _07199_, _07196_);
  and (_07201_, _07198_, _07194_);
  nand (_07202_, _07184_, _07185_);
  or (_07203_, _07202_, _07201_);
  nand (_07204_, _07202_, _07201_);
  and (_07205_, _07204_, _07203_);
  nand (_07206_, _07205_, _07200_);
  or (_07208_, _07200_, _07193_);
  nand (_07209_, _07208_, _07206_);
  nand (_07210_, _07209_, _06314_);
  and (_07211_, _06287_, _06114_);
  and (_07212_, _06899_, _06896_);
  and (_07213_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  nand (_07214_, _07213_, _07212_);
  and (_07215_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_07216_, _07215_, _07214_);
  or (_07217_, _07214_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_07218_, _07217_, _07216_);
  nand (_07219_, _07218_, _07211_);
  not (_07220_, _06604_);
  and (_07221_, _06672_, _07220_);
  nor (_07222_, _06672_, _07220_);
  nor (_07224_, _07222_, _07221_);
  and (_07225_, _07224_, _06581_);
  not (_07226_, _07225_);
  nor (_07227_, _06710_, _06604_);
  and (_07228_, _06710_, _06604_);
  or (_07229_, _07228_, _07227_);
  and (_07230_, _07229_, _06677_);
  nor (_07231_, _06714_, _06600_);
  nor (_07232_, _07231_, _06142_);
  and (_07233_, _07232_, _06730_);
  nor (_07234_, _07233_, _06720_);
  and (_07235_, _07234_, _06600_);
  nor (_07236_, _07234_, _06600_);
  nor (_07237_, _07236_, _07235_);
  nor (_07238_, _07237_, _06724_);
  and (_07239_, _06368_, _06750_);
  and (_07240_, _06142_, _06736_);
  nor (_07241_, _07240_, _07239_);
  nor (_07242_, _06600_, _06119_);
  and (_07243_, _06500_, _06131_);
  nor (_07244_, _07243_, _07242_);
  and (_07245_, _07244_, _07241_);
  and (_07246_, _07245_, _06806_);
  and (_07247_, _07246_, _06803_);
  not (_07248_, _07247_);
  nor (_07249_, _07248_, _07238_);
  and (_07250_, _07249_, _06800_);
  not (_07251_, _07250_);
  nor (_07252_, _07251_, _07230_);
  and (_07253_, _07252_, _07226_);
  and (_07254_, _07253_, _07219_);
  nand (_07255_, _07254_, _07210_);
  nand (_07257_, _07255_, _06973_);
  not (_07258_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_07259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05545_);
  and (_07260_, _07259_, _07258_);
  not (_07261_, _07260_);
  nor (_07262_, _06001_, _05958_);
  and (_07263_, _07262_, _06775_);
  and (_07264_, _07263_, _06767_);
  and (_07265_, _07264_, _06771_);
  and (_07266_, _07265_, _06763_);
  and (_07267_, _07262_, _06767_);
  and (_07269_, _07267_, _06775_);
  and (_07270_, _07269_, _06771_);
  nor (_07271_, _07270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_07272_, _07271_, _06973_);
  or (_07273_, _07272_, _07266_);
  and (_07274_, _07273_, _07261_);
  nand (_07275_, _07274_, _07257_);
  nor (_07276_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07277_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06085_);
  nor (_07278_, _07277_, _07276_);
  nor (_07279_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07280_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06170_);
  nor (_07281_, _07280_, _07279_);
  nor (_07282_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07283_, _06192_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07284_, _07283_, _07282_);
  not (_07285_, _07284_);
  nor (_07286_, _07285_, _06712_);
  nor (_07288_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_07289_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06235_);
  nor (_07290_, _07289_, _07288_);
  and (_07291_, _07290_, _07286_);
  nor (_07292_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_07293_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06219_);
  nor (_07294_, _07293_, _07292_);
  and (_07295_, _07294_, _07291_);
  and (_07296_, _07295_, _07281_);
  nor (_07297_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07298_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06148_);
  nor (_07299_, _07298_, _07297_);
  and (_07300_, _07299_, _07296_);
  and (_07301_, _07300_, _07278_);
  nor (_07302_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07303_, _06487_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07304_, _07303_, _07302_);
  and (_07305_, _07304_, _07301_);
  nor (_07306_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_07308_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06590_);
  nor (_07309_, _07308_, _07306_);
  or (_07310_, _07309_, _07305_);
  nand (_07311_, _07309_, _07305_);
  and (_07312_, _07311_, _07310_);
  nand (_07313_, _07312_, _06677_);
  and (_07314_, _06878_, _06877_);
  not (_07315_, _07314_);
  and (_07316_, _07315_, _06879_);
  and (_07317_, _07316_, _07211_);
  nor (_07318_, _06600_, _06386_);
  and (_07319_, _07318_, _06793_);
  and (_07320_, _07319_, _06635_);
  and (_07321_, _07320_, _06631_);
  and (_07322_, _07321_, _06534_);
  and (_07323_, _07322_, _06625_);
  nor (_07325_, _07323_, _06142_);
  and (_07326_, _06789_, _06600_);
  and (_07327_, _06351_, _06386_);
  and (_07328_, _06337_, _06373_);
  and (_07329_, _07328_, _07327_);
  and (_07330_, _07329_, _07326_);
  and (_07331_, _07330_, _06379_);
  nor (_07332_, _07331_, _06253_);
  nor (_07333_, _07332_, _07325_);
  nor (_07334_, _06279_, _06142_);
  nor (_07335_, _07334_, _06296_);
  and (_07336_, _07335_, _07333_);
  nor (_07337_, _06399_, _06142_);
  and (_07339_, _06399_, _06142_);
  nor (_07340_, _07339_, _07337_);
  and (_07342_, _07340_, _07336_);
  and (_07343_, _07342_, _06583_);
  nor (_07344_, _07342_, _06583_);
  nor (_07345_, _07344_, _07343_);
  and (_07346_, _07345_, _06266_);
  and (_07347_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_07348_, _06785_, _06142_);
  or (_07349_, _07348_, _06118_);
  and (_07350_, _07349_, _06583_);
  or (_07351_, _07350_, _07347_);
  and (_07352_, _06184_, _06746_);
  and (_07353_, _06725_, _06295_);
  or (_07354_, _07353_, _07352_);
  nor (_07355_, _07354_, _07351_);
  not (_07356_, _07355_);
  nor (_07357_, _07356_, _07346_);
  not (_07358_, _07357_);
  nor (_07359_, _07358_, _07317_);
  nand (_07360_, _07359_, _07313_);
  or (_07362_, _07360_, _07261_);
  and (_07363_, _07362_, _07275_);
  and (_05610_, _07363_, _05552_);
  and (_07364_, _06532_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_07365_, _06251_, _06142_);
  nor (_07366_, _07365_, _06258_);
  and (_07367_, _07366_, _06164_);
  nor (_07368_, _07366_, _06164_);
  nor (_07369_, _07368_, _07367_);
  and (_07370_, _07369_, _06266_);
  and (_07371_, _06379_, _06142_);
  nor (_07372_, _07371_, _06785_);
  not (_07373_, _07372_);
  nor (_07374_, _07373_, _06163_);
  nor (_07375_, _07374_, _07370_);
  and (_07376_, _06162_, _06134_);
  not (_07377_, _07376_);
  and (_07378_, _06628_, _06300_);
  not (_07379_, _07378_);
  nor (_07380_, _06627_, _06283_);
  not (_07381_, _07380_);
  and (_07382_, _06626_, _06288_);
  nor (_07383_, _06291_, _06162_);
  nor (_07384_, _07383_, _07382_);
  and (_07385_, _07384_, _07381_);
  and (_07386_, _07385_, _07379_);
  and (_07387_, _07386_, _07377_);
  and (_07388_, _07387_, _07375_);
  nor (_07389_, _07388_, _06532_);
  nor (_07390_, _07389_, _07364_);
  not (_07391_, _07390_);
  and (_07392_, _06562_, _05669_);
  and (_07393_, _07392_, _07391_);
  and (_07394_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_07395_, _06562_, _05818_);
  and (_07396_, _07395_, _07391_);
  and (_07397_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_07398_, _07397_, _07394_);
  nor (_07399_, _06562_, _05818_);
  and (_07400_, _07399_, _07391_);
  and (_07401_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor (_07402_, _06562_, _05669_);
  and (_07403_, _07402_, _07391_);
  and (_07404_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_07405_, _07404_, _07401_);
  and (_07406_, _07405_, _07398_);
  and (_07407_, _07395_, _07390_);
  and (_07408_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_07410_, _07392_, _07390_);
  and (_07411_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_07412_, _07411_, _07408_);
  and (_07413_, _07399_, _07390_);
  and (_07414_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_07416_, _07402_, _07390_);
  and (_07417_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_07418_, _07417_, _07414_);
  and (_07419_, _07418_, _07412_);
  and (_07420_, _07419_, _07406_);
  nor (_07421_, _07390_, _06527_);
  and (_07422_, _07390_, _06527_);
  nor (_07423_, _07422_, _07421_);
  and (_07424_, _06562_, _06064_);
  nor (_07425_, _06059_, _05669_);
  not (_07426_, _07425_);
  and (_07427_, _06068_, _06054_);
  and (_07428_, _07427_, _06001_);
  and (_07429_, _07428_, _05972_);
  nand (_07430_, _07429_, _07426_);
  nor (_07431_, _07430_, _07424_);
  nor (_07432_, _06562_, _06064_);
  and (_07433_, _06043_, _06031_);
  nor (_07434_, _07433_, _05818_);
  nor (_07435_, _07434_, _07432_);
  and (_07436_, _07435_, _07431_);
  and (_07437_, _07436_, _07423_);
  nor (_07438_, _07437_, _07420_);
  not (_07439_, _06811_);
  and (_07440_, _07437_, _07439_);
  nor (_07441_, _07440_, _07438_);
  nor (_05672_, _07441_, rst);
  and (_07442_, _06525_, _06054_);
  and (_07443_, _06910_, _06766_);
  and (_07444_, _07443_, _07442_);
  and (_07445_, _07444_, _06770_);
  nand (_07446_, _07199_, _07196_);
  or (_07447_, _07172_, _07145_);
  and (_07448_, _07171_, _07168_);
  nor (_07449_, _07448_, _07447_);
  and (_07450_, _07448_, _07447_);
  nor (_07451_, _07450_, _07449_);
  or (_07452_, _07451_, _07446_);
  or (_07453_, _07200_, _07144_);
  and (_07454_, _07453_, _07452_);
  nand (_07455_, _07454_, _06314_);
  nand (_07456_, _06895_, _07211_);
  and (_07457_, _06694_, _06687_);
  or (_07458_, _07457_, _06678_);
  nor (_07459_, _07458_, _06695_);
  not (_07460_, _07459_);
  and (_07461_, _06662_, _06649_);
  nor (_07462_, _07461_, _06663_);
  nor (_07463_, _07462_, _06582_);
  and (_07464_, _06184_, _06118_);
  and (_07465_, _06227_, _06131_);
  nor (_07466_, _07465_, _07464_);
  nor (_07467_, _06717_, _06724_);
  not (_07468_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_07469_, _06249_, _07468_);
  or (_07470_, _07469_, _06184_);
  nand (_07471_, _07470_, _07467_);
  nand (_07472_, _06162_, _06128_);
  and (_07473_, _07472_, _06555_);
  and (_07474_, _07473_, _07471_);
  and (_07475_, _07474_, _07466_);
  and (_07476_, _07475_, _06543_);
  and (_07477_, _07476_, _06552_);
  not (_07478_, _07477_);
  nor (_07479_, _07478_, _07463_);
  and (_07481_, _07479_, _07460_);
  and (_07482_, _07481_, _07456_);
  nand (_07483_, _07482_, _07455_);
  and (_07484_, _07483_, _07445_);
  and (_07485_, _07259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_07486_, _07445_);
  and (_07487_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_07488_, _07487_, _07485_);
  or (_07489_, _07488_, _07484_);
  and (_07490_, _06534_, _06118_);
  nor (_07491_, _07321_, _06142_);
  and (_07492_, _07327_, _07326_);
  and (_07493_, _07492_, _06373_);
  nor (_07494_, _07493_, _06253_);
  or (_07495_, _07494_, _07491_);
  and (_07496_, _07495_, _06337_);
  nor (_07497_, _07495_, _06337_);
  nor (_07498_, _07497_, _07496_);
  and (_07499_, _07498_, _06266_);
  and (_07500_, _06295_, _06184_);
  or (_07501_, _07500_, _07499_);
  or (_07503_, _07501_, _06748_);
  and (_07504_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_07505_, _07295_, _07281_);
  nor (_07506_, _07505_, _07296_);
  and (_07507_, _07506_, _06677_);
  and (_07508_, _06462_, _06459_);
  not (_07509_, _07508_);
  and (_07510_, _07509_, _06463_);
  and (_07511_, _07510_, _07211_);
  or (_07512_, _07511_, _07507_);
  or (_07513_, _07512_, _07504_);
  or (_07514_, _07513_, _07503_);
  nor (_07515_, _07514_, _07490_);
  nand (_07516_, _07515_, _07485_);
  and (_07517_, _07516_, _05552_);
  and (_05863_, _07517_, _07489_);
  or (_07518_, _07183_, _07116_);
  nand (_07519_, _07518_, _07184_);
  nand (_07520_, _07519_, _07200_);
  or (_07521_, _07200_, _07112_);
  and (_07522_, _07521_, _07520_);
  nand (_07523_, _07522_, _06314_);
  or (_07524_, _07213_, _07212_);
  and (_07525_, _07524_, _07214_);
  nand (_07526_, _07525_, _07211_);
  nor (_07527_, _06670_, _06620_);
  nor (_07528_, _07527_, _06671_);
  nor (_07529_, _07528_, _06582_);
  not (_07530_, _07529_);
  nor (_07531_, _06706_, _06700_);
  nor (_07532_, _07531_, _06678_);
  and (_07533_, _07532_, _06708_);
  nor (_07534_, _06498_, _06142_);
  or (_07535_, _07534_, _07339_);
  and (_07536_, _07535_, _06295_);
  or (_07537_, _06792_, _06500_);
  and (_07538_, _07537_, _06794_);
  and (_07539_, _06252_, _06433_);
  nor (_07540_, _06498_, _07539_);
  or (_07542_, _07540_, _06789_);
  and (_07543_, _07542_, _06142_);
  or (_07544_, _07543_, _07538_);
  and (_07545_, _07544_, _06266_);
  nor (_07546_, _07545_, _07536_);
  nor (_07547_, _07233_, _06719_);
  and (_07548_, _07547_, _06433_);
  and (_07549_, _07548_, _06498_);
  nor (_07550_, _07548_, _06498_);
  nor (_07551_, _07550_, _07549_);
  nor (_07552_, _07551_, _06724_);
  and (_07553_, _06611_, _06300_);
  and (_07554_, _06608_, _06288_);
  nor (_07555_, _06609_, _06283_);
  and (_07556_, _06498_, _06290_);
  or (_07557_, _07556_, _07555_);
  or (_07558_, _07557_, _07554_);
  nor (_07559_, _07558_, _07553_);
  not (_07560_, _06128_);
  or (_07561_, _06600_, _07560_);
  and (_07562_, _06131_, _06111_);
  nor (_07563_, _06498_, _06119_);
  nor (_07564_, _07563_, _07562_);
  and (_07565_, _07564_, _07561_);
  and (_07566_, _07565_, _07559_);
  not (_07567_, _07566_);
  nor (_07568_, _07567_, _07552_);
  and (_07569_, _07568_, _07546_);
  not (_07570_, _07569_);
  nor (_07571_, _07570_, _07533_);
  and (_07572_, _07571_, _07530_);
  and (_07573_, _07572_, _07526_);
  nand (_07574_, _07573_, _07523_);
  and (_07575_, _07574_, _07445_);
  and (_07576_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_07577_, _07576_, _07485_);
  or (_07578_, _07577_, _07575_);
  not (_07579_, _07485_);
  and (_07580_, _06399_, _06118_);
  and (_07581_, _06227_, _06746_);
  and (_07582_, _07336_, _06606_);
  nor (_07583_, _07336_, _06606_);
  or (_07584_, _07583_, _07582_);
  and (_07585_, _07584_, _06266_);
  and (_07586_, _06498_, _06142_);
  not (_07587_, _07586_);
  nor (_07588_, _07337_, _06785_);
  and (_07589_, _07588_, _07587_);
  or (_07590_, _07589_, _07585_);
  or (_07591_, _07590_, _07581_);
  and (_07592_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_07593_, _07304_, _07301_);
  nor (_07594_, _07593_, _07305_);
  and (_07595_, _07594_, _06677_);
  and (_07596_, _06521_, _07211_);
  or (_07597_, _07596_, _07595_);
  or (_07598_, _07597_, _07592_);
  or (_07599_, _07598_, _07591_);
  or (_07600_, _07599_, _07580_);
  or (_07601_, _07600_, _07579_);
  and (_07602_, _07601_, _05552_);
  and (_05866_, _07602_, _07578_);
  nand (_07603_, _07178_, _07176_);
  and (_07604_, _07603_, _07132_);
  nand (_07605_, _07134_, _07604_);
  or (_07606_, _07134_, _07604_);
  and (_07607_, _07606_, _07605_);
  or (_07608_, _07607_, _07446_);
  or (_07609_, _07200_, _07124_);
  and (_07610_, _07609_, _07608_);
  and (_07611_, _07610_, _06314_);
  and (_07612_, _06905_, _07211_);
  nor (_07613_, _06669_, _06624_);
  nor (_07614_, _07613_, _06670_);
  nor (_07616_, _07614_, _06582_);
  nor (_07617_, _06626_, _06301_);
  nor (_07618_, _07617_, _06702_);
  or (_07619_, _07618_, _06699_);
  nor (_07620_, _06700_, _06678_);
  and (_07621_, _07620_, _07619_);
  nor (_07622_, _07547_, _06433_);
  or (_07623_, _07622_, _07548_);
  and (_07624_, _07623_, _06716_);
  and (_07625_, _06118_, _06111_);
  and (_07626_, _06162_, _06131_);
  nor (_07627_, _06498_, _07560_);
  or (_07628_, _07627_, _07626_);
  or (_07629_, _07628_, _07625_);
  or (_07630_, _07629_, _07624_);
  or (_07631_, _07630_, _06305_);
  or (_07632_, _07631_, _07621_);
  or (_07633_, _07632_, _07616_);
  or (_07634_, _07633_, _07612_);
  or (_07635_, _07634_, _07611_);
  and (_07636_, _07635_, _07445_);
  and (_07637_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_07638_, _07637_, _07485_);
  or (_07639_, _07638_, _07636_);
  or (_07640_, _07300_, _07278_);
  nor (_07641_, _07301_, _06678_);
  and (_07642_, _07641_, _07640_);
  and (_07643_, _06473_, _06470_);
  nand (_07644_, _07643_, _06450_);
  or (_07645_, _07643_, _06450_);
  and (_07646_, _07645_, _07644_);
  and (_07647_, _07646_, _07211_);
  nand (_07648_, _07333_, _06279_);
  or (_07649_, _07333_, _06279_);
  and (_07650_, _07649_, _06266_);
  and (_07651_, _07650_, _07648_);
  and (_07652_, _06248_, _06746_);
  or (_07653_, _06253_, _06111_);
  nor (_07654_, _07334_, _06785_);
  and (_07655_, _07654_, _07653_);
  and (_07656_, _06279_, _06118_);
  and (_07657_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_07658_, _07657_, _07656_);
  or (_07659_, _07658_, _07655_);
  or (_07660_, _07659_, _07652_);
  or (_07661_, _07660_, _07651_);
  or (_07662_, _07661_, _07647_);
  or (_07663_, _07662_, _07642_);
  or (_07664_, _07663_, _07579_);
  and (_07665_, _07664_, _05552_);
  and (_05871_, _07665_, _07639_);
  nor (_07666_, _06043_, _06031_);
  and (_07667_, _07444_, _07666_);
  nor (_07668_, _07667_, _07485_);
  or (_07669_, _07668_, _07483_);
  not (_07670_, _07668_);
  or (_07671_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_07672_, _07671_, _05552_);
  and (_05899_, _07672_, _07669_);
  nand (_07674_, _07200_, _07059_);
  and (_07675_, _07674_, _07157_);
  nor (_07676_, _07674_, _07157_);
  or (_07677_, _07676_, _07675_);
  nand (_07678_, _07677_, _06314_);
  nor (_07679_, _06658_, _06142_);
  nor (_07680_, _07679_, _06688_);
  nor (_07681_, _06677_, _06581_);
  not (_07682_, _07681_);
  and (_07683_, _07682_, _07680_);
  not (_07684_, _07683_);
  and (_07685_, _06656_, _06288_);
  and (_07686_, _06290_, _06206_);
  nor (_07687_, _07686_, _07685_);
  and (_07688_, _06639_, _06295_);
  and (_07689_, _06266_, _06206_);
  nor (_07690_, _07689_, _07688_);
  and (_07691_, _06747_, _06732_);
  and (_07692_, _06142_, _06746_);
  nor (_07693_, _07692_, _07691_);
  and (_07694_, _07693_, _07690_);
  and (_07695_, _07694_, _07687_);
  not (_07696_, _06887_);
  and (_07697_, _06882_, _06880_);
  nor (_07698_, _07697_, _07696_);
  and (_07699_, _07698_, _07211_);
  nor (_07700_, _06656_, _06546_);
  nor (_07701_, _07700_, _06282_);
  or (_07702_, _07701_, _06657_);
  and (_07703_, _06248_, _06128_);
  nor (_07704_, _06716_, _06118_);
  nor (_07705_, _07704_, _06206_);
  nor (_07706_, _07705_, _07703_);
  nand (_07707_, _07706_, _07702_);
  nor (_07708_, _07707_, _07699_);
  and (_07709_, _07708_, _07695_);
  and (_07710_, _07709_, _07684_);
  nand (_07711_, _07710_, _07678_);
  or (_07712_, _07711_, _07668_);
  or (_07713_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_07714_, _07713_, _05552_);
  and (_05929_, _07714_, _07712_);
  or (_07715_, _07668_, _07574_);
  or (_07716_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_07717_, _07716_, _05552_);
  and (_05932_, _07717_, _07715_);
  and (_06005_, _06402_, _05552_);
  or (_07718_, _06472_, _06464_);
  and (_07719_, _07718_, _06473_);
  and (_06007_, _07719_, _05552_);
  and (_06013_, _07510_, _05552_);
  and (_07720_, _06458_, _06456_);
  not (_07721_, _07720_);
  and (_07722_, _07721_, _06459_);
  and (_06017_, _07722_, _05552_);
  and (_07723_, _06366_, _06368_);
  not (_07724_, _07723_);
  and (_07725_, _07724_, _06411_);
  nor (_07726_, _07725_, _06403_);
  and (_06036_, _07726_, _05552_);
  and (_07727_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_07728_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05552_);
  and (_07729_, _07728_, _05917_);
  or (_06264_, _07729_, _07727_);
  nor (_07730_, _05575_, _05562_);
  or (_07731_, _07730_, _05556_);
  and (_07732_, _07731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_07733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_07734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_07735_, _07734_, _07733_);
  and (_07736_, _05562_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_07737_, _07736_, _07735_);
  or (_07738_, _07737_, _07732_);
  and (_06338_, _07738_, _05552_);
  and (_07740_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_06460_, _07740_, _05558_);
  nor (_07741_, _05547_, _06584_);
  and (_07742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_07743_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_07744_, _05616_, _07743_);
  nor (_07745_, _05624_, _05768_);
  or (_07746_, _07745_, _07744_);
  and (_07747_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_07748_, _05631_, _05762_);
  or (_07749_, _07748_, _07747_);
  or (_07750_, _07749_, _07746_);
  and (_07751_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_07752_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_07753_, _07752_, _07751_);
  or (_07754_, _07753_, _07750_);
  and (_07755_, _07754_, _05671_);
  or (_07756_, _07755_, _07742_);
  and (_07757_, _07756_, _05547_);
  nor (_07758_, _07757_, _07741_);
  nor (_06468_, _07758_, rst);
  and (_07759_, _05777_, _05729_);
  and (_07760_, _05799_, _05752_);
  and (_07761_, _07760_, _07759_);
  nor (_07762_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_07763_, _07762_, _05608_);
  and (_07764_, _07763_, _05706_);
  and (_07765_, _05660_, _05636_);
  and (_07766_, _07765_, _07764_);
  and (_07767_, _07766_, _05685_);
  and (_06484_, _07767_, _07761_);
  and (_06548_, _07316_, _05552_);
  not (_07768_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_07769_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07768_);
  and (_07770_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_07771_, _07770_, _07769_);
  and (_06592_, _07771_, _05552_);
  nor (_07772_, _05710_, _05689_);
  not (_07773_, _05665_);
  nor (_07774_, _07773_, _05641_);
  and (_07775_, _07774_, _07772_);
  not (_07776_, _05781_);
  and (_07777_, _05803_, _07776_);
  and (_07778_, _05756_, _05733_);
  and (_07779_, _07778_, _07777_);
  and (_07780_, _07779_, _07775_);
  not (_07781_, _05756_);
  and (_07782_, _07781_, _05733_);
  nor (_07783_, _05803_, _05781_);
  and (_07784_, _07783_, _07782_);
  and (_07785_, _07784_, _07775_);
  nor (_07786_, _07785_, _07780_);
  not (_07787_, _05803_);
  and (_07788_, _07787_, _05781_);
  and (_07789_, _05689_, _05641_);
  nor (_07790_, _05733_, _05710_);
  and (_07791_, _07790_, _07789_);
  and (_07792_, _07791_, _07788_);
  not (_07793_, _07792_);
  nor (_07794_, _07781_, _05733_);
  and (_07795_, _07794_, _07788_);
  and (_07796_, _07795_, _05710_);
  nor (_07797_, _05665_, _05641_);
  and (_07798_, _07797_, _07772_);
  nor (_07799_, _07798_, _07796_);
  and (_07800_, _07799_, _07793_);
  and (_07801_, _07800_, _07786_);
  nor (_07802_, _05710_, _07773_);
  not (_07803_, _05689_);
  nor (_07804_, _07803_, _05641_);
  and (_07805_, _07804_, _07802_);
  not (_07806_, _07805_);
  and (_07807_, _07782_, _07777_);
  not (_07808_, _07807_);
  and (_07809_, _07788_, _07778_);
  and (_07810_, _07783_, _07781_);
  nor (_07811_, _07810_, _07809_);
  and (_07812_, _07811_, _07808_);
  nor (_07813_, _07812_, _07806_);
  not (_07814_, _05710_);
  and (_07815_, _07804_, _07814_);
  and (_07816_, _07815_, _07773_);
  not (_07817_, _07816_);
  nor (_07818_, _05756_, _05733_);
  and (_07819_, _05803_, _05781_);
  and (_07820_, _07819_, _07818_);
  and (_07821_, _07783_, _05756_);
  nor (_07823_, _07821_, _07820_);
  nor (_07824_, _07823_, _07817_);
  nor (_07825_, _07824_, _07813_);
  and (_07826_, _07825_, _07801_);
  and (_07827_, _07819_, _07782_);
  and (_07828_, _07827_, _07816_);
  not (_07830_, _07828_);
  and (_07831_, _07803_, _05641_);
  nor (_07832_, _07831_, _07804_);
  not (_07833_, _07832_);
  and (_07834_, _07777_, _07781_);
  and (_07835_, _07834_, _07790_);
  and (_07836_, _07835_, _07833_);
  and (_07837_, _07816_, _07810_);
  nor (_07838_, _07837_, _07836_);
  and (_07839_, _07838_, _07830_);
  and (_07840_, _07795_, _07775_);
  and (_07841_, _05733_, _07814_);
  and (_07842_, _07841_, _07789_);
  nor (_07843_, _05803_, _05756_);
  and (_07844_, _07843_, _05781_);
  or (_07845_, _07834_, _07844_);
  and (_07846_, _07845_, _07842_);
  nor (_07847_, _07846_, _07840_);
  and (_07848_, _07788_, _07782_);
  and (_07849_, _07848_, _07775_);
  not (_07850_, _07775_);
  and (_07851_, _07794_, _07777_);
  nor (_07852_, _07851_, _07834_);
  nor (_07853_, _07852_, _07850_);
  nor (_07854_, _07853_, _07849_);
  and (_07855_, _07854_, _07847_);
  and (_07856_, _07855_, _07839_);
  and (_07857_, _07856_, _07826_);
  nor (_07859_, _07794_, _07782_);
  and (_07860_, _07859_, _07783_);
  and (_07861_, _07860_, _07775_);
  and (_07862_, _07819_, _07778_);
  and (_07863_, _07862_, _07816_);
  nor (_07864_, _07863_, _07861_);
  and (_07865_, _07831_, _07802_);
  and (_07866_, _07865_, _07821_);
  not (_07867_, _07866_);
  or (_07868_, _07807_, _07795_);
  and (_07869_, _07868_, _07816_);
  and (_07870_, _07848_, _07805_);
  nor (_07871_, _07870_, _07869_);
  and (_07872_, _07871_, _07867_);
  and (_07873_, _07872_, _07864_);
  not (_07874_, _07865_);
  and (_07875_, _07819_, _07794_);
  nor (_07876_, _07875_, _07848_);
  nor (_07877_, _07876_, _07874_);
  and (_07878_, _05803_, _05756_);
  and (_07879_, _07878_, _05781_);
  and (_07880_, _07818_, _07788_);
  nor (_07881_, _07880_, _07879_);
  nor (_07882_, _07881_, _07850_);
  nor (_07883_, _07882_, _07877_);
  nor (_07884_, _07875_, _07809_);
  nor (_07885_, _07884_, _07817_);
  nor (_07886_, _07862_, _07807_);
  nor (_07887_, _07886_, _07874_);
  nor (_07888_, _07887_, _07885_);
  and (_07889_, _07888_, _07883_);
  and (_07890_, _07889_, _07873_);
  and (_07891_, _07890_, _07857_);
  and (_07892_, _07833_, _07802_);
  nor (_07893_, _07892_, _07816_);
  not (_07894_, _07893_);
  and (_07895_, _07894_, _07851_);
  not (_07896_, _07895_);
  and (_07897_, _07831_, _07814_);
  and (_07898_, _07897_, _07773_);
  and (_07899_, _07851_, _07898_);
  and (_07900_, _07809_, _07775_);
  nor (_07901_, _07900_, _07899_);
  not (_07902_, _07901_);
  and (_07903_, _07848_, _07816_);
  and (_07904_, _07898_, _07779_);
  or (_07905_, _07904_, _07903_);
  nor (_07906_, _07905_, _07902_);
  and (_07907_, _07906_, _07896_);
  and (_07908_, _07865_, _07788_);
  and (_07909_, _07908_, _07859_);
  and (_07910_, _07908_, _07794_);
  nor (_07911_, _07910_, _07909_);
  not (_07912_, _07844_);
  and (_07913_, _07886_, _07912_);
  nor (_07914_, _07913_, _07814_);
  and (_07915_, _07894_, _07779_);
  nor (_07916_, _07915_, _07914_);
  and (_07917_, _07916_, _07911_);
  and (_07918_, _07917_, _07907_);
  and (_07919_, _07918_, _07891_);
  and (_07920_, _07818_, _07777_);
  and (_07921_, _07920_, _07898_);
  or (_07922_, _07789_, _05710_);
  and (_07923_, _07922_, _07848_);
  or (_07924_, _07923_, _07785_);
  nor (_07925_, _07924_, _07921_);
  nand (_07926_, _07925_, _07901_);
  nor (_07928_, _07926_, _07905_);
  nand (_07929_, _07928_, _07873_);
  nor (_07930_, _07929_, _07919_);
  nor (_07931_, _07930_, _05548_);
  nand (_07932_, _07931_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_07933_, rst, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_07934_, _07931_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07935_, _07934_, _07933_);
  and (_06607_, _07935_, _07932_);
  and (_07936_, _06528_, _05972_);
  and (_07937_, _07936_, _06057_);
  and (_07938_, _07937_, _06068_);
  not (_07939_, _07938_);
  and (_07940_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_07941_, _06206_, _06133_);
  not (_07942_, _07941_);
  and (_07943_, _07942_, _07690_);
  and (_07944_, _07943_, _07687_);
  and (_07945_, _07944_, _07702_);
  nor (_07946_, _07945_, _06955_);
  and (_07947_, _07946_, _07937_);
  or (_07948_, _07947_, _07940_);
  and (_06610_, _07948_, _05552_);
  and (_07949_, _07936_, _06061_);
  and (_07950_, _07949_, _06068_);
  not (_07951_, _07950_);
  and (_07952_, _07951_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_07953_, _06635_, _06295_);
  and (_07954_, _06206_, _06254_);
  nor (_07955_, _06255_, _07954_);
  and (_07956_, _07955_, _06253_);
  nor (_07957_, _07955_, _06253_);
  or (_07958_, _07957_, _07956_);
  and (_07959_, _07958_, _06266_);
  nor (_07960_, _07959_, _07953_);
  nor (_07961_, _06254_, _06133_);
  not (_07962_, _07961_);
  and (_07963_, _06638_, _06300_);
  not (_07964_, _07963_);
  nor (_07965_, _06637_, _06283_);
  not (_07966_, _07965_);
  and (_07967_, _06636_, _06288_);
  nor (_07969_, _06291_, _06248_);
  nor (_07970_, _07969_, _07967_);
  and (_07971_, _07970_, _07966_);
  and (_07972_, _07971_, _07964_);
  and (_07974_, _07972_, _07962_);
  and (_07975_, _07974_, _07960_);
  nor (_07976_, _07975_, _06955_);
  and (_07977_, _07976_, _07949_);
  or (_07978_, _07977_, _07952_);
  and (_06623_, _07978_, _05552_);
  and (_06691_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _05552_);
  and (_06780_, _05781_, _05552_);
  or (_07979_, _06674_, _06672_);
  not (_07980_, _06601_);
  nand (_07981_, _06672_, _07980_);
  and (_07982_, _07981_, _06581_);
  and (_07983_, _07982_, _07979_);
  nand (_07984_, _06710_, _06679_);
  and (_07985_, _06711_, _06677_);
  and (_07986_, _07985_, _07984_);
  and (_07987_, _06379_, _06340_);
  and (_07988_, _07987_, _07088_);
  and (_07989_, _07988_, _07329_);
  nand (_07990_, _07989_, _06314_);
  nand (_07991_, _07990_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_07992_, _07991_, _07986_);
  or (_07993_, _07992_, _07983_);
  nand (_07994_, _06888_, _06861_);
  and (_07995_, _07994_, _06889_);
  or (_07996_, _07995_, _07698_);
  or (_07997_, _06890_, _06868_);
  and (_07998_, _07997_, _06891_);
  or (_07999_, _07998_, _07996_);
  or (_08000_, _07999_, _06895_);
  or (_08001_, _08000_, _06908_);
  or (_08002_, _07525_, _06905_);
  or (_08003_, _08002_, _07218_);
  or (_08004_, _08003_, _08001_);
  and (_08005_, _08004_, _07211_);
  or (_08006_, _08005_, _07993_);
  nor (_08007_, _06764_, _05958_);
  and (_08008_, _08007_, _06775_);
  and (_08009_, _08008_, _06915_);
  nor (_08010_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_08011_, _08010_, _08009_);
  and (_08012_, _08011_, _08006_);
  and (_08013_, _07666_, _06054_);
  not (_08014_, _08013_);
  nor (_08015_, _08014_, _06763_);
  and (_08016_, _08014_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_08017_, _08016_, _08015_);
  and (_08018_, _08017_, _08009_);
  or (_08019_, _08018_, _06531_);
  or (_08020_, _08019_, _08012_);
  nor (_08021_, _06255_, _06142_);
  nor (_08022_, _07954_, _06253_);
  nor (_08023_, _08022_, _08021_);
  nor (_08024_, _08023_, _06227_);
  and (_08025_, _08023_, _06227_);
  nor (_08026_, _08025_, _08024_);
  and (_08027_, _08026_, _06266_);
  and (_08028_, _06631_, _06295_);
  nor (_08029_, _08028_, _08027_);
  and (_08030_, _06632_, _06288_);
  nor (_08031_, _06291_, _06227_);
  nor (_08033_, _08031_, _08030_);
  not (_08034_, _06227_);
  nor (_08035_, _08034_, _06133_);
  and (_08036_, _06634_, _06300_);
  nor (_08037_, _06633_, _06283_);
  or (_08038_, _08037_, _08036_);
  nor (_08039_, _08038_, _08035_);
  and (_08040_, _08039_, _08033_);
  and (_08041_, _08040_, _08029_);
  nand (_08042_, _08041_, _06531_);
  and (_08043_, _08042_, _05552_);
  and (_06894_, _08043_, _08020_);
  not (_08044_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_08045_, _08009_, _06056_);
  nor (_08046_, _08045_, _08044_);
  or (_08047_, _08046_, _06531_);
  not (_08048_, _06763_);
  and (_08049_, _08045_, _08048_);
  or (_08050_, _08049_, _08047_);
  nand (_08051_, _07975_, _06531_);
  and (_08052_, _08051_, _05552_);
  and (_06900_, _08052_, _08050_);
  nor (_06907_, _05665_, rst);
  and (_06909_, _05641_, _05552_);
  and (_06912_, _05689_, _05552_);
  and (_06914_, _05710_, _05552_);
  and (_06917_, _05733_, _05552_);
  nor (_06920_, _05756_, rst);
  and (_06923_, _05803_, _05552_);
  nand (_08053_, _07975_, _06949_);
  or (_08054_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_08055_, _08054_, _08053_);
  and (_06961_, _08055_, _05552_);
  not (_08056_, _08009_);
  and (_08057_, _06059_, _06769_);
  nor (_08058_, _06059_, _06769_);
  nor (_08059_, _08058_, _08057_);
  or (_08060_, _08059_, _08056_);
  and (_08061_, _08060_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_08062_, _08057_, _08048_);
  and (_08063_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_08064_, _08063_, _08062_);
  and (_08065_, _08064_, _08009_);
  or (_08066_, _08065_, _08061_);
  and (_08067_, _08066_, _06532_);
  or (_08068_, _08067_, _07389_);
  and (_06964_, _08068_, _05552_);
  or (_08069_, _07159_, _07154_);
  and (_08070_, _08069_, _07160_);
  or (_08071_, _08070_, _07446_);
  or (_08072_, _07200_, _07151_);
  and (_08073_, _08072_, _08071_);
  nand (_08074_, _08073_, _06314_);
  nand (_08075_, _07995_, _07211_);
  nor (_08076_, _06659_, _06655_);
  nor (_08077_, _08076_, _06660_);
  nor (_08078_, _08077_, _06582_);
  not (_08079_, _08078_);
  nand (_08080_, _06227_, _06128_);
  and (_08081_, _06368_, _06131_);
  and (_08082_, _06248_, _06118_);
  nor (_08083_, _08082_, _08081_);
  and (_08084_, _08083_, _08080_);
  and (_08085_, _08084_, _07972_);
  and (_08086_, _08085_, _07960_);
  nor (_08087_, _06717_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_08088_, _08087_, _06248_);
  nor (_08089_, _08087_, _06248_);
  nor (_08090_, _08089_, _08088_);
  nor (_08091_, _08090_, _06724_);
  nor (_08092_, _06656_, _06638_);
  or (_08093_, _08092_, _06681_);
  and (_08094_, _08093_, _06688_);
  nor (_08095_, _08093_, _06688_);
  or (_08096_, _08095_, _08094_);
  and (_08097_, _08096_, _06677_);
  nor (_08098_, _08097_, _08091_);
  and (_08099_, _08098_, _08086_);
  and (_08100_, _08099_, _08079_);
  and (_08101_, _08100_, _08075_);
  nand (_08102_, _08101_, _08074_);
  or (_08103_, _08102_, _07668_);
  or (_08104_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_08105_, _08104_, _05552_);
  and (_07080_, _08105_, _08103_);
  and (_08106_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_08107_, _08106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_07083_, _08107_, _05552_);
  and (_08108_, _07170_, _07161_);
  not (_08109_, _08108_);
  and (_08110_, _08109_, _07171_);
  or (_08111_, _08110_, _07446_);
  or (_08112_, _07200_, _07167_);
  and (_08113_, _08112_, _08111_);
  nand (_08114_, _08113_, _06314_);
  nand (_08115_, _07998_, _07211_);
  nor (_08116_, _06660_, _06652_);
  nor (_08117_, _08116_, _06661_);
  nor (_08118_, _08117_, _06582_);
  not (_08120_, _08118_);
  nor (_08121_, _06692_, _06689_);
  not (_08122_, _08121_);
  nor (_08123_, _06693_, _06678_);
  and (_08124_, _08123_, _08122_);
  not (_08125_, _08124_);
  and (_08126_, _06249_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_08127_, _08089_, _08034_);
  nor (_08128_, _08127_, _08126_);
  nor (_08129_, _08128_, _06724_);
  nor (_08130_, _08129_, _08038_);
  nand (_08131_, _06184_, _06128_);
  and (_08132_, _06248_, _06131_);
  not (_08133_, _08132_);
  and (_08134_, _08133_, _08131_);
  and (_08135_, _06227_, _06118_);
  not (_08136_, _08135_);
  and (_08137_, _08136_, _08033_);
  and (_08138_, _08137_, _08134_);
  and (_08139_, _08138_, _08029_);
  and (_08140_, _08139_, _08130_);
  and (_08141_, _08140_, _08125_);
  and (_08142_, _08141_, _08120_);
  and (_08143_, _08142_, _08115_);
  nand (_08144_, _08143_, _08114_);
  or (_08145_, _08144_, _07668_);
  or (_08146_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_08147_, _08146_, _05552_);
  and (_07085_, _08147_, _08145_);
  and (_08148_, _08102_, _07445_);
  and (_08149_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_08150_, _08149_, _07485_);
  or (_08151_, _08150_, _08148_);
  and (_08152_, _06635_, _06118_);
  and (_08153_, _06746_, _06111_);
  and (_08154_, _07326_, _06386_);
  nor (_08155_, _08154_, _06253_);
  nor (_08156_, _07319_, _06142_);
  nor (_08157_, _08156_, _08155_);
  nor (_08158_, _08157_, _06635_);
  and (_08159_, _08157_, _06635_);
  or (_08160_, _08159_, _06267_);
  nor (_08161_, _08160_, _08158_);
  and (_08162_, _06295_, _06248_);
  or (_08163_, _08162_, _08161_);
  or (_08164_, _08163_, _08153_);
  and (_08165_, _07117_, _06314_);
  nor (_08166_, _07290_, _07286_);
  nor (_08167_, _08166_, _07291_);
  and (_08168_, _08167_, _06677_);
  and (_08169_, _07726_, _07211_);
  or (_08170_, _08169_, _08168_);
  or (_08171_, _08170_, _08165_);
  or (_08172_, _08171_, _08164_);
  nor (_08173_, _08172_, _08152_);
  nand (_08174_, _08173_, _07485_);
  and (_08175_, _08174_, _05552_);
  and (_07107_, _08175_, _08151_);
  and (_08176_, _08144_, _07445_);
  and (_08177_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_08178_, _08177_, _07485_);
  or (_08179_, _08178_, _08176_);
  and (_08180_, _06631_, _06118_);
  and (_08181_, _06500_, _06746_);
  nor (_08182_, _07492_, _06253_);
  nor (_08183_, _07320_, _06142_);
  nor (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _06373_);
  nor (_08186_, _08184_, _06373_);
  nor (_08187_, _08186_, _08185_);
  nor (_08188_, _08187_, _06267_);
  and (_08189_, _06295_, _06227_);
  or (_08190_, _08189_, _08188_);
  or (_08191_, _08190_, _08181_);
  and (_08192_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_08193_, _07294_, _07291_);
  nor (_08194_, _08193_, _07295_);
  and (_08195_, _08194_, _06677_);
  and (_08196_, _07722_, _07211_);
  or (_08197_, _08196_, _08195_);
  or (_08198_, _08197_, _08192_);
  or (_08199_, _08198_, _08191_);
  nor (_08200_, _08199_, _08180_);
  nand (_08201_, _08200_, _07485_);
  and (_08202_, _08201_, _05552_);
  and (_07109_, _08202_, _08179_);
  and (_08203_, _07711_, _07445_);
  and (_08204_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_08205_, _08204_, _07485_);
  or (_08206_, _08205_, _08203_);
  and (_08207_, _07285_, _06712_);
  nor (_08208_, _08207_, _07286_);
  and (_08209_, _08208_, _06677_);
  nand (_08210_, _07200_, _06314_);
  nor (_08211_, _06783_, _06725_);
  not (_08212_, _08211_);
  nor (_08213_, _08212_, _06795_);
  nor (_08214_, _08213_, _06639_);
  and (_08215_, _08213_, _06639_);
  nor (_08216_, _08215_, _08214_);
  and (_08217_, _08216_, _06266_);
  and (_08218_, _06639_, _06118_);
  and (_08219_, _06402_, _07211_);
  and (_08220_, _06162_, _06746_);
  nor (_08221_, _06785_, _06206_);
  or (_08222_, _08221_, _08220_);
  or (_08223_, _08222_, _08219_);
  nor (_08224_, _08223_, _08218_);
  not (_08225_, _08224_);
  nor (_08226_, _08225_, _08217_);
  nand (_08227_, _08226_, _08210_);
  or (_08228_, _08227_, _08209_);
  or (_08229_, _08228_, _07579_);
  and (_08230_, _08229_, _05552_);
  and (_07113_, _08230_, _08206_);
  nor (_08232_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08233_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _07768_);
  nor (_08234_, _08233_, _08232_);
  not (_08235_, \oc8051_symbolic_cxrom1.regvalid [5]);
  not (_08236_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_08237_, _05550_, _08236_);
  and (_08238_, _08237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08239_, _08237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08240_, _08239_, _08238_);
  nor (_08241_, _08240_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08242_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _07768_);
  nor (_08243_, _08242_, _08241_);
  nor (_08244_, _08243_, _08235_);
  and (_08245_, _08243_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_08246_, _08245_, _08244_);
  not (_08247_, _08246_);
  nor (_08248_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08249_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _07768_);
  nor (_08250_, _08249_, _08248_);
  not (_08251_, _08250_);
  and (_08252_, _05550_, _08236_);
  nor (_08253_, _08252_, _08237_);
  nor (_08254_, _08253_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08255_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _07768_);
  nor (_08256_, _08255_, _08254_);
  and (_08257_, _08256_, _08251_);
  nand (_08258_, _08257_, _08247_);
  and (_08259_, _08258_, _08234_);
  nor (_08260_, _08256_, _08251_);
  not (_08261_, _08260_);
  not (_08262_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_08263_, _08243_, _08262_);
  and (_08264_, _08243_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08265_, _08264_, _08263_);
  nor (_08266_, _08265_, _08261_);
  and (_08267_, _08256_, _08250_);
  not (_08268_, _08267_);
  nor (_08269_, _08243_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_08270_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_08271_, _08243_, _08270_);
  or (_08272_, _08271_, _08269_);
  nor (_08273_, _08272_, _08268_);
  nor (_08274_, _08273_, _08266_);
  and (_08275_, _08243_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not (_08276_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_08277_, _08243_, _08276_);
  nor (_08278_, _08277_, _08275_);
  nor (_08279_, _08256_, _08250_);
  not (_08280_, _08279_);
  or (_08281_, _08280_, _08278_);
  and (_08282_, _08281_, _08274_);
  and (_08283_, _08282_, _08259_);
  and (_08284_, _08243_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08285_, _08284_, _08260_);
  not (_08286_, _08243_);
  and (_08288_, _08260_, _08286_);
  and (_08289_, _08288_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08290_, _08289_, _08234_);
  or (_08291_, _08290_, _08285_);
  and (_08292_, _08243_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not (_08293_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08294_, _08243_, _08293_);
  nor (_08295_, _08294_, _08292_);
  nor (_08296_, _08295_, _08280_);
  nor (_08297_, _08243_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_08298_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08299_, _08243_, _08298_);
  or (_08300_, _08299_, _08297_);
  nor (_08301_, _08300_, _08268_);
  not (_08302_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08303_, _08243_, _08302_);
  nor (_08304_, _08243_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08305_, _08304_, _08303_);
  not (_08306_, _08305_);
  and (_08307_, _08306_, _08257_);
  or (_08308_, _08307_, _08301_);
  or (_08309_, _08308_, _08296_);
  nor (_08310_, _08309_, _08291_);
  nor (_08311_, _08310_, _08283_);
  not (_08312_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_08313_, _08234_, _08312_);
  or (_08314_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_08315_, _08314_, _08313_);
  and (_08316_, _08315_, _08267_);
  not (_08317_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_08318_, _08234_, _08317_);
  or (_08319_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_08320_, _08319_, _08318_);
  and (_08321_, _08320_, _08260_);
  or (_08322_, _08321_, _08316_);
  not (_08323_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_08324_, _08234_, _08323_);
  or (_08325_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_08326_, _08325_, _08324_);
  and (_08327_, _08326_, _08257_);
  not (_08328_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_08329_, _08234_, _08328_);
  or (_08330_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_08331_, _08330_, _08329_);
  and (_08332_, _08331_, _08279_);
  or (_08333_, _08332_, _08327_);
  or (_08334_, _08333_, _08322_);
  and (_08335_, _08334_, _08243_);
  not (_08336_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_08337_, _08234_, _08336_);
  or (_08338_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_08339_, _08338_, _08337_);
  and (_08340_, _08339_, _08260_);
  not (_08341_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_08342_, _08234_, _08341_);
  or (_08343_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_08344_, _08343_, _08342_);
  and (_08345_, _08344_, _08267_);
  or (_08346_, _08345_, _08340_);
  not (_08347_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_08348_, _08234_, _08347_);
  or (_08349_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_08350_, _08349_, _08348_);
  and (_08351_, _08350_, _08257_);
  not (_08352_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_08353_, _08234_, _08352_);
  or (_08354_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_08355_, _08354_, _08353_);
  and (_08356_, _08355_, _08279_);
  or (_08357_, _08356_, _08351_);
  or (_08358_, _08357_, _08346_);
  and (_08359_, _08358_, _08286_);
  or (_08360_, _08359_, _08335_);
  and (_08361_, _08360_, _08311_);
  not (_08362_, _08311_);
  and (_08363_, _08362_, word_in[7]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08363_, _08361_);
  nor (_08364_, _06054_, _06043_);
  and (_08365_, _08364_, _06030_);
  not (_08366_, _08365_);
  nor (_08367_, _08366_, _06763_);
  or (_08368_, _08365_, _07468_);
  nand (_08369_, _08368_, _08009_);
  or (_08370_, _08369_, _08367_);
  and (_08371_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_08372_, _08371_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_08373_, _06668_, _06581_);
  and (_08374_, _06698_, _06677_);
  nand (_08375_, _06118_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_08376_, _08375_, _08371_);
  or (_08377_, _08376_, _08374_);
  or (_08378_, _08377_, _08373_);
  and (_08379_, _08378_, _08372_);
  or (_08380_, _08379_, _08009_);
  and (_08381_, _08380_, _08370_);
  or (_08382_, _08381_, _06531_);
  nor (_08383_, _06498_, _06133_);
  not (_08384_, _08383_);
  and (_08385_, _08384_, _07559_);
  and (_08386_, _08385_, _07546_);
  nand (_08387_, _08386_, _06531_);
  and (_08388_, _08387_, _05552_);
  and (_07139_, _08388_, _08382_);
  not (_08389_, _08234_);
  and (_08390_, _08250_, _08389_);
  not (_08391_, _08390_);
  and (_08392_, _08250_, _08234_);
  nor (_08393_, _08392_, _08256_);
  and (_08394_, _08392_, _08256_);
  nor (_08395_, _08394_, _08393_);
  not (_08396_, _08395_);
  nor (_08397_, _08396_, _08272_);
  and (_08398_, _08394_, _08286_);
  or (_08399_, _08394_, _08286_);
  not (_08400_, _08399_);
  nor (_08401_, _08400_, _08398_);
  nor (_08402_, _08401_, _08395_);
  and (_08403_, _08402_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08404_, _08393_, _08286_);
  and (_08405_, _08394_, _08243_);
  nor (_08406_, _08405_, _08404_);
  nor (_08407_, _08406_, _08262_);
  or (_08408_, _08407_, _08403_);
  nor (_08409_, _08408_, _08397_);
  nor (_08410_, _08409_, _08391_);
  not (_08411_, _08392_);
  nor (_08412_, _08396_, _08305_);
  nor (_08413_, _08406_, _08293_);
  nor (_08414_, _08413_, _08412_);
  or (_08415_, _08414_, _08411_);
  nand (_08416_, _08398_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08417_, _08416_, _08415_);
  not (_08418_, _08417_);
  nor (_08419_, _08418_, _08410_);
  and (_08420_, _08251_, _08234_);
  not (_08421_, _08420_);
  nor (_08422_, _08396_, _08300_);
  and (_08423_, _08402_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_08424_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_08425_, _08406_, _08424_);
  or (_08426_, _08425_, _08423_);
  nor (_08427_, _08426_, _08422_);
  nor (_08428_, _08427_, _08421_);
  nor (_08429_, _08250_, _08234_);
  not (_08430_, _08429_);
  nor (_08431_, _08396_, _08246_);
  and (_08432_, _08402_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_08433_, _08406_, _08276_);
  or (_08434_, _08433_, _08432_);
  nor (_08436_, _08434_, _08431_);
  nor (_08437_, _08436_, _08430_);
  nor (_08438_, _08437_, _08428_);
  and (_08439_, _08438_, _08419_);
  or (_08440_, _08429_, _08392_);
  not (_08441_, _08440_);
  not (_08442_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_08443_, _08234_, _08442_);
  or (_08445_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_08446_, _08445_, _08443_);
  and (_08447_, _08446_, _08441_);
  not (_08448_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_08449_, _08234_, _08448_);
  or (_08450_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_08451_, _08450_, _08449_);
  and (_08452_, _08451_, _08440_);
  or (_08453_, _08452_, _08447_);
  and (_08454_, _08453_, _08402_);
  not (_08455_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_08456_, _08234_, _08455_);
  or (_08457_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_08458_, _08457_, _08456_);
  and (_08459_, _08458_, _08441_);
  not (_08460_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_08461_, _08234_, _08460_);
  or (_08462_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_08463_, _08462_, _08461_);
  and (_08464_, _08463_, _08440_);
  nor (_08465_, _08464_, _08459_);
  nor (_08466_, _08465_, _08406_);
  and (_08467_, _08395_, _08286_);
  not (_08468_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_08469_, _08234_, _08468_);
  or (_08470_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_08471_, _08470_, _08469_);
  and (_08472_, _08471_, _08441_);
  not (_08473_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_08474_, _08234_, _08473_);
  or (_08475_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_08476_, _08475_, _08474_);
  and (_08477_, _08476_, _08440_);
  or (_08478_, _08477_, _08472_);
  and (_08479_, _08478_, _08467_);
  and (_08480_, _08395_, _08243_);
  not (_08481_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_08482_, _08234_, _08481_);
  or (_08483_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_08484_, _08483_, _08482_);
  and (_08485_, _08484_, _08441_);
  not (_08486_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_08487_, _08234_, _08486_);
  or (_08488_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_08489_, _08488_, _08487_);
  and (_08490_, _08489_, _08440_);
  or (_08491_, _08490_, _08485_);
  and (_08492_, _08491_, _08480_);
  or (_08493_, _08492_, _08479_);
  or (_08494_, _08493_, _08466_);
  nor (_08495_, _08494_, _08454_);
  nor (_08496_, _08495_, _08439_);
  and (_08497_, _08439_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08497_, _08496_);
  nor (_08498_, _08279_, _08267_);
  not (_08499_, _08498_);
  and (_08500_, _08268_, _08243_);
  and (_08501_, _08267_, _08286_);
  nor (_08502_, _08501_, _08500_);
  and (_08503_, _08502_, _08499_);
  and (_08504_, _08503_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_08505_, _08504_);
  nor (_08506_, _08499_, _08246_);
  nor (_08507_, _08502_, _08498_);
  and (_08508_, _08507_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_08509_, _08508_, _08506_);
  and (_08510_, _08509_, _08505_);
  nor (_08511_, _08510_, _08411_);
  and (_08512_, _08503_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_08513_, _08512_);
  nor (_08514_, _08499_, _08272_);
  and (_08515_, _08507_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08516_, _08515_, _08514_);
  and (_08517_, _08516_, _08513_);
  nor (_08518_, _08517_, _08421_);
  nor (_08519_, _08518_, _08511_);
  nor (_08520_, _08499_, _08300_);
  and (_08521_, _08507_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08522_, _08503_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08523_, _08522_, _08521_);
  nor (_08524_, _08523_, _08520_);
  nor (_08525_, _08524_, _08430_);
  nor (_08526_, _08499_, _08305_);
  and (_08527_, _08507_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08528_, _08503_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_08529_, _08528_, _08527_);
  nor (_08530_, _08529_, _08526_);
  nor (_08531_, _08530_, _08391_);
  nor (_08532_, _08531_, _08525_);
  and (_08533_, _08532_, _08519_);
  and (_08534_, _08344_, _08257_);
  and (_08535_, _08355_, _08267_);
  or (_08536_, _08535_, _08534_);
  and (_08537_, _08350_, _08260_);
  and (_08538_, _08339_, _08279_);
  or (_08539_, _08538_, _08537_);
  or (_08540_, _08539_, _08536_);
  and (_08541_, _08540_, _08502_);
  and (_08542_, _08320_, _08279_);
  and (_08543_, _08331_, _08267_);
  or (_08544_, _08543_, _08542_);
  and (_08545_, _08315_, _08257_);
  and (_08546_, _08326_, _08260_);
  or (_08547_, _08546_, _08545_);
  nor (_08548_, _08547_, _08544_);
  nor (_08549_, _08548_, _08502_);
  nor (_08550_, _08549_, _08541_);
  nor (_08552_, _08550_, _08533_);
  and (_08553_, _08533_, word_in[23]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08553_, _08552_);
  and (_08554_, _08256_, _08243_);
  and (_08555_, _08554_, _08420_);
  and (_08556_, _08555_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08557_, _08430_, _08256_);
  not (_08558_, _08557_);
  nand (_08559_, _08430_, _08256_);
  and (_08561_, _08559_, _08558_);
  not (_08562_, _08561_);
  nor (_08563_, _08305_, _08562_);
  and (_08564_, _08559_, _08243_);
  nor (_08565_, _08559_, _08243_);
  nor (_08566_, _08565_, _08564_);
  nor (_08567_, _08566_, _08561_);
  and (_08568_, _08567_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08569_, _08568_, _08563_);
  nor (_08570_, _08569_, _08421_);
  nor (_08571_, _08300_, _08562_);
  and (_08572_, _08566_, _08562_);
  and (_08573_, _08572_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_08574_, _08567_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08575_, _08574_, _08573_);
  nor (_08576_, _08575_, _08571_);
  nor (_08577_, _08576_, _08411_);
  or (_08578_, _08577_, _08570_);
  nor (_08579_, _08578_, _08556_);
  nor (_08580_, _08562_, _08246_);
  and (_08581_, _08567_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08582_, _08572_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08583_, _08582_, _08581_);
  nor (_08584_, _08583_, _08580_);
  nor (_08585_, _08584_, _08391_);
  nor (_08587_, _08562_, _08272_);
  and (_08588_, _08567_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08589_, _08588_, _08587_);
  nor (_08590_, _08589_, _08430_);
  and (_08592_, _08557_, _08263_);
  or (_08593_, _08592_, _08590_);
  nor (_08594_, _08593_, _08585_);
  and (_08595_, _08594_, _08579_);
  and (_08596_, _08451_, _08441_);
  and (_08598_, _08446_, _08440_);
  or (_08599_, _08598_, _08596_);
  and (_08601_, _08599_, _08567_);
  and (_08602_, _08463_, _08441_);
  and (_08603_, _08458_, _08440_);
  or (_08604_, _08603_, _08602_);
  and (_08605_, _08604_, _08572_);
  and (_08607_, _08561_, _08286_);
  and (_08608_, _08476_, _08441_);
  and (_08609_, _08471_, _08440_);
  or (_08610_, _08609_, _08608_);
  and (_08611_, _08610_, _08607_);
  and (_08613_, _08561_, _08243_);
  and (_08615_, _08489_, _08441_);
  and (_08616_, _08484_, _08440_);
  or (_08618_, _08616_, _08615_);
  and (_08620_, _08618_, _08613_);
  or (_08621_, _08620_, _08611_);
  or (_08622_, _08621_, _08605_);
  nor (_08623_, _08622_, _08601_);
  nor (_08624_, _08623_, _08595_);
  and (_08625_, _08595_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08625_, _08624_);
  and (_08626_, _07731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_08627_, _07733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_08628_, _08627_, _05593_);
  or (_08629_, _08628_, _08626_);
  and (_08630_, _07733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_08631_, _08630_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_08632_, _08631_, _05552_);
  and (_07180_, _08632_, _08629_);
  or (_08633_, _08554_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_07207_, _08633_, _05552_);
  not (_08634_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_08635_, _07433_, _06769_);
  and (_08636_, _08009_, _08635_);
  nor (_08637_, _08636_, _08634_);
  or (_08638_, _08637_, _06531_);
  and (_08639_, _08636_, _08048_);
  or (_08640_, _08639_, _08638_);
  nand (_08641_, _06531_, _06306_);
  and (_08642_, _08641_, _05552_);
  and (_07223_, _08642_, _08640_);
  and (_08643_, _08498_, _08243_);
  and (_08644_, _08533_, _05552_);
  and (_08645_, _08644_, _08420_);
  and (_08646_, _08645_, _08643_);
  not (_08647_, _08646_);
  and (_08648_, _08439_, _05552_);
  and (_08649_, _08648_, _08390_);
  and (_08650_, _08649_, _08480_);
  and (_08651_, _08283_, _05552_);
  and (_08652_, _08651_, _08250_);
  nor (_08653_, _08311_, rst);
  and (_08654_, _08653_, _08554_);
  and (_08655_, _08654_, _08652_);
  and (_08656_, _08653_, word_in[7]);
  and (_08657_, _08656_, _08655_);
  nor (_08658_, _08655_, _08312_);
  nor (_08659_, _08658_, _08657_);
  nor (_08660_, _08659_, _08650_);
  and (_08661_, _08650_, word_in[15]);
  or (_08662_, _08661_, _08660_);
  and (_08663_, _08662_, _08647_);
  and (_08664_, _08595_, _05552_);
  and (_08665_, _08664_, _08429_);
  and (_08666_, _08665_, _08554_);
  and (_08667_, _08644_, word_in[23]);
  and (_08668_, _08667_, _08646_);
  or (_08669_, _08668_, _08666_);
  or (_08670_, _08669_, _08663_);
  not (_08671_, _08666_);
  and (_08672_, _08664_, word_in[31]);
  or (_08673_, _08672_, _08671_);
  and (_13877_, _08673_, _08670_);
  or (_08674_, _08572_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_07256_, _08674_, _05552_);
  not (_08675_, _05546_);
  or (_08676_, _05641_, _08675_);
  or (_08677_, _05546_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_08678_, _08677_, _05552_);
  and (_07268_, _08678_, _08676_);
  or (_08679_, _08280_, _08243_);
  not (_08680_, _08679_);
  nor (_08681_, _08405_, _08680_);
  and (_08682_, _08554_, _08390_);
  nor (_08683_, _08682_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand (_08684_, _08683_, _08681_);
  and (_07287_, _08684_, _05552_);
  and (_08685_, _08404_, _08250_);
  nor (_08686_, _08685_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_08687_, _08686_, _08681_);
  and (_07324_, _08687_, _05552_);
  or (_08688_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not (_08689_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_08690_, _05550_, _08689_);
  and (_08691_, _08690_, _05552_);
  and (_07338_, _08691_, _08688_);
  or (_08692_, _05733_, _08675_);
  or (_08693_, _05546_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_08694_, _08693_, _05552_);
  and (_07341_, _08694_, _08692_);
  or (_08695_, _08411_, _08243_);
  nor (_08696_, _08695_, _08256_);
  or (_08697_, _08256_, _08243_);
  or (_08698_, _08697_, _08390_);
  and (_08699_, _08698_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_08700_, _08699_, _08696_);
  and (_08701_, _08700_, _08406_);
  and (_08702_, _08279_, _08263_);
  or (_08703_, _08702_, _08685_);
  or (_08704_, _08703_, _08701_);
  and (_08706_, _08704_, _08681_);
  or (_08707_, _08702_, _08700_);
  and (_08708_, _08707_, _08405_);
  or (_08710_, _08708_, _08680_);
  or (_08711_, _08710_, _08706_);
  and (_07361_, _08711_, _05552_);
  nand (_08713_, _05665_, _05546_);
  or (_08714_, _05546_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_08716_, _08714_, _05552_);
  and (_07409_, _08716_, _08713_);
  not (_08718_, _08256_);
  nor (_08720_, _08718_, _08243_);
  and (_08722_, _08720_, _08429_);
  or (_08723_, _08696_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08725_, _08723_, _08722_);
  and (_08726_, _08725_, _08406_);
  or (_08727_, _08722_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_08728_, _08727_, _08405_);
  and (_08729_, _08420_, _08607_);
  and (_08730_, _08557_, _08286_);
  and (_08731_, _08730_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08732_, _08731_, _08729_);
  or (_08733_, _08732_, _08728_);
  or (_08734_, _08733_, _08685_);
  or (_08735_, _08734_, _08726_);
  and (_07415_, _08735_, _05552_);
  nor (_08736_, _08267_, _08243_);
  not (_08737_, _08736_);
  or (_08738_, _08722_, _08696_);
  or (_08739_, _08738_, _08737_);
  and (_08740_, _08739_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08741_, _08420_, _08720_);
  and (_08742_, _08393_, _08244_);
  or (_08743_, _08742_, _08741_);
  or (_08744_, _08743_, _08740_);
  or (_08745_, _08400_, _08565_);
  and (_08746_, _08745_, _08744_);
  and (_08747_, _08561_, _08244_);
  or (_08748_, _08747_, _08722_);
  or (_08749_, _08748_, _08746_);
  and (_08750_, _08749_, _08682_);
  or (_08751_, _08720_, _08500_);
  and (_08752_, _08749_, _08751_);
  and (_08753_, _08744_, _08405_);
  nor (_08754_, _08679_, _08235_);
  or (_08755_, _08754_, _08685_);
  or (_08756_, _08755_, _08696_);
  or (_08757_, _08756_, _08753_);
  or (_08758_, _08757_, _08752_);
  or (_08759_, _08758_, _08750_);
  and (_07480_, _08759_, _05552_);
  and (_08760_, _06569_, _05822_);
  and (_08761_, _06569_, _05737_);
  nand (_08762_, _06576_, _08761_);
  or (_08763_, _08762_, _06572_);
  and (_08764_, _08763_, _01436_);
  or (_07502_, _08764_, _08760_);
  and (_08765_, _08720_, _08390_);
  or (_08766_, _08765_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08767_, _08765_, _08243_);
  and (_08768_, _08256_, _08234_);
  and (_08769_, _08404_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08770_, _08769_, _08768_);
  or (_08771_, _08770_, _08767_);
  and (_08772_, _08771_, _08766_);
  and (_08773_, _08772_, _08737_);
  and (_08774_, _08738_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08775_, _08774_, _08741_);
  or (_08776_, _08775_, _08773_);
  and (_08777_, _08776_, _08745_);
  and (_08778_, _08766_, _08405_);
  or (_08779_, _08769_, _08696_);
  or (_08780_, _08779_, _08722_);
  or (_08781_, _08780_, _08778_);
  or (_08782_, _08781_, _08777_);
  and (_07541_, _08782_, _05552_);
  and (_08783_, _08243_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08784_, _08730_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08785_, _08607_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_08786_, _08785_, _08722_);
  or (_08787_, _08786_, _08784_);
  or (_08788_, _08741_, _08765_);
  or (_08789_, _08788_, _08787_);
  or (_08790_, _08789_, _08398_);
  or (_08791_, _08790_, _08783_);
  and (_07615_, _08791_, _05552_);
  nor (_08792_, _08607_, _08567_);
  or (_08793_, _08792_, _08398_);
  and (_08794_, _08793_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08795_, _08557_, _08243_);
  not (_08796_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08797_, _08440_, _08796_);
  and (_08798_, _08797_, _08607_);
  and (_08799_, _08738_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08800_, _08799_, _08798_);
  or (_08802_, _08800_, _08795_);
  or (_08803_, _08802_, _08794_);
  and (_08804_, _08803_, _08243_);
  not (_08806_, _08768_);
  and (_08807_, _08736_, _08806_);
  and (_08808_, _08807_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08809_, _08741_, _08398_);
  or (_08811_, _08809_, _08808_);
  or (_08812_, _08811_, _08765_);
  or (_08813_, _08812_, _08804_);
  and (_07673_, _08813_, _05552_);
  nor (_08815_, _08399_, _08557_);
  and (_08816_, _08501_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08818_, _08420_, _08613_);
  or (_08819_, _08818_, _08275_);
  or (_08820_, _08819_, _08816_);
  and (_08821_, _08820_, _08815_);
  or (_08823_, _08741_, _08607_);
  and (_08824_, _08823_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08826_, _08816_, _08795_);
  or (_08827_, _08826_, _08824_);
  or (_08828_, _08827_, _08821_);
  and (_08829_, _08828_, _08400_);
  and (_08830_, _08736_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08831_, _08830_, _08765_);
  and (_08832_, _08820_, _08405_);
  or (_08833_, _08832_, _08398_);
  or (_08834_, _08833_, _08831_);
  or (_08835_, _08834_, _08829_);
  and (_07739_, _08835_, _05552_);
  not (_08836_, rxd_i);
  and (_08837_, _07734_, _05564_);
  and (_08838_, _07736_, _08837_);
  nand (_08839_, _08838_, _08836_);
  or (_08840_, _08838_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_08841_, _08840_, _05552_);
  and (_07822_, _08841_, _08839_);
  and (_08842_, _08280_, _08243_);
  and (_08843_, _08765_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08844_, _08738_, _08741_);
  and (_08846_, _08844_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08847_, _08846_, _08843_);
  and (_08848_, _08730_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08849_, _08643_, _08390_);
  or (_08850_, _08256_, _08234_);
  and (_08851_, _08850_, _08284_);
  or (_08852_, _08851_, _08849_);
  or (_08853_, _08852_, _08848_);
  and (_08854_, _08441_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08855_, _08854_, _08607_);
  or (_08856_, _08795_, _08398_);
  and (_08857_, _08856_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08858_, _08857_, _08855_);
  or (_08859_, _08858_, _08853_);
  or (_08860_, _08859_, _08847_);
  and (_08861_, _08860_, _08842_);
  and (_08862_, _08498_, _08286_);
  and (_08863_, _08862_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08864_, _08680_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08865_, _08864_, _08398_);
  or (_08866_, _08865_, _08843_);
  or (_08867_, _08866_, _08863_);
  or (_08868_, _08867_, _08818_);
  or (_08869_, _08868_, _08861_);
  or (_08870_, _08869_, _08795_);
  and (_07829_, _08870_, _05552_);
  or (_08871_, _08628_, _07731_);
  and (_08872_, _08871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  and (_08873_, _08627_, _05563_);
  and (_08874_, _07736_, _08873_);
  or (_08875_, _08874_, _08872_);
  and (_07858_, _08875_, _05552_);
  and (_08876_, _08730_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08877_, _08467_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08878_, _08398_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08879_, _08440_, _08697_);
  and (_08880_, _08879_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08881_, _08880_, _08878_);
  or (_08882_, _08881_, _08877_);
  or (_08883_, _08882_, _08795_);
  or (_08884_, _08883_, _08876_);
  or (_08885_, _08405_, _08480_);
  and (_08886_, _08680_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08887_, _08720_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08888_, _08887_, _08886_);
  and (_08889_, _08288_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08890_, _08260_, _08243_);
  or (_08891_, _08234_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08892_, _08891_, _08890_);
  and (_08893_, _08264_, _08261_);
  or (_08894_, _08893_, _08892_);
  or (_08895_, _08894_, _08889_);
  or (_08896_, _08895_, _08888_);
  and (_08897_, _08896_, _08885_);
  or (_08898_, _08897_, _08884_);
  or (_08900_, _08898_, _08818_);
  or (_08901_, _08900_, _08849_);
  and (_07927_, _08901_, _05552_);
  nand (_08903_, _07600_, _07260_);
  or (_08904_, _07574_, _06972_);
  nor (_08905_, _07264_, _06396_);
  nor (_08906_, _08905_, _06973_);
  nor (_08908_, _08365_, _06396_);
  nor (_08909_, _08908_, _08367_);
  and (_08910_, _07261_, _06972_);
  and (_08911_, _08910_, _07269_);
  not (_08913_, _08911_);
  or (_08914_, _08913_, _08909_);
  and (_08915_, _08914_, _08906_);
  nor (_08917_, _08915_, _07260_);
  nand (_08918_, _08917_, _08904_);
  nand (_08920_, _08918_, _08903_);
  and (_07968_, _08920_, _05552_);
  nand (_08921_, _08102_, _06973_);
  and (_08923_, _08910_, _07264_);
  not (_08924_, _08923_);
  not (_08925_, _06056_);
  nor (_08926_, _06763_, _08925_);
  nor (_08927_, _06056_, _06243_);
  nor (_08928_, _08927_, _08926_);
  or (_08929_, _08928_, _08924_);
  and (_08930_, _06020_, _05989_);
  and (_08931_, _07262_, _08930_);
  and (_08932_, _08931_, _06911_);
  and (_08933_, _08932_, _06775_);
  not (_08934_, _08933_);
  and (_08935_, _08934_, _08910_);
  and (_08936_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_08937_, _08936_, _07260_);
  and (_08938_, _08937_, _08929_);
  nand (_08939_, _08938_, _08921_);
  and (_08940_, _08173_, _07260_);
  not (_08941_, _08940_);
  and (_08942_, _08941_, _08939_);
  and (_07973_, _08942_, _05552_);
  and (_08943_, _08554_, _08430_);
  and (_08944_, _08943_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08945_, _08795_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08946_, _08643_, _08806_);
  or (_08947_, _08946_, _08945_);
  and (_08948_, _08250_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08949_, _08948_, _08607_);
  nor (_08950_, _08679_, _08302_);
  and (_08951_, _08720_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_08952_, _08951_, _08818_);
  or (_08953_, _08952_, _08950_);
  or (_08954_, _08953_, _08949_);
  or (_08955_, _08954_, _08947_);
  or (_08956_, _08955_, _08944_);
  and (_08032_, _08956_, _05552_);
  nand (_08957_, _08411_, _08243_);
  and (_08958_, _08957_, _08695_);
  nor (_08959_, _08958_, _08806_);
  nor (_08960_, _08959_, _08393_);
  and (_08961_, _08718_, _08243_);
  or (_08962_, _08961_, _08398_);
  or (_08963_, _08962_, _08960_);
  and (_08964_, _08963_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_08965_, _08964_, _08251_);
  and (_08966_, _08965_, _08554_);
  not (_08967_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_08968_, _08842_, _08967_);
  or (_08969_, _08968_, _08890_);
  or (_08970_, _08969_, _08966_);
  and (_08119_, _08970_, _05552_);
  or (_08971_, _08480_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08231_, _08971_, _05552_);
  not (_08972_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_08973_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor (_08974_, _08973_, _08972_);
  and (_08975_, _08973_, _08972_);
  nor (_08976_, _08975_, _08974_);
  not (_08977_, _08976_);
  and (_08978_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_08979_, _08978_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_08980_, _08978_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_08981_, _08980_, _08979_);
  or (_08982_, _08981_, _08973_);
  and (_08983_, _08982_, _08977_);
  nor (_08984_, _08974_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_08985_, _08974_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_08986_, _08985_, _08984_);
  or (_08987_, _08979_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_10089_, _08987_, _05552_);
  and (_08988_, _10089_, _08986_);
  and (_08435_, _08988_, _08983_);
  nor (_08989_, _06967_, _06020_);
  and (_08990_, _08989_, _06060_);
  and (_08991_, _08990_, _07443_);
  not (_08992_, _08991_);
  not (_08993_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_08994_, _08993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not (_08995_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_08996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_08997_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_08998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_08999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _08998_);
  nor (_09000_, _08999_, _08997_);
  nor (_09001_, _09000_, _08996_);
  or (_09002_, _09001_, _08995_);
  and (_09003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _08998_);
  and (_09004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_09005_, _09004_, _09003_);
  nor (_09006_, _09005_, _08996_);
  not (_09007_, _09006_);
  and (_09008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_09009_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _08998_);
  nor (_09010_, _09009_, _09008_);
  nor (_09012_, _09010_, _08996_);
  nand (_09013_, _09012_, _09007_);
  or (_09014_, _09013_, _09002_);
  and (_09015_, _09014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_09017_, _09015_, _08994_);
  nor (_09018_, _06054_, _06020_);
  and (_09019_, _09018_, _07433_);
  and (_09020_, _09019_, _07443_);
  and (_09021_, _09020_, _06775_);
  or (_09022_, _09021_, _09017_);
  and (_09023_, _09022_, _08992_);
  nand (_09024_, _09021_, _06763_);
  and (_09025_, _09024_, _09023_);
  nor (_09026_, _08992_, _06306_);
  or (_09027_, _09026_, _09025_);
  and (_08444_, _09027_, _05552_);
  and (_09028_, _07936_, _06308_);
  and (_09029_, _09028_, _06068_);
  not (_09030_, _09029_);
  and (_09031_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_09032_, _09028_, _07946_);
  or (_09033_, _09032_, _09031_);
  and (_08551_, _09033_, _05552_);
  and (_09035_, _05552_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_09036_, _09035_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_09038_, _05547_, _05671_);
  not (_09039_, _09038_);
  not (_09040_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_09041_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_09042_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_09043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_09044_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_09045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_09046_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_09047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_09048_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_09049_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_09050_, _09049_, _09048_);
  and (_09051_, _09050_, _09047_);
  and (_09052_, _09051_, _09046_);
  and (_09053_, _09052_, _09045_);
  and (_09054_, _09053_, _09044_);
  and (_09055_, _09054_, _09043_);
  and (_09056_, _09055_, _09042_);
  and (_09057_, _09056_, _09041_);
  and (_09058_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_09059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_09060_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_09061_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_09062_, _09061_, _09059_);
  and (_09063_, _09062_, _09060_);
  nor (_09064_, _09063_, _09059_);
  nor (_09065_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_09066_, _09065_, _09058_);
  not (_09067_, _09066_);
  nor (_09068_, _09067_, _09064_);
  nor (_09069_, _09068_, _09058_);
  and (_09070_, _09069_, _09057_);
  and (_09071_, _09070_, _09040_);
  nor (_09072_, _09071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_09073_, _09071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_09074_, _09073_, _09072_);
  not (_09075_, _09074_);
  nor (_09076_, _09070_, _09040_);
  nor (_09077_, _09076_, _09071_);
  not (_09078_, _09077_);
  not (_09079_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_09080_, _09069_, _09054_);
  and (_09081_, _09080_, _09043_);
  and (_09082_, _09081_, _09042_);
  and (_09083_, _09082_, _09079_);
  nor (_09084_, _09083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_09085_, _09083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_09086_, _09085_, _09084_);
  nor (_09087_, _09082_, _09079_);
  nor (_09088_, _09087_, _09083_);
  not (_09089_, _09088_);
  nor (_09090_, _09081_, _09042_);
  or (_09091_, _09090_, _09082_);
  nor (_09092_, _09080_, _09043_);
  nor (_09093_, _09092_, _09081_);
  not (_09094_, _09093_);
  and (_09095_, _09069_, _09053_);
  nor (_09096_, _09095_, _09044_);
  nor (_09097_, _09096_, _09080_);
  not (_09098_, _09097_);
  and (_09099_, _09069_, _09051_);
  nor (_09100_, _09099_, _09046_);
  and (_09101_, _09069_, _09052_);
  or (_09102_, _09101_, _09100_);
  and (_09103_, _09069_, _09050_);
  nor (_09104_, _09103_, _09047_);
  or (_09105_, _09104_, _09099_);
  not (_09106_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_09107_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_09108_, _09069_, _09048_);
  and (_09109_, _09108_, _09107_);
  nor (_09111_, _09109_, _09106_);
  or (_09112_, _09111_, _09103_);
  nor (_09113_, _09069_, _09048_);
  nor (_09114_, _09113_, _09108_);
  not (_09116_, _09114_);
  nor (_09117_, _09062_, _09060_);
  nor (_09118_, _09117_, _09063_);
  not (_09119_, _09118_);
  nor (_09121_, _09119_, _07919_);
  not (_09122_, _09121_);
  not (_09123_, _07930_);
  nor (_09124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_09126_, _09124_, _09060_);
  and (_09127_, _09126_, _09123_);
  and (_09128_, _09119_, _07919_);
  nor (_09130_, _09128_, _09121_);
  nand (_09131_, _09130_, _09127_);
  and (_09132_, _09131_, _09122_);
  not (_09133_, _09132_);
  and (_09135_, _09067_, _09064_);
  nor (_09136_, _09135_, _09068_);
  and (_09137_, _09136_, _09133_);
  and (_09139_, _09137_, _09116_);
  nor (_09140_, _09108_, _09107_);
  or (_09142_, _09140_, _09109_);
  and (_09143_, _09142_, _09139_);
  and (_09144_, _09143_, _09112_);
  and (_09145_, _09144_, _09105_);
  and (_09146_, _09145_, _09102_);
  nor (_09147_, _09101_, _09045_);
  or (_09148_, _09147_, _09095_);
  and (_09149_, _09148_, _09146_);
  and (_09150_, _09149_, _09098_);
  and (_09151_, _09150_, _09094_);
  and (_09152_, _09151_, _09091_);
  and (_09153_, _09152_, _09089_);
  and (_09154_, _09153_, _09086_);
  and (_09155_, _09154_, _09078_);
  nor (_09156_, _09155_, _09075_);
  and (_09157_, _09155_, _09075_);
  or (_09158_, _09157_, _09156_);
  or (_09159_, _09158_, _09039_);
  or (_09160_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_09161_, _09160_, _07933_);
  and (_09162_, _09161_, _09159_);
  or (_08560_, _09162_, _09036_);
  and (_09163_, _08653_, _08250_);
  nor (_09165_, _09163_, _08651_);
  and (_09166_, _08653_, _08697_);
  not (_09167_, _09166_);
  and (_09168_, _09167_, _09165_);
  and (_09169_, _09168_, _08653_);
  not (_09170_, _09169_);
  and (_09171_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_09172_, _08653_, word_in[0]);
  and (_09173_, _09172_, _09168_);
  or (_09174_, _09173_, _09171_);
  and (_09175_, _08648_, _08405_);
  not (_09176_, _09175_);
  and (_09177_, _09176_, _09174_);
  and (_09178_, _08644_, _08682_);
  and (_09179_, _08405_, word_in[8]);
  and (_09180_, _09179_, _08648_);
  or (_09181_, _09180_, _09178_);
  or (_09182_, _09181_, _09177_);
  and (_09183_, _08664_, _08555_);
  not (_09184_, _09183_);
  not (_09185_, _09178_);
  or (_09186_, _09185_, word_in[16]);
  and (_09187_, _09186_, _09184_);
  and (_09188_, _09187_, _09182_);
  and (_09189_, _08664_, word_in[24]);
  and (_09190_, _09189_, _08555_);
  or (_08586_, _09190_, _09188_);
  and (_09191_, _08664_, word_in[25]);
  and (_09192_, _09191_, _08555_);
  and (_09193_, _09178_, word_in[17]);
  and (_09194_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_09195_, _08653_, word_in[1]);
  and (_09196_, _09195_, _09168_);
  or (_09197_, _09196_, _09194_);
  or (_09198_, _09197_, _09175_);
  or (_09199_, _09176_, word_in[9]);
  and (_09200_, _09199_, _09185_);
  and (_09201_, _09200_, _09198_);
  or (_09202_, _09201_, _09193_);
  and (_09203_, _09202_, _09184_);
  or (_08591_, _09203_, _09192_);
  and (_09204_, _08664_, word_in[26]);
  and (_09205_, _09204_, _08555_);
  and (_09206_, _09178_, word_in[18]);
  and (_09207_, _08653_, word_in[2]);
  and (_09208_, _09207_, _09168_);
  and (_09209_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  or (_09210_, _09209_, _09208_);
  or (_09211_, _09210_, _09175_);
  or (_09212_, _09176_, word_in[10]);
  and (_09213_, _09212_, _09185_);
  and (_09214_, _09213_, _09211_);
  or (_09215_, _09214_, _09206_);
  and (_09216_, _09215_, _09184_);
  or (_08597_, _09216_, _09205_);
  and (_09218_, _08664_, word_in[27]);
  and (_09219_, _09218_, _08555_);
  and (_09221_, _09178_, word_in[19]);
  and (_09222_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_09223_, _08653_, word_in[3]);
  and (_09225_, _09223_, _09168_);
  or (_09226_, _09225_, _09222_);
  or (_09227_, _09226_, _09175_);
  or (_09228_, _09176_, word_in[11]);
  and (_09230_, _09228_, _09185_);
  and (_09231_, _09230_, _09227_);
  or (_09232_, _09231_, _09221_);
  and (_09234_, _09232_, _09184_);
  or (_08600_, _09234_, _09219_);
  and (_09236_, _08664_, word_in[28]);
  and (_09237_, _09236_, _08555_);
  and (_09239_, _09178_, word_in[20]);
  and (_09240_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_09241_, _08653_, word_in[4]);
  and (_09243_, _09241_, _09169_);
  or (_09244_, _09243_, _09240_);
  or (_09245_, _09244_, _09175_);
  or (_09246_, _09176_, word_in[12]);
  and (_09247_, _09246_, _09185_);
  and (_09248_, _09247_, _09245_);
  or (_09249_, _09248_, _09239_);
  and (_09250_, _09249_, _09184_);
  or (_08606_, _09250_, _09237_);
  and (_09251_, _08664_, word_in[29]);
  and (_09252_, _09251_, _08555_);
  and (_09253_, _08653_, word_in[5]);
  and (_09254_, _09253_, _09168_);
  and (_09255_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  or (_09256_, _09255_, _09254_);
  or (_09257_, _09256_, _09175_);
  or (_09258_, _09176_, word_in[13]);
  and (_09259_, _09258_, _09185_);
  and (_09260_, _09259_, _09257_);
  and (_09261_, _09178_, word_in[21]);
  or (_09262_, _09261_, _09260_);
  and (_09263_, _09262_, _09184_);
  or (_08612_, _09263_, _09252_);
  and (_09264_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_09265_, _09028_, _07976_);
  or (_09266_, _09265_, _09264_);
  and (_08614_, _09266_, _05552_);
  and (_09267_, _08664_, word_in[30]);
  and (_09268_, _09267_, _08555_);
  and (_09269_, _08653_, word_in[6]);
  and (_09270_, _09269_, _09168_);
  and (_09271_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or (_09272_, _09271_, _09270_);
  or (_09273_, _09272_, _09175_);
  or (_09274_, _09176_, word_in[14]);
  and (_09275_, _09274_, _09185_);
  and (_09276_, _09275_, _09273_);
  and (_09277_, _09178_, word_in[22]);
  or (_09278_, _09277_, _09276_);
  and (_09279_, _09278_, _09184_);
  or (_08617_, _09279_, _09268_);
  and (_09280_, _09178_, word_in[23]);
  not (_09281_, word_in[15]);
  nand (_09282_, _09175_, _09281_);
  and (_09283_, _09282_, _09185_);
  and (_09284_, _09169_, word_in[7]);
  nor (_09285_, _09169_, _08460_);
  or (_09286_, _09285_, _09284_);
  or (_09287_, _09286_, _09175_);
  and (_09288_, _09287_, _09283_);
  or (_09289_, _09288_, _09280_);
  and (_09290_, _09289_, _09184_);
  and (_09291_, _09183_, word_in[31]);
  or (_08619_, _09291_, _09290_);
  and (_09292_, _08664_, _08682_);
  not (_09293_, _09292_);
  and (_09294_, _08644_, _08392_);
  and (_09295_, _09294_, _08503_);
  not (_09296_, _09295_);
  not (_09297_, _08406_);
  and (_09298_, _08648_, _08429_);
  and (_09299_, _09298_, _09297_);
  and (_09300_, _08651_, _08251_);
  not (_09301_, _09300_);
  nor (_09302_, _09301_, _09166_);
  and (_09303_, _09302_, _09172_);
  not (_09304_, _09302_);
  and (_09305_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_09306_, _09305_, _09303_);
  nor (_09307_, _09306_, _09299_);
  and (_09308_, _09299_, word_in[8]);
  or (_09309_, _09308_, _09307_);
  and (_09310_, _09309_, _09296_);
  and (_09311_, _08644_, word_in[16]);
  and (_09312_, _09295_, _09311_);
  or (_09313_, _09312_, _09310_);
  and (_09314_, _09313_, _09293_);
  and (_09315_, _09292_, word_in[24]);
  or (_08705_, _09315_, _09314_);
  and (_09316_, _08644_, word_in[17]);
  and (_09317_, _09295_, _09316_);
  and (_09318_, _09302_, _09195_);
  and (_09319_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_09320_, _09319_, _09318_);
  nor (_09321_, _09320_, _09299_);
  and (_09322_, _09299_, word_in[9]);
  or (_09323_, _09322_, _09321_);
  and (_09324_, _09323_, _09296_);
  or (_09325_, _09324_, _09317_);
  and (_09326_, _09325_, _09293_);
  and (_09327_, _09292_, word_in[25]);
  or (_08709_, _09327_, _09326_);
  and (_09328_, _09302_, _09207_);
  and (_09329_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_09330_, _09329_, _09328_);
  nor (_09331_, _09330_, _09299_);
  and (_09332_, _09299_, word_in[10]);
  or (_09333_, _09332_, _09331_);
  and (_09334_, _09333_, _09296_);
  and (_09335_, _08644_, word_in[18]);
  and (_09336_, _09295_, _09335_);
  or (_09337_, _09336_, _09334_);
  and (_09338_, _09337_, _09293_);
  and (_09339_, _09292_, word_in[26]);
  or (_08712_, _09339_, _09338_);
  and (_09340_, _08644_, word_in[19]);
  and (_09341_, _09295_, _09340_);
  and (_09342_, _09302_, _09223_);
  and (_09343_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_09344_, _09343_, _09342_);
  nor (_09345_, _09344_, _09299_);
  and (_09346_, _09299_, word_in[11]);
  or (_09347_, _09346_, _09345_);
  and (_09348_, _09347_, _09296_);
  or (_09349_, _09348_, _09341_);
  and (_09350_, _09349_, _09293_);
  and (_09351_, _09292_, word_in[27]);
  or (_08715_, _09351_, _09350_);
  and (_09352_, _09302_, _09241_);
  and (_09353_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_09354_, _09353_, _09352_);
  nor (_09355_, _09354_, _09299_);
  and (_09356_, _09299_, word_in[12]);
  or (_09357_, _09356_, _09355_);
  and (_09358_, _09357_, _09296_);
  and (_09359_, _08644_, word_in[20]);
  and (_09360_, _09295_, _09359_);
  or (_09361_, _09360_, _09358_);
  and (_09362_, _09361_, _09293_);
  and (_09363_, _09292_, word_in[28]);
  or (_08717_, _09363_, _09362_);
  and (_09364_, _08644_, word_in[21]);
  and (_09365_, _09295_, _09364_);
  and (_09366_, _09302_, _09253_);
  and (_09367_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_09368_, _09367_, _09366_);
  nor (_09369_, _09368_, _09299_);
  and (_09370_, _09299_, word_in[13]);
  or (_09371_, _09370_, _09369_);
  and (_09372_, _09371_, _09296_);
  or (_09373_, _09372_, _09365_);
  and (_09374_, _09373_, _09293_);
  and (_09375_, _09292_, word_in[29]);
  or (_08719_, _09375_, _09374_);
  and (_09376_, _09302_, _09269_);
  and (_09377_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_09378_, _09377_, _09376_);
  nor (_09379_, _09378_, _09299_);
  and (_09380_, _09299_, word_in[14]);
  or (_09381_, _09380_, _09379_);
  and (_09382_, _09381_, _09296_);
  and (_09383_, _08644_, word_in[22]);
  and (_09384_, _09295_, _09383_);
  or (_09385_, _09384_, _09382_);
  and (_09386_, _09385_, _09293_);
  and (_09387_, _09292_, word_in[30]);
  or (_08721_, _09387_, _09386_);
  nor (_09388_, _09302_, _08352_);
  and (_09389_, _09302_, _08656_);
  or (_09390_, _09389_, _09388_);
  or (_09391_, _09390_, _09299_);
  nand (_09392_, _09299_, _09281_);
  and (_09393_, _09392_, _09391_);
  or (_09394_, _09393_, _09295_);
  or (_09395_, _09296_, _08667_);
  and (_09396_, _09395_, _09293_);
  and (_09397_, _09396_, _09394_);
  and (_09398_, _09292_, word_in[31]);
  or (_08724_, _09398_, _09397_);
  and (_09399_, _08664_, _08392_);
  and (_09400_, _09399_, _08572_);
  and (_09401_, _08644_, _08429_);
  and (_09402_, _09401_, _08503_);
  not (_09404_, _09402_);
  and (_09405_, _08648_, _08420_);
  and (_09406_, _09405_, _09297_);
  not (_09407_, _08697_);
  not (_09409_, _08651_);
  and (_09410_, _09163_, _09409_);
  and (_09411_, _09410_, _09407_);
  or (_09412_, _09411_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not (_09413_, _09411_);
  or (_09414_, _09413_, _09172_);
  and (_09415_, _09414_, _09412_);
  or (_09416_, _09415_, _09406_);
  not (_09417_, _09406_);
  or (_09418_, _09417_, word_in[8]);
  and (_09419_, _09418_, _09416_);
  and (_09420_, _09419_, _09404_);
  and (_09421_, _09402_, _09311_);
  or (_09422_, _09421_, _09420_);
  or (_09423_, _09422_, _09400_);
  not (_09424_, _09400_);
  or (_09425_, _09424_, word_in[24]);
  and (_08801_, _09425_, _09423_);
  and (_09426_, _09411_, _09195_);
  and (_09427_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  or (_09428_, _09427_, _09426_);
  and (_09429_, _09428_, _09417_);
  and (_09430_, _09406_, word_in[9]);
  or (_09431_, _09430_, _09429_);
  and (_09432_, _09431_, _09404_);
  and (_09433_, _09402_, _09316_);
  or (_09434_, _09433_, _09400_);
  or (_09435_, _09434_, _09432_);
  or (_09436_, _09424_, word_in[25]);
  and (_08805_, _09436_, _09435_);
  and (_09437_, _09402_, _09335_);
  and (_09438_, _09411_, _09207_);
  and (_09439_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  or (_09440_, _09439_, _09438_);
  or (_09441_, _09440_, _09406_);
  or (_09442_, _09417_, word_in[10]);
  and (_09443_, _09442_, _09404_);
  and (_09444_, _09443_, _09441_);
  or (_09445_, _09444_, _09437_);
  and (_09446_, _09445_, _09424_);
  and (_09447_, _09400_, word_in[26]);
  or (_08810_, _09447_, _09446_);
  and (_09448_, _09411_, _09223_);
  and (_09449_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  or (_09450_, _09449_, _09448_);
  or (_09451_, _09450_, _09406_);
  or (_09452_, _09417_, word_in[11]);
  and (_09453_, _09452_, _09404_);
  and (_09454_, _09453_, _09451_);
  and (_09455_, _09402_, _09340_);
  or (_09456_, _09455_, _09454_);
  and (_09457_, _09456_, _09424_);
  and (_09458_, _09400_, word_in[27]);
  or (_08814_, _09458_, _09457_);
  and (_09459_, _09411_, _09241_);
  and (_09460_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  or (_09461_, _09460_, _09459_);
  or (_09462_, _09461_, _09406_);
  or (_09463_, _09417_, word_in[12]);
  and (_09464_, _09463_, _09404_);
  and (_09465_, _09464_, _09462_);
  and (_09466_, _09402_, _09359_);
  or (_09467_, _09466_, _09400_);
  or (_09468_, _09467_, _09465_);
  or (_09469_, _09424_, word_in[28]);
  and (_08817_, _09469_, _09468_);
  and (_09470_, _09411_, _09253_);
  and (_09471_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or (_09472_, _09471_, _09470_);
  or (_09473_, _09472_, _09406_);
  or (_09474_, _09417_, word_in[13]);
  and (_09475_, _09474_, _09404_);
  and (_09476_, _09475_, _09473_);
  and (_09477_, _09402_, _09364_);
  or (_09478_, _09477_, _09400_);
  or (_09479_, _09478_, _09476_);
  or (_09480_, _09424_, word_in[29]);
  and (_13878_, _09480_, _09479_);
  and (_09481_, _09411_, _09269_);
  and (_09482_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  or (_09483_, _09482_, _09481_);
  or (_09484_, _09483_, _09406_);
  or (_09485_, _09417_, word_in[14]);
  and (_09486_, _09485_, _09404_);
  and (_09487_, _09486_, _09484_);
  and (_09488_, _09402_, _09383_);
  or (_09489_, _09488_, _09400_);
  or (_09490_, _09489_, _09487_);
  or (_09491_, _09424_, word_in[30]);
  and (_08822_, _09491_, _09490_);
  and (_09492_, _09402_, _08667_);
  and (_09493_, _09411_, _08656_);
  nor (_09494_, _09411_, _08455_);
  or (_09495_, _09494_, _09493_);
  or (_09496_, _09495_, _09406_);
  nand (_09497_, _09406_, _09281_);
  and (_09498_, _09497_, _09404_);
  and (_09499_, _09498_, _09496_);
  or (_09500_, _09499_, _09492_);
  and (_09501_, _09500_, _09424_);
  and (_09502_, _09400_, word_in[31]);
  or (_08825_, _09502_, _09501_);
  nor (_09503_, _07949_, _07937_);
  and (_09504_, _07936_, _06065_);
  not (_09505_, _09504_);
  nand (_09506_, _09505_, _09503_);
  nor (_09507_, _09506_, _06069_);
  or (_09508_, _09507_, _06955_);
  and (_09509_, _09508_, _09030_);
  or (_09510_, _09509_, _06069_);
  and (_09511_, _09510_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_09512_, _09030_, _06306_);
  and (_09513_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_09514_, _09513_, _09506_);
  or (_09515_, _09514_, _09512_);
  or (_09516_, _09515_, _09511_);
  and (_08845_, _09516_, _05552_);
  and (_09517_, _08645_, _08503_);
  not (_09518_, _09517_);
  and (_09519_, _08649_, _09297_);
  not (_09520_, _08652_);
  nor (_09521_, _09166_, _09520_);
  and (_09522_, _09521_, _09172_);
  not (_09523_, _09521_);
  and (_09524_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_09525_, _09524_, _09522_);
  nor (_09526_, _09525_, _09519_);
  and (_09527_, _09519_, word_in[8]);
  or (_09528_, _09527_, _09526_);
  and (_09529_, _09528_, _09518_);
  and (_09530_, _08665_, _08572_);
  and (_09531_, _09517_, _09311_);
  or (_09532_, _09531_, _09530_);
  or (_09533_, _09532_, _09529_);
  not (_09534_, _09530_);
  or (_09535_, _09534_, word_in[24]);
  and (_13879_, _09535_, _09533_);
  and (_09536_, _09521_, _09195_);
  and (_09537_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_09538_, _09537_, _09536_);
  nor (_09539_, _09538_, _09519_);
  and (_09540_, _09519_, word_in[9]);
  or (_09541_, _09540_, _09539_);
  and (_09542_, _09541_, _09518_);
  and (_09543_, _09517_, _09316_);
  or (_09544_, _09543_, _09530_);
  or (_09545_, _09544_, _09542_);
  or (_09546_, _09534_, word_in[25]);
  and (_08899_, _09546_, _09545_);
  and (_09547_, _09521_, _09207_);
  and (_09548_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_09549_, _09548_, _09547_);
  nor (_09550_, _09549_, _09519_);
  and (_09551_, _09519_, word_in[10]);
  or (_09552_, _09551_, _09550_);
  and (_09553_, _09552_, _09518_);
  and (_09554_, _09517_, _09335_);
  or (_09555_, _09554_, _09530_);
  or (_09556_, _09555_, _09553_);
  or (_09557_, _09534_, word_in[26]);
  and (_08902_, _09557_, _09556_);
  and (_09558_, _09521_, _09223_);
  and (_09559_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_09560_, _09559_, _09558_);
  nor (_09561_, _09560_, _09519_);
  and (_09562_, _09519_, word_in[11]);
  or (_09563_, _09562_, _09561_);
  and (_09564_, _09563_, _09518_);
  and (_09565_, _09517_, _09340_);
  or (_09566_, _09565_, _09564_);
  and (_09567_, _09566_, _09534_);
  and (_09568_, _09530_, word_in[27]);
  or (_08907_, _09568_, _09567_);
  and (_09569_, _09521_, _09241_);
  and (_09570_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_09571_, _09570_, _09569_);
  nor (_09572_, _09571_, _09519_);
  and (_09573_, _09519_, word_in[12]);
  or (_09574_, _09573_, _09572_);
  and (_09575_, _09574_, _09518_);
  and (_09576_, _09517_, _09359_);
  or (_09577_, _09576_, _09530_);
  or (_09578_, _09577_, _09575_);
  or (_09579_, _09534_, word_in[28]);
  and (_08912_, _09579_, _09578_);
  or (_09580_, _09521_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  or (_09581_, _09523_, _09253_);
  and (_09582_, _09581_, _09580_);
  or (_09583_, _09582_, _09519_);
  not (_09584_, word_in[13]);
  nand (_09585_, _09519_, _09584_);
  and (_09586_, _09585_, _09583_);
  and (_09587_, _09586_, _09518_);
  and (_09588_, _09517_, _09364_);
  or (_09589_, _09588_, _09530_);
  or (_09590_, _09589_, _09587_);
  or (_09591_, _09534_, word_in[29]);
  and (_08916_, _09591_, _09590_);
  and (_09592_, _09521_, _09269_);
  and (_09593_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_09594_, _09593_, _09592_);
  nor (_09595_, _09594_, _09519_);
  and (_09596_, _09519_, word_in[14]);
  or (_09597_, _09596_, _09595_);
  and (_09598_, _09597_, _09518_);
  and (_09599_, _09517_, _09383_);
  or (_09600_, _09599_, _09530_);
  or (_09601_, _09600_, _09598_);
  or (_09602_, _09534_, word_in[30]);
  and (_08919_, _09602_, _09601_);
  nor (_09603_, _09521_, _08336_);
  and (_09604_, _09521_, _08656_);
  or (_09605_, _09604_, _09603_);
  or (_09606_, _09605_, _09519_);
  nand (_09607_, _09519_, _09281_);
  and (_09608_, _09607_, _09606_);
  or (_09609_, _09608_, _09517_);
  or (_09610_, _09518_, _08667_);
  and (_09611_, _09610_, _09534_);
  and (_09612_, _09611_, _09609_);
  and (_09613_, _09530_, word_in[31]);
  or (_08922_, _09613_, _09612_);
  and (_09614_, _08644_, _08685_);
  not (_09615_, _09614_);
  and (_09616_, _08648_, _08696_);
  not (_09617_, _09616_);
  and (_09618_, _08653_, _08720_);
  and (_09619_, _09618_, _09165_);
  not (_09620_, _09619_);
  and (_09621_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_09622_, _09619_, word_in[0]);
  or (_09623_, _09622_, _09621_);
  and (_09624_, _09623_, _09617_);
  and (_09625_, _09616_, word_in[8]);
  or (_09626_, _09625_, _09624_);
  and (_09627_, _09626_, _09615_);
  and (_09628_, _08664_, _08561_);
  and (_09629_, _09628_, _08566_);
  and (_09630_, _09629_, _08420_);
  and (_09631_, _09614_, _09311_);
  or (_09632_, _09631_, _09630_);
  or (_09633_, _09632_, _09627_);
  not (_09634_, _09630_);
  or (_09635_, _09634_, _09189_);
  and (_09011_, _09635_, _09633_);
  and (_09636_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_09637_, _09619_, word_in[1]);
  or (_09638_, _09637_, _09636_);
  and (_09639_, _09638_, _09617_);
  and (_09640_, _09616_, word_in[9]);
  or (_09641_, _09640_, _09639_);
  or (_09642_, _09641_, _09614_);
  nor (_09643_, _09615_, _09316_);
  nor (_09644_, _09643_, _09630_);
  and (_09645_, _09644_, _09642_);
  and (_09646_, _09630_, _09191_);
  or (_09016_, _09646_, _09645_);
  and (_09647_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_09648_, _09619_, word_in[2]);
  or (_09649_, _09648_, _09647_);
  and (_09650_, _09649_, _09617_);
  and (_09651_, _09616_, word_in[10]);
  or (_09652_, _09651_, _09650_);
  and (_09653_, _09652_, _09615_);
  and (_09654_, _09614_, _09335_);
  or (_09655_, _09654_, _09630_);
  or (_09656_, _09655_, _09653_);
  or (_09657_, _09634_, _09204_);
  and (_13880_, _09657_, _09656_);
  and (_09658_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_09659_, _09619_, word_in[3]);
  or (_09660_, _09659_, _09658_);
  and (_09661_, _09660_, _09617_);
  and (_09662_, _09616_, word_in[11]);
  or (_09663_, _09662_, _09661_);
  and (_09664_, _09663_, _09615_);
  and (_09665_, _09614_, _09340_);
  or (_09666_, _09665_, _09630_);
  or (_09667_, _09666_, _09664_);
  or (_09668_, _09634_, _09218_);
  and (_13881_, _09668_, _09667_);
  and (_09669_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_09670_, _09619_, word_in[4]);
  or (_09671_, _09670_, _09669_);
  and (_09672_, _09671_, _09617_);
  and (_09673_, _09616_, word_in[12]);
  or (_09674_, _09673_, _09672_);
  and (_09675_, _09674_, _09615_);
  and (_09676_, _09614_, _09359_);
  or (_09677_, _09676_, _09630_);
  or (_09678_, _09677_, _09675_);
  or (_09679_, _09634_, _09236_);
  and (_13882_, _09679_, _09678_);
  and (_09680_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_09681_, _09619_, word_in[5]);
  or (_09682_, _09681_, _09680_);
  and (_09683_, _09682_, _09617_);
  and (_09684_, _09616_, word_in[13]);
  or (_09685_, _09684_, _09683_);
  and (_09686_, _09685_, _09615_);
  and (_09687_, _09614_, _09364_);
  or (_09688_, _09687_, _09630_);
  or (_09689_, _09688_, _09686_);
  or (_09690_, _09634_, _09251_);
  and (_13883_, _09690_, _09689_);
  and (_09691_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_09692_, _09619_, word_in[6]);
  or (_09693_, _09692_, _09691_);
  and (_09694_, _09693_, _09617_);
  and (_09695_, _09616_, word_in[14]);
  or (_09696_, _09695_, _09694_);
  and (_09697_, _09696_, _09615_);
  and (_09698_, _09614_, _09383_);
  or (_09699_, _09698_, _09630_);
  or (_09700_, _09699_, _09697_);
  or (_09701_, _09634_, _09267_);
  and (_09034_, _09701_, _09700_);
  nor (_09702_, _09619_, _08473_);
  and (_09703_, _09619_, word_in[7]);
  or (_09704_, _09703_, _09702_);
  or (_09705_, _09704_, _09616_);
  nand (_09706_, _09616_, _09281_);
  and (_09707_, _09706_, _09705_);
  or (_09708_, _09707_, _09614_);
  or (_09709_, _09615_, _08667_);
  and (_09710_, _09709_, _09708_);
  or (_09711_, _09710_, _09630_);
  or (_09712_, _09634_, _08672_);
  and (_09037_, _09712_, _09711_);
  and (_09713_, _09629_, _08390_);
  not (_09714_, _09713_);
  and (_09715_, _09294_, _08862_);
  and (_09716_, _09715_, _09311_);
  not (_09717_, _09715_);
  and (_09718_, _09298_, _08467_);
  and (_09719_, _09618_, _09300_);
  and (_09720_, _09719_, _09172_);
  not (_09721_, _09719_);
  and (_09722_, _09721_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_09723_, _09722_, _09720_);
  nor (_09724_, _09723_, _09718_);
  and (_09725_, _09718_, word_in[8]);
  or (_09726_, _09725_, _09724_);
  and (_09727_, _09726_, _09717_);
  or (_09728_, _09727_, _09716_);
  and (_09729_, _09728_, _09714_);
  and (_09730_, _09713_, word_in[24]);
  or (_09110_, _09730_, _09729_);
  and (_09731_, _09715_, _09316_);
  and (_09732_, _09719_, _09195_);
  and (_09733_, _09721_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_09734_, _09733_, _09732_);
  nor (_09735_, _09734_, _09718_);
  and (_09736_, _09718_, word_in[9]);
  or (_09737_, _09736_, _09735_);
  and (_09738_, _09737_, _09717_);
  or (_09739_, _09738_, _09731_);
  and (_09740_, _09739_, _09714_);
  and (_09741_, _09713_, word_in[25]);
  or (_09115_, _09741_, _09740_);
  or (_09742_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  or (_09743_, _09721_, _09207_);
  and (_09744_, _09743_, _09742_);
  or (_09745_, _09744_, _09718_);
  not (_09746_, _09718_);
  or (_09747_, _09746_, word_in[10]);
  and (_09748_, _09747_, _09745_);
  or (_09749_, _09748_, _09715_);
  or (_09750_, _09717_, _09335_);
  and (_09752_, _09750_, _09749_);
  or (_09753_, _09752_, _09713_);
  or (_09754_, _09714_, word_in[26]);
  and (_09120_, _09754_, _09753_);
  or (_09756_, _09717_, _09340_);
  or (_09757_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  or (_09759_, _09721_, _09223_);
  and (_09761_, _09759_, _09757_);
  or (_09763_, _09761_, _09718_);
  or (_09764_, _09746_, word_in[11]);
  and (_09766_, _09764_, _09763_);
  or (_09767_, _09766_, _09715_);
  and (_09768_, _09767_, _09756_);
  or (_09770_, _09768_, _09713_);
  or (_09771_, _09714_, word_in[27]);
  and (_09125_, _09771_, _09770_);
  and (_09773_, _09719_, _09241_);
  and (_09774_, _09721_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_09775_, _09774_, _09773_);
  nor (_09776_, _09775_, _09718_);
  and (_09777_, _09718_, word_in[12]);
  or (_09778_, _09777_, _09776_);
  and (_09779_, _09778_, _09717_);
  and (_09780_, _09715_, _09359_);
  or (_09781_, _09780_, _09713_);
  or (_09782_, _09781_, _09779_);
  or (_09783_, _09714_, word_in[28]);
  and (_09129_, _09783_, _09782_);
  or (_09784_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or (_09785_, _09721_, _09253_);
  and (_09786_, _09785_, _09784_);
  or (_09787_, _09786_, _09718_);
  nand (_09788_, _09718_, _09584_);
  and (_09789_, _09788_, _09787_);
  or (_09790_, _09789_, _09715_);
  or (_09791_, _09717_, _09364_);
  and (_09792_, _09791_, _09790_);
  or (_09793_, _09792_, _09713_);
  or (_09794_, _09714_, word_in[29]);
  and (_09134_, _09794_, _09793_);
  or (_09795_, _09717_, _09383_);
  or (_09796_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or (_09797_, _09721_, _09269_);
  and (_09798_, _09797_, _09796_);
  or (_09799_, _09798_, _09718_);
  or (_09800_, _09746_, word_in[14]);
  and (_09801_, _09800_, _09799_);
  or (_09802_, _09801_, _09715_);
  and (_09803_, _09802_, _09795_);
  or (_09804_, _09803_, _09713_);
  or (_09805_, _09714_, word_in[30]);
  and (_09138_, _09805_, _09804_);
  or (_09806_, _09717_, _08667_);
  nor (_09807_, _09719_, _08347_);
  and (_09808_, _09719_, _08656_);
  or (_09809_, _09808_, _09807_);
  or (_09810_, _09809_, _09718_);
  nand (_09811_, _09718_, _09281_);
  and (_09812_, _09811_, _09810_);
  or (_09813_, _09812_, _09715_);
  and (_09814_, _09813_, _09806_);
  or (_09815_, _09814_, _09713_);
  or (_09816_, _09714_, word_in[31]);
  and (_09141_, _09816_, _09815_);
  and (_09817_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand (_09818_, _09817_, _05556_);
  nand (_09819_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_09164_, _09819_, _09818_);
  and (_09820_, _09401_, _08862_);
  not (_09821_, _09820_);
  and (_09822_, _09405_, _08467_);
  not (_09823_, _09822_);
  and (_09824_, _09618_, _09410_);
  not (_09825_, _09824_);
  and (_09826_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_09827_, _09824_, word_in[0]);
  or (_09828_, _09827_, _09826_);
  and (_09829_, _09828_, _09823_);
  and (_09830_, _09822_, word_in[8]);
  or (_09831_, _09830_, _09829_);
  and (_09833_, _09831_, _09821_);
  and (_09834_, _09629_, _08392_);
  and (_09835_, _09820_, _09311_);
  or (_09837_, _09835_, _09834_);
  or (_09838_, _09837_, _09833_);
  not (_09839_, _09834_);
  or (_09841_, _09839_, word_in[24]);
  and (_09217_, _09841_, _09838_);
  and (_09843_, _09824_, word_in[1]);
  and (_09844_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  or (_09846_, _09844_, _09843_);
  and (_09848_, _09846_, _09823_);
  and (_09849_, _09822_, word_in[9]);
  or (_09851_, _09849_, _09848_);
  and (_09852_, _09851_, _09821_);
  and (_09853_, _09820_, _09316_);
  or (_09854_, _09853_, _09834_);
  or (_09855_, _09854_, _09852_);
  or (_09856_, _09839_, word_in[25]);
  and (_09220_, _09856_, _09855_);
  or (_09857_, _09821_, _09335_);
  or (_09858_, _09824_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  or (_09859_, _09825_, word_in[2]);
  and (_09860_, _09859_, _09858_);
  or (_09861_, _09860_, _09822_);
  or (_09862_, _09823_, word_in[10]);
  and (_09863_, _09862_, _09861_);
  or (_09864_, _09863_, _09820_);
  and (_09865_, _09864_, _09857_);
  or (_09866_, _09865_, _09834_);
  or (_09867_, _09839_, word_in[26]);
  and (_09224_, _09867_, _09866_);
  and (_09868_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_09869_, _09824_, word_in[3]);
  or (_09870_, _09869_, _09868_);
  and (_09871_, _09870_, _09823_);
  and (_09872_, _09822_, word_in[11]);
  or (_09873_, _09872_, _09871_);
  and (_09874_, _09873_, _09821_);
  and (_09875_, _09820_, _09340_);
  or (_09876_, _09875_, _09834_);
  or (_09877_, _09876_, _09874_);
  or (_09878_, _09839_, word_in[27]);
  and (_09229_, _09878_, _09877_);
  and (_09879_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_09880_, _09824_, word_in[4]);
  or (_09881_, _09880_, _09879_);
  and (_09882_, _09881_, _09823_);
  and (_09883_, _09822_, word_in[12]);
  or (_09884_, _09883_, _09882_);
  and (_09885_, _09884_, _09821_);
  and (_09886_, _09820_, _09359_);
  or (_09887_, _09886_, _09834_);
  or (_09888_, _09887_, _09885_);
  or (_09889_, _09839_, word_in[28]);
  and (_09233_, _09889_, _09888_);
  or (_09890_, _09821_, _09364_);
  and (_09891_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_09892_, _09824_, word_in[5]);
  or (_09893_, _09892_, _09891_);
  or (_09894_, _09893_, _09822_);
  nand (_09895_, _09822_, _09584_);
  and (_09896_, _09895_, _09894_);
  or (_09897_, _09896_, _09820_);
  and (_09898_, _09897_, _09890_);
  or (_09899_, _09898_, _09834_);
  or (_09900_, _09839_, word_in[29]);
  and (_09235_, _09900_, _09899_);
  and (_09901_, _09824_, word_in[6]);
  and (_09902_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or (_09903_, _09902_, _09901_);
  and (_09904_, _09903_, _09823_);
  and (_09905_, _09822_, word_in[14]);
  or (_09906_, _09905_, _09904_);
  and (_09907_, _09906_, _09821_);
  and (_09908_, _09820_, _09383_);
  or (_09909_, _09908_, _09834_);
  or (_09911_, _09909_, _09907_);
  or (_09912_, _09839_, word_in[30]);
  and (_09238_, _09912_, _09911_);
  nor (_09913_, _09824_, _08468_);
  and (_09914_, _09824_, word_in[7]);
  or (_09915_, _09914_, _09913_);
  or (_09916_, _09915_, _09822_);
  nand (_09917_, _09822_, _09281_);
  and (_09918_, _09917_, _09916_);
  and (_09919_, _09918_, _09821_);
  and (_09920_, _09820_, _08667_);
  or (_09921_, _09920_, _09834_);
  or (_09922_, _09921_, _09919_);
  or (_09924_, _09839_, word_in[31]);
  and (_09242_, _09924_, _09922_);
  and (_09927_, _08664_, _08722_);
  and (_09928_, _08649_, _08467_);
  and (_09930_, _09618_, _08652_);
  or (_09931_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  not (_09933_, _09930_);
  or (_09934_, _09933_, _09172_);
  and (_09936_, _09934_, _09931_);
  or (_09937_, _09936_, _09928_);
  not (_09938_, _09928_);
  or (_09940_, _09938_, word_in[8]);
  and (_09942_, _09940_, _09937_);
  and (_09943_, _08644_, _08498_);
  and (_09944_, _09943_, _08502_);
  and (_09945_, _09944_, _08420_);
  or (_09946_, _09945_, _09942_);
  nand (_09947_, _08862_, _08645_);
  or (_09948_, _09947_, _09311_);
  and (_09949_, _09948_, _09946_);
  or (_09950_, _09949_, _09927_);
  not (_09951_, _09927_);
  or (_09952_, _09951_, word_in[24]);
  and (_13884_, _09952_, _09950_);
  or (_09953_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  or (_09954_, _09933_, _09195_);
  and (_09955_, _09954_, _09953_);
  or (_09956_, _09955_, _09928_);
  or (_09957_, _09938_, word_in[9]);
  and (_09958_, _09957_, _09956_);
  or (_09959_, _09958_, _09945_);
  or (_09960_, _09947_, _09316_);
  and (_09961_, _09960_, _09959_);
  or (_09962_, _09961_, _09927_);
  or (_09963_, _09951_, word_in[25]);
  and (_13885_, _09963_, _09962_);
  or (_09964_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  or (_09965_, _09933_, _09207_);
  and (_09966_, _09965_, _09964_);
  or (_09967_, _09966_, _09928_);
  or (_09968_, _09938_, word_in[10]);
  and (_09969_, _09968_, _09967_);
  or (_09970_, _09969_, _09945_);
  or (_09971_, _09947_, _09335_);
  and (_09972_, _09971_, _09970_);
  or (_09973_, _09972_, _09927_);
  or (_09974_, _09951_, word_in[26]);
  and (_13886_, _09974_, _09973_);
  or (_09975_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  or (_09976_, _09933_, _09223_);
  and (_09977_, _09976_, _09975_);
  or (_09978_, _09977_, _09928_);
  or (_09979_, _09938_, word_in[11]);
  and (_09980_, _09979_, _09978_);
  or (_09981_, _09980_, _09945_);
  or (_09982_, _09947_, _09340_);
  and (_09983_, _09982_, _09981_);
  or (_09984_, _09983_, _09927_);
  or (_09985_, _09951_, word_in[27]);
  and (_13887_, _09985_, _09984_);
  and (_09986_, _09933_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_09987_, _09930_, _09241_);
  nor (_09988_, _09987_, _09986_);
  nor (_09989_, _09988_, _09928_);
  and (_09990_, _09928_, word_in[12]);
  or (_09991_, _09990_, _09989_);
  and (_09992_, _09991_, _09947_);
  and (_09993_, _09945_, _09359_);
  or (_09994_, _09993_, _09992_);
  and (_09995_, _09994_, _09951_);
  and (_09996_, _09927_, word_in[28]);
  or (_13888_, _09996_, _09995_);
  or (_09997_, _09947_, _09364_);
  or (_09998_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  or (_09999_, _09933_, _09253_);
  and (_10000_, _09999_, _09998_);
  or (_10001_, _10000_, _09928_);
  nand (_10002_, _09928_, _09584_);
  and (_10003_, _10002_, _10001_);
  or (_10004_, _10003_, _09945_);
  and (_10005_, _10004_, _09997_);
  or (_10006_, _10005_, _09927_);
  or (_10007_, _09951_, word_in[29]);
  and (_13889_, _10007_, _10006_);
  or (_10008_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  or (_10009_, _09933_, _09269_);
  and (_10010_, _10009_, _10008_);
  or (_10011_, _10010_, _09928_);
  or (_10012_, _09938_, word_in[14]);
  and (_10013_, _10012_, _10011_);
  or (_10014_, _10013_, _09945_);
  or (_10015_, _09947_, _09383_);
  and (_10016_, _10015_, _10014_);
  or (_10017_, _10016_, _09927_);
  or (_10018_, _09951_, word_in[30]);
  and (_13890_, _10018_, _10017_);
  nand (_10019_, _09928_, _09281_);
  nor (_10020_, _09930_, _08341_);
  and (_10021_, _09930_, _08656_);
  or (_10022_, _10021_, _10020_);
  nor (_10023_, _10022_, _09928_);
  nor (_10024_, _10023_, _09945_);
  and (_10025_, _10024_, _10019_);
  and (_10026_, _09945_, _08667_);
  or (_10027_, _10026_, _10025_);
  and (_10028_, _10027_, _09951_);
  and (_10029_, _09927_, word_in[31]);
  or (_13891_, _10029_, _10028_);
  and (_10030_, _08664_, _08741_);
  not (_10031_, _10030_);
  and (_10032_, _08644_, _08765_);
  and (_10034_, _10032_, word_in[16]);
  not (_10035_, _10032_);
  and (_10036_, _08648_, _08398_);
  not (_10037_, _10036_);
  and (_10038_, _08653_, _08961_);
  and (_10039_, _10038_, _09165_);
  and (_10040_, _10039_, word_in[0]);
  not (_10041_, _10039_);
  and (_10042_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or (_10043_, _10042_, _10040_);
  and (_10044_, _10043_, _10037_);
  and (_10045_, _10036_, word_in[8]);
  or (_10046_, _10045_, _10044_);
  and (_10047_, _10046_, _10035_);
  or (_10048_, _10047_, _10034_);
  and (_10049_, _10048_, _10031_);
  and (_10050_, _10030_, word_in[24]);
  or (_09403_, _10050_, _10049_);
  and (_10051_, _10032_, word_in[17]);
  and (_10052_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_10053_, _10039_, word_in[1]);
  or (_10054_, _10053_, _10052_);
  and (_10055_, _10054_, _10037_);
  and (_10056_, _10036_, word_in[9]);
  or (_10057_, _10056_, _10055_);
  and (_10058_, _10057_, _10035_);
  or (_10059_, _10058_, _10051_);
  and (_10060_, _10059_, _10031_);
  and (_10061_, _10030_, word_in[25]);
  or (_09408_, _10061_, _10060_);
  and (_10062_, _10032_, word_in[18]);
  and (_10063_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_10064_, _10039_, word_in[2]);
  or (_10065_, _10064_, _10063_);
  and (_10066_, _10065_, _10037_);
  and (_10067_, _10036_, word_in[10]);
  or (_10068_, _10067_, _10066_);
  and (_10069_, _10068_, _10035_);
  or (_10070_, _10069_, _10062_);
  and (_10071_, _10070_, _10031_);
  and (_10072_, _10030_, word_in[26]);
  or (_13892_, _10072_, _10071_);
  and (_10073_, _10032_, word_in[19]);
  and (_10074_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_10075_, _10039_, word_in[3]);
  or (_10076_, _10075_, _10074_);
  and (_10077_, _10076_, _10037_);
  and (_10078_, _10036_, word_in[11]);
  or (_10079_, _10078_, _10077_);
  and (_10080_, _10079_, _10035_);
  or (_10081_, _10080_, _10073_);
  and (_10082_, _10081_, _10031_);
  and (_10083_, _10030_, word_in[27]);
  or (_13893_, _10083_, _10082_);
  and (_10084_, _10032_, word_in[20]);
  and (_10085_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_10086_, _10039_, word_in[4]);
  or (_10087_, _10086_, _10085_);
  and (_10088_, _10087_, _10037_);
  and (_10090_, _10036_, word_in[12]);
  or (_10091_, _10090_, _10088_);
  and (_10092_, _10091_, _10035_);
  or (_10093_, _10092_, _10084_);
  and (_10094_, _10093_, _10031_);
  and (_10095_, _10030_, word_in[28]);
  or (_13894_, _10095_, _10094_);
  and (_10096_, _10032_, word_in[21]);
  and (_10097_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_10098_, _10039_, word_in[5]);
  or (_10099_, _10098_, _10097_);
  and (_10100_, _10099_, _10037_);
  and (_10101_, _10036_, word_in[13]);
  or (_10102_, _10101_, _10100_);
  and (_10103_, _10102_, _10035_);
  or (_10104_, _10103_, _10096_);
  and (_10105_, _10104_, _10031_);
  and (_10106_, _10030_, word_in[29]);
  or (_13895_, _10106_, _10105_);
  and (_10107_, _10032_, word_in[22]);
  and (_10108_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_10109_, _10039_, word_in[6]);
  or (_10110_, _10109_, _10108_);
  and (_10111_, _10110_, _10037_);
  and (_10112_, _10036_, word_in[14]);
  or (_10113_, _10112_, _10111_);
  and (_10114_, _10113_, _10035_);
  or (_10115_, _10114_, _10107_);
  and (_10116_, _10115_, _10031_);
  and (_10117_, _10030_, word_in[30]);
  or (_13896_, _10117_, _10116_);
  nor (_10118_, _10039_, _08448_);
  and (_10120_, _10039_, word_in[7]);
  or (_10121_, _10120_, _10118_);
  and (_10122_, _10121_, _10037_);
  and (_10123_, _10036_, word_in[15]);
  or (_10124_, _10123_, _10122_);
  and (_10125_, _10124_, _10035_);
  and (_10126_, _10032_, word_in[23]);
  or (_10127_, _10126_, _10125_);
  and (_10128_, _10127_, _10031_);
  and (_10129_, _10030_, word_in[31]);
  or (_13897_, _10129_, _10128_);
  and (_10130_, _09294_, _08507_);
  and (_10131_, _09298_, _08402_);
  and (_10132_, _10038_, _09300_);
  or (_10133_, _10132_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  not (_10134_, _10132_);
  or (_10135_, _10134_, word_in[0]);
  and (_10136_, _10135_, _10133_);
  or (_10137_, _10136_, _10131_);
  not (_10138_, _10131_);
  or (_10139_, _10138_, word_in[8]);
  and (_10140_, _10139_, _10137_);
  or (_10141_, _10140_, _10130_);
  and (_10142_, _08664_, _08567_);
  and (_10143_, _10142_, _08390_);
  not (_10144_, _10143_);
  not (_10145_, _10130_);
  or (_10146_, _10145_, _09311_);
  and (_10147_, _10146_, _10144_);
  and (_10148_, _10147_, _10141_);
  and (_10149_, _10143_, word_in[24]);
  or (_13898_, _10149_, _10148_);
  and (_10150_, _10130_, _09316_);
  and (_10151_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_10152_, _10132_, word_in[1]);
  nor (_10153_, _10152_, _10151_);
  nor (_10154_, _10153_, _10131_);
  and (_10155_, _10131_, word_in[9]);
  or (_10156_, _10155_, _10154_);
  and (_10157_, _10156_, _10145_);
  or (_10158_, _10157_, _10150_);
  and (_10159_, _10158_, _10144_);
  and (_10160_, _10143_, word_in[25]);
  or (_13899_, _10160_, _10159_);
  and (_10161_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_10162_, _10132_, word_in[2]);
  nor (_10163_, _10162_, _10161_);
  nor (_10164_, _10163_, _10131_);
  and (_10165_, _10131_, word_in[10]);
  or (_10166_, _10165_, _10164_);
  and (_10167_, _10166_, _10145_);
  and (_10168_, _10130_, _09335_);
  or (_10169_, _10168_, _10167_);
  and (_10170_, _10169_, _10144_);
  and (_10171_, _10143_, word_in[26]);
  or (_13900_, _10171_, _10170_);
  and (_10172_, _10132_, word_in[3]);
  and (_10173_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_10174_, _10173_, _10172_);
  nor (_10175_, _10174_, _10131_);
  and (_10176_, _10131_, word_in[11]);
  or (_10177_, _10176_, _10175_);
  and (_10178_, _10177_, _10145_);
  and (_10179_, _10130_, _09340_);
  or (_10180_, _10179_, _10143_);
  or (_10181_, _10180_, _10178_);
  or (_10182_, _10144_, word_in[27]);
  and (_13901_, _10182_, _10181_);
  and (_10183_, _10132_, word_in[4]);
  and (_10184_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_10185_, _10184_, _10183_);
  nor (_10186_, _10185_, _10131_);
  and (_10187_, _10131_, word_in[12]);
  or (_10188_, _10187_, _10186_);
  and (_10189_, _10188_, _10145_);
  and (_10190_, _10130_, _09359_);
  or (_10191_, _10190_, _10189_);
  and (_10192_, _10191_, _10144_);
  and (_10193_, _10143_, word_in[28]);
  or (_13902_, _10193_, _10192_);
  and (_10194_, _10132_, word_in[5]);
  and (_10195_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_10196_, _10195_, _10194_);
  nor (_10197_, _10196_, _10131_);
  and (_10198_, _10131_, word_in[13]);
  or (_10199_, _10198_, _10197_);
  and (_10200_, _10199_, _10145_);
  and (_10201_, _10130_, _09364_);
  or (_10202_, _10201_, _10200_);
  and (_10203_, _10202_, _10144_);
  and (_10204_, _10143_, word_in[29]);
  or (_13903_, _10204_, _10203_);
  or (_10205_, _10132_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or (_10206_, _10134_, word_in[6]);
  and (_10207_, _10206_, _10205_);
  or (_10208_, _10207_, _10131_);
  or (_10209_, _10138_, word_in[14]);
  and (_10210_, _10209_, _10208_);
  or (_10211_, _10210_, _10130_);
  or (_10212_, _10145_, _09383_);
  and (_10213_, _10212_, _10144_);
  and (_10214_, _10213_, _10211_);
  and (_10215_, _10143_, word_in[30]);
  or (_13904_, _10215_, _10214_);
  and (_10216_, _10132_, word_in[7]);
  nor (_10217_, _10132_, _08328_);
  nor (_10218_, _10217_, _10216_);
  nor (_10219_, _10218_, _10131_);
  and (_10220_, _10131_, word_in[15]);
  or (_10221_, _10220_, _10219_);
  and (_10222_, _10221_, _10145_);
  and (_10223_, _10130_, _08667_);
  or (_10224_, _10223_, _10222_);
  and (_10225_, _10224_, _10144_);
  and (_10226_, _10143_, word_in[31]);
  or (_13905_, _10226_, _10225_);
  and (_10227_, _09401_, _08507_);
  and (_10228_, _09405_, _08402_);
  and (_10229_, _09410_, _08961_);
  not (_10230_, _10229_);
  and (_10231_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_10232_, _10229_, word_in[0]);
  or (_10233_, _10232_, _10231_);
  or (_10234_, _10233_, _10228_);
  not (_10235_, _10228_);
  or (_10236_, _10235_, word_in[8]);
  and (_10237_, _10236_, _10234_);
  or (_10238_, _10237_, _10227_);
  and (_10239_, _10142_, _08392_);
  not (_10240_, _10239_);
  not (_10241_, _10227_);
  or (_10242_, _10241_, _09311_);
  and (_10243_, _10242_, _10240_);
  and (_10244_, _10243_, _10238_);
  and (_10245_, _10239_, word_in[24]);
  or (_13853_, _10245_, _10244_);
  or (_10246_, _10229_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  or (_10248_, _10230_, word_in[1]);
  and (_10249_, _10248_, _10246_);
  or (_10250_, _10249_, _10228_);
  or (_10251_, _10235_, word_in[9]);
  and (_10252_, _10251_, _10250_);
  or (_10253_, _10252_, _10227_);
  or (_10255_, _10241_, _09316_);
  and (_10256_, _10255_, _10253_);
  and (_10258_, _10256_, _10240_);
  and (_10259_, _10239_, word_in[25]);
  or (_13854_, _10259_, _10258_);
  or (_10260_, _10229_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  or (_10261_, _10230_, word_in[2]);
  and (_10262_, _10261_, _10260_);
  or (_10264_, _10262_, _10228_);
  or (_10265_, _10235_, word_in[10]);
  and (_10266_, _10265_, _10264_);
  or (_10267_, _10266_, _10227_);
  or (_10268_, _10241_, _09335_);
  and (_10270_, _10268_, _10240_);
  and (_10271_, _10270_, _10267_);
  and (_10272_, _10239_, word_in[26]);
  or (_13855_, _10272_, _10271_);
  and (_10273_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_10274_, _10229_, word_in[3]);
  or (_10275_, _10274_, _10273_);
  or (_10276_, _10275_, _10228_);
  or (_10277_, _10235_, word_in[11]);
  and (_10278_, _10277_, _10276_);
  or (_10279_, _10278_, _10227_);
  or (_10280_, _10241_, _09340_);
  and (_10281_, _10280_, _10240_);
  and (_10283_, _10281_, _10279_);
  and (_10284_, _10239_, word_in[27]);
  or (_13856_, _10284_, _10283_);
  and (_10285_, _10227_, _09359_);
  and (_10286_, _10229_, word_in[4]);
  and (_10287_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  or (_10288_, _10287_, _10286_);
  or (_10289_, _10288_, _10228_);
  or (_10290_, _10235_, word_in[12]);
  and (_10291_, _10290_, _10241_);
  and (_10292_, _10291_, _10289_);
  or (_10293_, _10292_, _10285_);
  and (_10294_, _10293_, _10240_);
  and (_10295_, _10239_, word_in[28]);
  or (_13857_, _10295_, _10294_);
  and (_10296_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_10297_, _10229_, word_in[5]);
  or (_10299_, _10297_, _10296_);
  or (_10300_, _10299_, _10228_);
  nand (_10301_, _10228_, _09584_);
  and (_10303_, _10301_, _10300_);
  or (_10304_, _10303_, _10227_);
  or (_10305_, _10241_, _09364_);
  and (_10306_, _10305_, _10240_);
  and (_10307_, _10306_, _10304_);
  and (_10308_, _10239_, word_in[29]);
  or (_13858_, _10308_, _10307_);
  or (_10309_, _10229_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or (_10310_, _10230_, word_in[6]);
  and (_10311_, _10310_, _10309_);
  or (_10312_, _10311_, _10228_);
  or (_10313_, _10235_, word_in[14]);
  and (_10314_, _10313_, _10312_);
  or (_10315_, _10314_, _10227_);
  or (_10316_, _10241_, _09383_);
  and (_10317_, _10316_, _10240_);
  and (_10318_, _10317_, _10315_);
  and (_10319_, _10239_, word_in[30]);
  or (_13859_, _10319_, _10318_);
  nor (_10320_, _10229_, _08442_);
  and (_10321_, _10229_, word_in[7]);
  or (_10322_, _10321_, _10320_);
  or (_10323_, _10322_, _10228_);
  nand (_10324_, _10228_, _09281_);
  and (_10325_, _10324_, _10323_);
  or (_10326_, _10325_, _10227_);
  or (_10327_, _10241_, _08667_);
  and (_10328_, _10327_, _10240_);
  and (_10329_, _10328_, _10326_);
  and (_10330_, _10239_, word_in[31]);
  or (_13860_, _10330_, _10329_);
  and (_10331_, _08645_, _08507_);
  not (_10332_, _10331_);
  and (_10333_, _08649_, _08402_);
  and (_10334_, _10038_, _08652_);
  and (_10335_, _10334_, word_in[0]);
  not (_10336_, _10334_);
  and (_10337_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_10338_, _10337_, _10335_);
  nor (_10339_, _10338_, _10333_);
  and (_10340_, _10333_, word_in[8]);
  or (_10341_, _10340_, _10339_);
  and (_10342_, _10341_, _10332_);
  and (_10343_, _10142_, _08429_);
  and (_10344_, _10331_, _09311_);
  or (_10345_, _10344_, _10343_);
  or (_10346_, _10345_, _10342_);
  not (_10347_, _10343_);
  or (_10348_, _10347_, _09189_);
  and (_13861_, _10348_, _10346_);
  and (_10349_, _10334_, word_in[1]);
  and (_10350_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_10351_, _10350_, _10349_);
  nor (_10352_, _10351_, _10333_);
  and (_10353_, _10333_, word_in[9]);
  or (_10354_, _10353_, _10352_);
  and (_10355_, _10354_, _10332_);
  and (_10356_, _10331_, _09316_);
  or (_10357_, _10356_, _10343_);
  or (_10358_, _10357_, _10355_);
  or (_10359_, _10347_, _09191_);
  and (_13862_, _10359_, _10358_);
  and (_10360_, _10331_, _09335_);
  and (_10362_, _10334_, word_in[2]);
  and (_10363_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_10364_, _10363_, _10362_);
  nor (_10365_, _10364_, _10333_);
  and (_10366_, _10333_, word_in[10]);
  or (_10367_, _10366_, _10365_);
  and (_10368_, _10367_, _10332_);
  or (_10369_, _10368_, _10360_);
  and (_10370_, _10369_, _10347_);
  and (_10371_, _10343_, word_in[26]);
  or (_13863_, _10371_, _10370_);
  or (_10372_, _10334_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  or (_10373_, _10336_, word_in[3]);
  and (_10374_, _10373_, _10372_);
  or (_10375_, _10374_, _10333_);
  not (_10376_, word_in[11]);
  nand (_10377_, _10333_, _10376_);
  and (_10378_, _10377_, _10375_);
  or (_10379_, _10378_, _10331_);
  or (_10380_, _10332_, _09340_);
  and (_10381_, _10380_, _10347_);
  and (_10382_, _10381_, _10379_);
  and (_10383_, _10343_, _09218_);
  or (_13864_, _10383_, _10382_);
  and (_10384_, _10334_, word_in[4]);
  and (_10385_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_10386_, _10385_, _10384_);
  nor (_10387_, _10386_, _10333_);
  and (_10388_, _10333_, word_in[12]);
  or (_10389_, _10388_, _10387_);
  and (_10390_, _10389_, _10332_);
  and (_10391_, _10331_, _09359_);
  or (_10392_, _10391_, _10390_);
  and (_10393_, _10392_, _10347_);
  and (_10394_, _10343_, word_in[28]);
  or (_13865_, _10394_, _10393_);
  and (_10395_, _10334_, word_in[5]);
  and (_10396_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_10397_, _10396_, _10395_);
  nor (_10398_, _10397_, _10333_);
  and (_10399_, _10333_, word_in[13]);
  or (_10400_, _10399_, _10398_);
  and (_10401_, _10400_, _10332_);
  and (_10402_, _10331_, _09364_);
  or (_10403_, _10402_, _10343_);
  or (_10404_, _10403_, _10401_);
  or (_10405_, _10347_, _09251_);
  and (_13866_, _10405_, _10404_);
  and (_10406_, _10334_, word_in[6]);
  and (_10407_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_10408_, _10407_, _10406_);
  nor (_10409_, _10408_, _10333_);
  and (_10410_, _10333_, word_in[14]);
  or (_10411_, _10410_, _10409_);
  and (_10412_, _10411_, _10332_);
  and (_10413_, _10331_, _09383_);
  or (_10414_, _10413_, _10412_);
  and (_10415_, _10414_, _10347_);
  and (_10416_, _10343_, word_in[30]);
  or (_13867_, _10416_, _10415_);
  and (_10417_, _10334_, word_in[7]);
  nor (_10418_, _10334_, _08317_);
  nor (_10419_, _10418_, _10417_);
  nor (_10420_, _10419_, _10333_);
  and (_10421_, _10333_, word_in[15]);
  or (_10422_, _10421_, _10420_);
  and (_10423_, _10422_, _10332_);
  and (_10424_, _10331_, _08667_);
  or (_10425_, _10424_, _10343_);
  or (_10426_, _10425_, _10423_);
  or (_10427_, _10347_, _08672_);
  and (_13868_, _10427_, _10426_);
  and (_10428_, _08644_, _08849_);
  not (_10429_, _10428_);
  and (_10430_, _08613_, _08392_);
  and (_10431_, _08648_, _10430_);
  not (_10432_, _10431_);
  and (_10433_, _09165_, _08654_);
  and (_10434_, _10433_, word_in[0]);
  not (_10435_, _10433_);
  and (_10436_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or (_10437_, _10436_, _10434_);
  and (_10438_, _10437_, _10432_);
  and (_10439_, _10431_, word_in[8]);
  or (_10440_, _10439_, _10438_);
  and (_10441_, _10440_, _10429_);
  not (_10442_, _08566_);
  and (_10443_, _09628_, _10442_);
  and (_10444_, _10443_, _08420_);
  and (_10445_, _10428_, word_in[16]);
  or (_10446_, _10445_, _10444_);
  or (_10447_, _10446_, _10441_);
  not (_10448_, _10444_);
  or (_10449_, _10448_, _09189_);
  and (_09751_, _10449_, _10447_);
  and (_10450_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_10451_, _10433_, word_in[1]);
  or (_10452_, _10451_, _10450_);
  and (_10453_, _10452_, _10432_);
  and (_10454_, _10431_, word_in[9]);
  or (_10455_, _10454_, _10453_);
  and (_10456_, _10455_, _10429_);
  and (_10457_, _10428_, word_in[17]);
  or (_10458_, _10457_, _10444_);
  or (_10459_, _10458_, _10456_);
  or (_10460_, _10448_, _09191_);
  and (_09755_, _10460_, _10459_);
  and (_10461_, _10433_, word_in[2]);
  and (_10462_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  or (_10463_, _10462_, _10461_);
  and (_10464_, _10463_, _10432_);
  and (_10465_, _10431_, word_in[10]);
  or (_10466_, _10465_, _10464_);
  and (_10467_, _10466_, _10429_);
  and (_10468_, _10428_, word_in[18]);
  or (_10469_, _10468_, _10444_);
  or (_10470_, _10469_, _10467_);
  or (_10471_, _10448_, _09204_);
  and (_09758_, _10471_, _10470_);
  and (_10472_, _10433_, word_in[3]);
  and (_10473_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  or (_10474_, _10473_, _10472_);
  and (_10475_, _10474_, _10432_);
  and (_10476_, _10431_, word_in[11]);
  or (_10477_, _10476_, _10475_);
  and (_10478_, _10477_, _10429_);
  and (_10479_, _10428_, word_in[19]);
  or (_10480_, _10479_, _10444_);
  or (_10481_, _10480_, _10478_);
  or (_10482_, _10448_, _09218_);
  and (_09760_, _10482_, _10481_);
  and (_10483_, _10433_, word_in[4]);
  and (_10484_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or (_10485_, _10484_, _10483_);
  and (_10486_, _10485_, _10432_);
  and (_10487_, _10431_, word_in[12]);
  or (_10488_, _10487_, _10486_);
  and (_10489_, _10488_, _10429_);
  and (_10490_, _10428_, word_in[20]);
  or (_10491_, _10490_, _10444_);
  or (_10492_, _10491_, _10489_);
  or (_10493_, _10448_, _09236_);
  and (_09762_, _10493_, _10492_);
  and (_10494_, _10433_, word_in[5]);
  and (_10495_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  or (_10496_, _10495_, _10494_);
  and (_10497_, _10496_, _10432_);
  and (_10498_, _10431_, word_in[13]);
  or (_10499_, _10498_, _10497_);
  and (_10500_, _10499_, _10429_);
  and (_10501_, _10428_, word_in[21]);
  or (_10502_, _10501_, _10444_);
  or (_10503_, _10502_, _10500_);
  or (_10504_, _10448_, _09251_);
  and (_09765_, _10504_, _10503_);
  and (_10505_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_10506_, _10433_, word_in[6]);
  or (_10507_, _10506_, _10505_);
  and (_10508_, _10507_, _10432_);
  and (_10509_, _10431_, word_in[14]);
  or (_10510_, _10509_, _10508_);
  and (_10511_, _10510_, _10429_);
  and (_10512_, _10428_, word_in[22]);
  or (_10513_, _10512_, _10444_);
  or (_10514_, _10513_, _10511_);
  or (_10515_, _10448_, _09267_);
  and (_09769_, _10515_, _10514_);
  nor (_10516_, _10433_, _08486_);
  and (_10517_, _10433_, word_in[7]);
  or (_10518_, _10517_, _10516_);
  and (_10519_, _10518_, _10432_);
  and (_10520_, _10431_, word_in[15]);
  or (_10521_, _10520_, _10519_);
  and (_10522_, _10521_, _10429_);
  and (_10523_, _10428_, word_in[23]);
  or (_10524_, _10523_, _10444_);
  or (_10525_, _10524_, _10522_);
  or (_10526_, _10448_, _08672_);
  and (_09772_, _10526_, _10525_);
  and (_10527_, _10443_, _08390_);
  and (_10528_, _09294_, _08643_);
  not (_10529_, _10528_);
  or (_10530_, _10529_, _09311_);
  and (_10531_, _09298_, _08480_);
  and (_10532_, _09300_, _08654_);
  not (_10533_, _10532_);
  and (_10534_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_10535_, _10532_, word_in[0]);
  or (_10536_, _10535_, _10534_);
  or (_10537_, _10536_, _10531_);
  not (_10538_, _10531_);
  or (_10539_, _10538_, word_in[8]);
  and (_10540_, _10539_, _10537_);
  or (_10541_, _10540_, _10528_);
  and (_10542_, _10541_, _10530_);
  or (_10543_, _10542_, _10527_);
  not (_10544_, _10527_);
  or (_10545_, _10544_, word_in[24]);
  and (_13869_, _10545_, _10543_);
  or (_10546_, _10529_, _09316_);
  or (_10547_, _10532_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  or (_10548_, _10533_, word_in[1]);
  and (_10549_, _10548_, _10547_);
  or (_10550_, _10549_, _10531_);
  or (_10551_, _10538_, word_in[9]);
  and (_10552_, _10551_, _10550_);
  or (_10553_, _10552_, _10528_);
  and (_10554_, _10553_, _10546_);
  or (_10555_, _10554_, _10527_);
  or (_10556_, _10544_, word_in[25]);
  and (_09832_, _10556_, _10555_);
  or (_10557_, _10529_, _09335_);
  or (_10558_, _10532_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  or (_10559_, _10533_, word_in[2]);
  and (_10560_, _10559_, _10558_);
  or (_10561_, _10560_, _10531_);
  or (_10562_, _10538_, word_in[10]);
  and (_10563_, _10562_, _10561_);
  or (_10564_, _10563_, _10528_);
  and (_10565_, _10564_, _10557_);
  or (_10566_, _10565_, _10527_);
  or (_10567_, _10544_, word_in[26]);
  and (_09836_, _10567_, _10566_);
  and (_10568_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_10569_, _10532_, word_in[3]);
  nor (_10570_, _10569_, _10568_);
  nor (_10571_, _10570_, _10531_);
  and (_10572_, _10531_, word_in[11]);
  or (_10573_, _10572_, _10571_);
  and (_10574_, _10573_, _10529_);
  and (_10575_, _10528_, _09340_);
  or (_10576_, _10575_, _10527_);
  or (_10577_, _10576_, _10574_);
  or (_10578_, _10544_, word_in[27]);
  and (_09840_, _10578_, _10577_);
  and (_10579_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_10580_, _10532_, word_in[4]);
  nor (_10581_, _10580_, _10579_);
  nor (_10582_, _10581_, _10531_);
  and (_10583_, _10531_, word_in[12]);
  or (_10584_, _10583_, _10582_);
  and (_10585_, _10584_, _10529_);
  and (_10586_, _10528_, _09359_);
  or (_10587_, _10586_, _10527_);
  or (_10588_, _10587_, _10585_);
  or (_10589_, _10544_, word_in[28]);
  and (_09842_, _10589_, _10588_);
  and (_10590_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_10591_, _10532_, word_in[5]);
  nor (_10592_, _10591_, _10590_);
  nor (_10593_, _10592_, _10531_);
  and (_10594_, _10531_, word_in[13]);
  or (_10595_, _10594_, _10593_);
  and (_10596_, _10595_, _10529_);
  and (_10597_, _10528_, _09364_);
  or (_10598_, _10597_, _10527_);
  or (_10599_, _10598_, _10596_);
  or (_10600_, _10544_, word_in[29]);
  and (_09845_, _10600_, _10599_);
  and (_10601_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_10602_, _10532_, word_in[6]);
  nor (_10603_, _10602_, _10601_);
  nor (_10605_, _10603_, _10531_);
  and (_10606_, _10531_, word_in[14]);
  or (_10607_, _10606_, _10605_);
  and (_10608_, _10607_, _10529_);
  and (_10609_, _10528_, _09383_);
  or (_10610_, _10609_, _10527_);
  or (_10611_, _10610_, _10608_);
  or (_10612_, _10544_, word_in[30]);
  and (_09847_, _10612_, _10611_);
  nor (_10613_, _10532_, _08323_);
  and (_10614_, _10532_, word_in[7]);
  nor (_10615_, _10614_, _10613_);
  nor (_10616_, _10615_, _10531_);
  and (_10617_, _10531_, word_in[15]);
  or (_10618_, _10617_, _10616_);
  and (_10619_, _10618_, _10529_);
  and (_10620_, _10528_, _08667_);
  or (_10621_, _10620_, _10527_);
  or (_10622_, _10621_, _10619_);
  or (_10624_, _10544_, word_in[31]);
  and (_09850_, _10624_, _10622_);
  and (_10626_, _08007_, _06766_);
  and (_10627_, _08989_, _08013_);
  and (_10629_, _10627_, _10626_);
  nand (_10630_, _10629_, _06811_);
  and (_10632_, _06770_, _06054_);
  and (_10633_, _08989_, _10632_);
  and (_10635_, _10633_, _10626_);
  not (_10636_, _10635_);
  and (_10638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_10639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_10641_, _10639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_10642_, _10641_, _10638_);
  not (_10643_, _10642_);
  and (_10644_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_10645_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_10646_, _10645_, _10644_);
  or (_10647_, _10629_, _10646_);
  and (_10648_, _10647_, _10636_);
  and (_10649_, _10648_, _10630_);
  and (_10650_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_10651_, _10650_, _10649_);
  and (_09910_, _10651_, _05552_);
  and (_10652_, _09401_, _08643_);
  not (_10653_, _10652_);
  and (_10654_, _09405_, _08480_);
  not (_10655_, _10654_);
  and (_10656_, _09410_, _08654_);
  not (_10657_, _10656_);
  and (_10658_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_10659_, _10656_, word_in[0]);
  or (_10660_, _10659_, _10658_);
  and (_10661_, _10660_, _10655_);
  and (_10662_, _10654_, word_in[8]);
  or (_10663_, _10662_, _10661_);
  and (_10664_, _10663_, _10653_);
  and (_10665_, _10443_, _08392_);
  and (_10666_, _10652_, _09311_);
  or (_10667_, _10666_, _10665_);
  or (_10668_, _10667_, _10664_);
  not (_10669_, _10665_);
  or (_10670_, _10669_, word_in[24]);
  and (_09923_, _10670_, _10668_);
  and (_10671_, _10656_, word_in[1]);
  and (_10672_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  or (_10673_, _10672_, _10671_);
  and (_10674_, _10673_, _10655_);
  and (_10675_, _10654_, word_in[9]);
  or (_10676_, _10675_, _10674_);
  and (_10677_, _10676_, _10653_);
  and (_10678_, _10652_, _09316_);
  or (_10679_, _10678_, _10665_);
  or (_10680_, _10679_, _10677_);
  or (_10681_, _10669_, word_in[25]);
  and (_09925_, _10681_, _10680_);
  and (_10682_, _10656_, word_in[2]);
  and (_10683_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  or (_10684_, _10683_, _10682_);
  and (_10685_, _10684_, _10655_);
  and (_10686_, _10654_, word_in[10]);
  or (_10687_, _10686_, _10685_);
  and (_10688_, _10687_, _10653_);
  and (_10689_, _10652_, _09335_);
  or (_10690_, _10689_, _10688_);
  and (_10691_, _10690_, _10669_);
  and (_10692_, _10665_, word_in[26]);
  or (_09926_, _10692_, _10691_);
  and (_10694_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_10696_, _10656_, word_in[3]);
  or (_10697_, _10696_, _10694_);
  and (_10698_, _10697_, _10655_);
  and (_10699_, _10654_, word_in[11]);
  or (_10700_, _10699_, _10698_);
  and (_10701_, _10700_, _10653_);
  and (_10702_, _10652_, _09340_);
  or (_10703_, _10702_, _10665_);
  or (_10704_, _10703_, _10701_);
  or (_10705_, _10669_, word_in[27]);
  and (_09929_, _10705_, _10704_);
  and (_10706_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_10707_, _10656_, word_in[4]);
  or (_10708_, _10707_, _10706_);
  and (_10709_, _10708_, _10655_);
  and (_10710_, _10654_, word_in[12]);
  or (_10711_, _10710_, _10709_);
  and (_10712_, _10711_, _10653_);
  and (_10713_, _10652_, _09359_);
  or (_10714_, _10713_, _10665_);
  or (_10715_, _10714_, _10712_);
  or (_10716_, _10669_, word_in[28]);
  and (_09932_, _10716_, _10715_);
  or (_10717_, _10653_, _09364_);
  or (_10718_, _10656_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  or (_10719_, _10657_, word_in[5]);
  and (_10720_, _10719_, _10718_);
  or (_10721_, _10720_, _10654_);
  nand (_10722_, _10654_, _09584_);
  and (_10723_, _10722_, _10721_);
  or (_10724_, _10723_, _10652_);
  and (_10725_, _10724_, _10717_);
  or (_10726_, _10725_, _10665_);
  or (_10727_, _10669_, word_in[29]);
  and (_09935_, _10727_, _10726_);
  and (_10728_, _10656_, word_in[6]);
  and (_10729_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or (_10730_, _10729_, _10728_);
  and (_10732_, _10730_, _10655_);
  and (_10733_, _10654_, word_in[14]);
  or (_10734_, _10733_, _10732_);
  and (_10735_, _10734_, _10653_);
  and (_10736_, _10652_, _09383_);
  or (_10737_, _10736_, _10665_);
  or (_10738_, _10737_, _10735_);
  or (_10739_, _10669_, word_in[30]);
  and (_09939_, _10739_, _10738_);
  nor (_10740_, _10656_, _08481_);
  and (_10741_, _10656_, word_in[7]);
  or (_10742_, _10741_, _10740_);
  or (_10743_, _10742_, _10654_);
  nand (_10744_, _10654_, _09281_);
  and (_10745_, _10744_, _10743_);
  or (_10746_, _10745_, _10652_);
  or (_10747_, _10653_, _08667_);
  and (_10748_, _10747_, _10746_);
  or (_10749_, _10748_, _10665_);
  or (_10750_, _10669_, word_in[31]);
  and (_09941_, _10750_, _10749_);
  not (_10751_, _08655_);
  and (_10752_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_10753_, _08655_, word_in[0]);
  nor (_10754_, _10753_, _10752_);
  nor (_10755_, _10754_, _08650_);
  and (_10756_, _08650_, word_in[8]);
  or (_10757_, _10756_, _10755_);
  and (_10758_, _10757_, _08647_);
  and (_10759_, _09311_, _08646_);
  or (_10760_, _10759_, _08666_);
  or (_10761_, _10760_, _10758_);
  or (_10762_, _08671_, word_in[24]);
  and (_13870_, _10762_, _10761_);
  and (_10763_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_10764_, _08655_, word_in[1]);
  nor (_10765_, _10764_, _10763_);
  nor (_10766_, _10765_, _08650_);
  and (_10767_, _08650_, word_in[9]);
  or (_10768_, _10767_, _10766_);
  and (_10769_, _10768_, _08647_);
  and (_10770_, _09316_, _08646_);
  or (_10771_, _10770_, _08666_);
  or (_10772_, _10771_, _10769_);
  or (_10773_, _08671_, word_in[25]);
  and (_13871_, _10773_, _10772_);
  and (_10774_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_10775_, _08655_, word_in[2]);
  nor (_10776_, _10775_, _10774_);
  nor (_10777_, _10776_, _08650_);
  and (_10778_, _08650_, word_in[10]);
  or (_10779_, _10778_, _10777_);
  and (_10780_, _10779_, _08647_);
  and (_10781_, _09335_, _08646_);
  or (_10782_, _10781_, _08666_);
  or (_10783_, _10782_, _10780_);
  or (_10784_, _08671_, word_in[26]);
  and (_13872_, _10784_, _10783_);
  and (_10785_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_10786_, _08655_, word_in[3]);
  nor (_10787_, _10786_, _10785_);
  nor (_10788_, _10787_, _08650_);
  and (_10789_, _08650_, word_in[11]);
  or (_10790_, _10789_, _10788_);
  and (_10791_, _10790_, _08647_);
  and (_10792_, _09340_, _08646_);
  or (_10793_, _10792_, _08666_);
  or (_10794_, _10793_, _10791_);
  or (_10795_, _08671_, word_in[27]);
  and (_13873_, _10795_, _10794_);
  and (_10796_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_10797_, _08655_, word_in[4]);
  nor (_10798_, _10797_, _10796_);
  nor (_10799_, _10798_, _08650_);
  and (_10800_, _08650_, word_in[12]);
  or (_10801_, _10800_, _10799_);
  and (_10802_, _10801_, _08647_);
  and (_10803_, _09359_, _08646_);
  or (_10804_, _10803_, _08666_);
  or (_10805_, _10804_, _10802_);
  or (_10806_, _08671_, word_in[28]);
  and (_13874_, _10806_, _10805_);
  or (_10808_, _09364_, _08647_);
  or (_10809_, _08655_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  or (_10811_, _10751_, word_in[5]);
  and (_10812_, _10811_, _10809_);
  or (_10814_, _10812_, _08650_);
  nand (_10815_, _08650_, _09584_);
  and (_10817_, _10815_, _10814_);
  or (_10818_, _10817_, _08646_);
  and (_10819_, _10818_, _10808_);
  or (_10820_, _10819_, _08666_);
  or (_10821_, _08671_, word_in[29]);
  and (_13875_, _10821_, _10820_);
  and (_10822_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_10823_, _08655_, word_in[6]);
  nor (_10824_, _10823_, _10822_);
  nor (_10825_, _10824_, _08650_);
  and (_10826_, _08650_, word_in[14]);
  or (_10827_, _10826_, _10825_);
  and (_10828_, _10827_, _08647_);
  and (_10829_, _09383_, _08646_);
  or (_10830_, _10829_, _08666_);
  or (_10831_, _10830_, _10828_);
  or (_10832_, _08671_, word_in[30]);
  and (_13876_, _10832_, _10831_);
  and (_10833_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_10834_, _05550_, _05677_);
  or (_10835_, _10834_, _10833_);
  and (_10033_, _10835_, _05552_);
  and (_10836_, _08009_, _10632_);
  nand (_10837_, _10836_, _06763_);
  or (_10838_, _10836_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_10839_, _10838_, _06532_);
  and (_10841_, _10839_, _10837_);
  or (_10842_, _10841_, _06561_);
  and (_10119_, _10842_, _05552_);
  and (_10843_, _05715_, _05819_);
  and (_10844_, _10843_, _05737_);
  and (_10845_, _10844_, _05837_);
  and (_10846_, _05875_, _05827_);
  and (_10847_, _10843_, _05809_);
  or (_10848_, _10847_, _10846_);
  or (_10849_, _10848_, _10845_);
  and (_10850_, _05851_, _05738_);
  and (_10851_, _10843_, _05814_);
  or (_10852_, _10851_, _10850_);
  or (_10853_, _10852_, _10849_);
  or (_10854_, _10853_, _05889_);
  and (_10855_, _10854_, _05547_);
  and (_10856_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_10857_, _10856_, _10855_);
  or (_10858_, _10857_, _05902_);
  and (_10247_, _10858_, _05552_);
  not (_10859_, _06775_);
  nor (_10860_, _10859_, _06020_);
  and (_10861_, _10860_, _07443_);
  nand (_10862_, _10861_, _06030_);
  and (_10863_, _10862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_10864_, _10863_, _08991_);
  nand (_10865_, _06030_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_10866_, _10865_, _08364_);
  or (_10867_, _10866_, _08367_);
  and (_10868_, _10867_, _10861_);
  or (_10869_, _10868_, _10864_);
  nand (_10870_, _08991_, _08386_);
  and (_10871_, _10870_, _05552_);
  and (_10254_, _10871_, _10869_);
  and (_10872_, _10861_, _06771_);
  nand (_10873_, _10872_, _06763_);
  nor (_10874_, _06326_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  nand (_10875_, _09010_, _09006_);
  or (_10876_, _10875_, _09002_);
  and (_10877_, _10876_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_10878_, _10877_, _10874_);
  or (_10879_, _10878_, _10872_);
  and (_10880_, _10879_, _10873_);
  or (_10881_, _10880_, _08991_);
  nand (_10882_, _08991_, _06811_);
  and (_10883_, _10882_, _05552_);
  and (_10257_, _10883_, _10881_);
  nor (_10884_, _09153_, _09086_);
  nor (_10885_, _10884_, _09154_);
  or (_10886_, _10885_, _09039_);
  or (_10887_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_10888_, _10887_, _05605_);
  and (_10890_, _10888_, _10886_);
  and (_10891_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_10892_, _10891_, _10890_);
  and (_10263_, _10892_, _05552_);
  and (_10893_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_10894_, _05550_, _05611_);
  or (_10895_, _10894_, _10893_);
  and (_10269_, _10895_, _05552_);
  and (_10896_, _05894_, _05830_);
  and (_10897_, _06567_, _05808_);
  and (_10898_, _05715_, _05646_);
  and (_10899_, _10898_, _05840_);
  or (_10901_, _10899_, _10897_);
  or (_10902_, _10901_, _10896_);
  not (_10904_, _05716_);
  and (_10905_, _05808_, _05760_);
  nor (_10906_, _10905_, _05877_);
  nor (_10907_, _10906_, _10904_);
  nor (_10908_, _10906_, _05714_);
  and (_10909_, _05852_, _05738_);
  and (_10910_, _10909_, _06567_);
  or (_10911_, _10910_, _10908_);
  or (_10912_, _10911_, _10907_);
  and (_10913_, _05850_, _05840_);
  or (_10914_, _05896_, _05878_);
  or (_10915_, _10914_, _10913_);
  and (_10917_, _05853_, _05737_);
  and (_10918_, _06567_, _10917_);
  or (_10919_, _10918_, _05838_);
  or (_10920_, _10919_, _10915_);
  or (_10921_, _10920_, _10912_);
  or (_10922_, _10921_, _10902_);
  nand (_10923_, _05894_, _05828_);
  not (_10924_, _10923_);
  and (_10925_, _05827_, _05815_);
  nor (_10926_, _10925_, _10924_);
  not (_10927_, _10926_);
  and (_10929_, _05894_, _06569_);
  or (_10930_, _10929_, _10927_);
  and (_10931_, _05894_, _05810_);
  or (_10932_, _05846_, _05824_);
  and (_10933_, _10932_, _05894_);
  or (_10934_, _10933_, _10931_);
  or (_10935_, _10934_, _05897_);
  or (_10936_, _10935_, _10930_);
  and (_10937_, _10843_, _05877_);
  and (_10938_, _05737_, _05820_);
  and (_10939_, _10938_, _05839_);
  and (_10940_, _10905_, _10843_);
  or (_10941_, _10940_, _10939_);
  or (_10942_, _10941_, _10937_);
  and (_10943_, _10843_, _05840_);
  or (_10944_, _10943_, _06569_);
  or (_10945_, _10938_, _10844_);
  and (_10946_, _10945_, _10944_);
  and (_10947_, _06568_, _05737_);
  or (_10948_, _10947_, _10946_);
  or (_10949_, _10948_, _10942_);
  or (_10950_, _10949_, _10936_);
  or (_10952_, _10950_, _10922_);
  and (_10953_, _10952_, _05547_);
  and (_10955_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_10956_, _06575_, _05893_);
  and (_10957_, _05896_, _05545_);
  and (_10958_, _05897_, _05545_);
  nor (_10959_, _10958_, _10957_);
  nor (_10960_, _10959_, _05546_);
  or (_10961_, _10960_, _10956_);
  or (_10962_, _10961_, _10955_);
  or (_10963_, _10962_, _10953_);
  and (_10282_, _10963_, _05552_);
  nor (_10964_, _09154_, _09078_);
  nor (_10965_, _10964_, _09155_);
  or (_10966_, _10965_, _09039_);
  or (_10967_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_10968_, _10967_, _05605_);
  and (_10969_, _10968_, _10966_);
  and (_10970_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_10971_, _10970_, _10969_);
  and (_10298_, _10971_, _05552_);
  nor (_10972_, _09152_, _09089_);
  nor (_10973_, _10972_, _09153_);
  or (_10974_, _10973_, _09039_);
  or (_10975_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_10976_, _10975_, _05605_);
  and (_10977_, _10976_, _10974_);
  and (_10978_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_10979_, _10978_, _10977_);
  and (_10302_, _10979_, _05552_);
  nor (_10980_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_10981_, _10980_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not (_10982_, _10981_);
  or (_10983_, _10982_, _08144_);
  or (_10984_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_10986_, _10984_, _05552_);
  and (_10604_, _10986_, _10983_);
  and (_10987_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_10988_, _05550_, _05921_);
  or (_10989_, _10988_, _10987_);
  and (_10623_, _10989_, _05552_);
  and (_10990_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not (_10991_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor (_10992_, _05550_, _10991_);
  or (_10993_, _10992_, _10990_);
  and (_10625_, _10993_, _05552_);
  and (_10994_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  not (_10995_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_10996_, _05550_, _10995_);
  or (_10997_, _10996_, _10994_);
  and (_10628_, _10997_, _05552_);
  and (_10998_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_10999_, _05550_, _05553_);
  or (_11000_, _10999_, _10998_);
  and (_10631_, _11000_, _05552_);
  and (_11001_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not (_11002_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_11003_, _05550_, _11002_);
  or (_11004_, _11003_, _11001_);
  and (_10634_, _11004_, _05552_);
  and (_11005_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not (_11006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_11007_, _05550_, _11006_);
  or (_11008_, _11007_, _11005_);
  and (_10637_, _11008_, _05552_);
  and (_11009_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_11010_, _05550_, _05748_);
  or (_11011_, _11010_, _11009_);
  and (_10640_, _11011_, _05552_);
  or (_11012_, _10918_, _10908_);
  and (_11014_, _05878_, _05818_);
  and (_11015_, _10898_, _10905_);
  and (_11016_, _11015_, _05738_);
  or (_11017_, _11016_, _11014_);
  or (_11018_, _11017_, _11012_);
  or (_11019_, _11018_, _05889_);
  and (_11020_, _11015_, _05737_);
  and (_11022_, _10898_, _05877_);
  or (_11023_, _11022_, _05896_);
  or (_11024_, _11023_, _06568_);
  or (_11025_, _11024_, _11020_);
  or (_11026_, _11025_, _10902_);
  or (_11027_, _11026_, _11019_);
  and (_11028_, _05894_, _05860_);
  and (_11029_, _05894_, _05853_);
  or (_11030_, _11029_, _11028_);
  and (_11031_, _08761_, _05716_);
  or (_11032_, _11031_, _11030_);
  and (_11033_, _10938_, _05837_);
  or (_11035_, _11033_, _10943_);
  or (_11036_, _11035_, _10845_);
  or (_11037_, _11036_, _11032_);
  or (_11038_, _11037_, _10942_);
  or (_11039_, _11038_, _10936_);
  or (_11040_, _11039_, _11027_);
  and (_11041_, _11040_, _05547_);
  and (_11042_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_11043_, _11042_, _10961_);
  or (_11045_, _11043_, _11041_);
  and (_10693_, _11045_, _05552_);
  or (_11046_, _10982_, _07483_);
  or (_11048_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_11050_, _11048_, _05552_);
  and (_10731_, _11050_, _11046_);
  and (_11051_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not (_11052_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor (_11053_, _05550_, _11052_);
  or (_11054_, _11053_, _11051_);
  and (_10807_, _11054_, _05552_);
  and (_11056_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  not (_11057_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_11058_, _05550_, _11057_);
  or (_11059_, _11058_, _11056_);
  and (_10810_, _11059_, _05552_);
  and (_11060_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_11061_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_11062_, _05550_, _11061_);
  or (_11063_, _11062_, _11060_);
  and (_10813_, _11063_, _05552_);
  nand (_11064_, _07388_, _06949_);
  or (_11065_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_11066_, _11065_, _05552_);
  and (_10816_, _11066_, _11064_);
  nor (_11067_, _07211_, _06341_);
  and (_11068_, _06346_, _07211_);
  or (_11069_, _11068_, _11067_);
  and (_10840_, _11069_, _05552_);
  and (_11070_, _05852_, _05850_);
  and (_11071_, _11070_, _05886_);
  not (_11072_, _11071_);
  and (_11073_, _05850_, _05738_);
  and (_11074_, _11073_, _10905_);
  and (_11075_, _05850_, _05737_);
  and (_11076_, _11075_, _05808_);
  nor (_11077_, _11076_, _11074_);
  not (_11078_, _11077_);
  and (_11079_, _11071_, _05761_);
  nor (_11080_, _11079_, _11078_);
  nor (_11081_, _11080_, _05892_);
  and (_11082_, _11081_, _11072_);
  and (_11083_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11084_, _05546_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11085_, _11084_);
  and (_11086_, _06567_, _05840_);
  not (_11087_, _11086_);
  and (_11088_, _05895_, _06567_);
  nor (_11089_, _11088_, _10918_);
  and (_11090_, _11089_, _11087_);
  and (_11091_, _11090_, _05898_);
  nor (_11092_, _11091_, _11085_);
  nor (_11093_, _11071_, _10960_);
  not (_11094_, _11093_);
  nor (_11095_, _11094_, _11092_);
  nor (_11097_, _11095_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11098_, _11097_, _11083_);
  and (_11099_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11100_, _10905_, _05823_);
  nand (_11101_, _11100_, _05885_);
  or (_11102_, _11101_, _05884_);
  or (_11103_, _10940_, _10937_);
  and (_11105_, _05850_, _05846_);
  or (_11106_, _11105_, _05876_);
  nor (_11107_, _11106_, _11103_);
  not (_11108_, _10847_);
  nand (_11109_, _10843_, _05828_);
  and (_11111_, _11109_, _11108_);
  nor (_11112_, _10943_, _10851_);
  and (_11113_, _11112_, _11111_);
  or (_11114_, _10909_, _06570_);
  and (_11115_, _11114_, _10843_);
  nor (_11116_, _11115_, _11100_);
  and (_11117_, _11116_, _11113_);
  and (_11118_, _11117_, _11107_);
  and (_11119_, _11090_, _11118_);
  nor (_11120_, _11119_, _11085_);
  and (_11121_, _10905_, _05738_);
  nand (_11122_, _11121_, _05850_);
  and (_11123_, _10905_, _05737_);
  and (_11124_, _11123_, _05850_);
  nor (_11125_, _11124_, _05887_);
  and (_11126_, _11125_, _11122_);
  and (_11127_, _05859_, _05850_);
  and (_11128_, _11127_, _05886_);
  not (_11129_, _11128_);
  and (_11130_, _11129_, _11126_);
  nor (_11131_, _11130_, _05892_);
  not (_11132_, _05886_);
  and (_11133_, _05853_, _05850_);
  nor (_11134_, _11133_, _11127_);
  nor (_11135_, _11134_, _11132_);
  not (_11136_, _11135_);
  nor (_11137_, _11136_, _11131_);
  nor (_11138_, _11137_, _11120_);
  and (_11139_, _11138_, _11102_);
  nor (_11140_, _11139_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11141_, _11140_, _11099_);
  not (_11142_, _11141_);
  and (_11144_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11145_, _05816_);
  nor (_11147_, _05861_, _05842_);
  and (_11148_, _11147_, _11145_);
  and (_11149_, _10898_, _05860_);
  and (_11150_, _11149_, _05669_);
  and (_11151_, _11075_, _05827_);
  or (_11152_, _11151_, _11150_);
  and (_11153_, _10917_, _05823_);
  and (_11154_, _11073_, _05827_);
  or (_11155_, _11154_, _11153_);
  or (_11157_, _11155_, _05833_);
  nor (_11158_, _11157_, _11152_);
  and (_11159_, _11158_, _11148_);
  and (_11160_, _05857_, _05823_);
  nor (_11161_, _11160_, _05878_);
  and (_11163_, _11161_, _11077_);
  and (_11164_, _05854_, _05716_);
  nor (_11166_, _11164_, _05845_);
  and (_11167_, _05846_, _05822_);
  and (_11169_, _11167_, _05818_);
  nor (_11170_, _11169_, _05841_);
  and (_11171_, _11170_, _11166_);
  and (_11172_, _11171_, _11163_);
  nor (_11173_, _11100_, _10907_);
  and (_11174_, _05895_, _05823_);
  and (_11175_, _05826_, _05815_);
  nor (_11176_, _11175_, _11174_);
  and (_11177_, _11176_, _11173_);
  and (_11178_, _06570_, _05716_);
  not (_11179_, _11178_);
  and (_11180_, _05895_, _05820_);
  nor (_11181_, _11180_, _10846_);
  and (_11182_, _11181_, _11179_);
  nor (_11183_, _05858_, _05811_);
  and (_11185_, _11183_, _05856_);
  and (_11186_, _11185_, _11182_);
  and (_11187_, _11186_, _11177_);
  and (_11188_, _11187_, _11172_);
  and (_11189_, _11188_, _11159_);
  nor (_11190_, _11189_, _11085_);
  nor (_11192_, _11190_, _11135_);
  and (_11193_, _11192_, _11102_);
  nor (_11194_, _11193_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11195_, _11194_, _11144_);
  and (_11196_, _11195_, _11142_);
  and (_11197_, _11196_, _11098_);
  and (_11198_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_11199_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_11200_, _11199_, _11198_);
  and (_11201_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_11202_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_11203_, _11202_, _11201_);
  and (_11204_, _11203_, _11200_);
  and (_11205_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_11206_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_11207_, _11206_, _11205_);
  and (_11208_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_11209_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_11210_, _11209_, _11208_);
  and (_11211_, _11210_, _11207_);
  and (_11212_, _11211_, _11204_);
  nor (_11213_, _11212_, _07437_);
  not (_11214_, _06560_);
  and (_11216_, _07437_, _11214_);
  nor (_11217_, _11216_, _11213_);
  not (_11218_, _11217_);
  and (_11219_, _11218_, _11197_);
  not (_11220_, _11219_);
  nor (_11221_, _11195_, _11141_);
  and (_11222_, _11098_, _11221_);
  and (_11223_, _07443_, _06057_);
  and (_11224_, _11223_, _06524_);
  not (_11225_, _11224_);
  nor (_11226_, _11225_, _06560_);
  and (_11227_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_11228_, _11226_, _11227_);
  and (_11230_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_11231_, _11225_, _08041_);
  nor (_11232_, _11231_, _11230_);
  and (_11233_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  not (_11234_, _07975_);
  and (_11235_, _11224_, _11234_);
  nor (_11236_, _11235_, _11233_);
  nor (_11237_, _11224_, _06025_);
  not (_11238_, _07945_);
  and (_11239_, _11224_, _11238_);
  nor (_11240_, _11239_, _11237_);
  and (_11241_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_11242_, _11241_, _11236_);
  and (_11243_, _11242_, _11232_);
  and (_11244_, _11243_, _11228_);
  nor (_11245_, _11243_, _11228_);
  nor (_11246_, _11245_, _11244_);
  nor (_11247_, _11246_, _05936_);
  nor (_11248_, _11247_, _06012_);
  nor (_11249_, _11248_, _11224_);
  nor (_11250_, _11249_, _11226_);
  not (_11251_, _11250_);
  and (_11252_, _11251_, _11222_);
  not (_11253_, _11252_);
  not (_11254_, _06562_);
  and (_11255_, _11098_, _11141_);
  and (_11256_, _11255_, _11195_);
  and (_11257_, _11256_, _11254_);
  not (_11258_, _11195_);
  and (_11260_, _11255_, _11258_);
  nor (_11261_, _05547_, _06165_);
  nor (_11262_, _05616_, _05699_);
  and (_11263_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_11264_, _11263_, _11262_);
  and (_11265_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_11266_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_11267_, _11266_, _11265_);
  nor (_11268_, _05613_, _11002_);
  nor (_11269_, _05624_, _05695_);
  nor (_11270_, _11269_, _11268_);
  and (_11271_, _11270_, _11267_);
  and (_11272_, _11271_, _11264_);
  nor (_11273_, _11272_, _09039_);
  nor (_11274_, _11273_, _11261_);
  not (_11275_, _11274_);
  and (_11276_, _11275_, _11260_);
  nor (_11277_, _11276_, _11257_);
  and (_11278_, _11277_, _11253_);
  and (_11279_, _11278_, _11220_);
  nor (_11280_, _11279_, _06064_);
  and (_11281_, _11279_, _06064_);
  nor (_11282_, _11281_, _11280_);
  and (_11283_, _11224_, _06811_);
  and (_11284_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_11285_, _11225_, _07388_);
  nor (_11286_, _11285_, _11284_);
  and (_11287_, _11286_, _11244_);
  and (_11288_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_11289_, _11225_, _06306_);
  nor (_11290_, _11289_, _11288_);
  and (_11291_, _11290_, _11287_);
  and (_11292_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_11294_, _11225_, _08386_);
  nor (_11296_, _11294_, _11292_);
  and (_11297_, _11296_, _11291_);
  nor (_11299_, _11224_, _05959_);
  nor (_11300_, _11299_, _11297_);
  and (_11301_, _11299_, _11297_);
  or (_11303_, _11301_, _11300_);
  nor (_11304_, _11303_, _05936_);
  nor (_11305_, _11224_, _05963_);
  not (_11306_, _11305_);
  nor (_11307_, _11306_, _11304_);
  nor (_11308_, _11307_, _11283_);
  and (_11309_, _11308_, _11221_);
  not (_11310_, _11309_);
  nor (_11311_, _11195_, _11142_);
  nor (_11312_, _05547_, _06359_);
  nor (_11313_, _05616_, _05762_);
  nor (_11315_, _05631_, _05768_);
  nor (_11316_, _11315_, _11313_);
  and (_11317_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_11318_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_11320_, _11318_, _11317_);
  nor (_11321_, _05613_, _07743_);
  nor (_11322_, _05624_, _05770_);
  nor (_11323_, _11322_, _11321_);
  and (_11324_, _11323_, _11320_);
  and (_11325_, _11324_, _11316_);
  nor (_11326_, _11325_, _09039_);
  nor (_11327_, _11326_, _11312_);
  not (_11328_, _11327_);
  and (_11329_, _11328_, _11311_);
  not (_11330_, _11098_);
  not (_11331_, _07441_);
  and (_11332_, _11196_, _11331_);
  or (_11333_, _11332_, _11330_);
  nor (_11334_, _11333_, _11329_);
  and (_11335_, _11334_, _11310_);
  nor (_11336_, _11335_, _06911_);
  and (_11337_, _11335_, _06911_);
  nor (_11338_, _11337_, _11336_);
  nor (_11339_, _11296_, _11291_);
  nor (_11340_, _11339_, _11297_);
  nor (_11341_, _11340_, _05936_);
  nor (_11342_, _11341_, _05940_);
  nor (_11343_, _11342_, _11224_);
  nor (_11344_, _11343_, _11294_);
  not (_11345_, _11344_);
  and (_11346_, _11345_, _11222_);
  not (_11347_, _11346_);
  and (_11348_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_11349_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_11351_, _11349_, _11348_);
  and (_11352_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_11353_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_11354_, _11353_, _11352_);
  and (_11356_, _11354_, _11351_);
  and (_11358_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_11359_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_11360_, _11359_, _11358_);
  and (_11361_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_11362_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_11363_, _11362_, _11361_);
  and (_11364_, _11363_, _11360_);
  and (_11365_, _11364_, _11356_);
  nor (_11366_, _11365_, _07437_);
  not (_11367_, _08386_);
  and (_11368_, _11367_, _07437_);
  nor (_11370_, _11368_, _11366_);
  not (_11371_, _11370_);
  and (_11372_, _11371_, _11197_);
  not (_11373_, _11372_);
  nor (_11374_, _11196_, _11098_);
  nor (_11376_, _05547_, _06394_);
  nor (_11377_, _05616_, _05786_);
  nor (_11378_, _05631_, _05791_);
  nor (_11379_, _11378_, _11377_);
  and (_11380_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_11381_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_11382_, _11381_, _11380_);
  not (_11383_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_11384_, _05613_, _11383_);
  and (_11385_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_11386_, _11385_, _11384_);
  and (_11387_, _11386_, _11382_);
  and (_11388_, _11387_, _11379_);
  nor (_11389_, _11388_, _09039_);
  nor (_11390_, _11389_, _11376_);
  not (_11391_, _11390_);
  and (_11392_, _11391_, _11260_);
  nor (_11393_, _11392_, _11374_);
  and (_11394_, _11393_, _11373_);
  and (_11395_, _11394_, _11347_);
  nor (_11396_, _11395_, _06925_);
  and (_11397_, _11395_, _06925_);
  nor (_11398_, _11397_, _11396_);
  and (_11399_, _11398_, _11338_);
  and (_11400_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_11401_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_11402_, _11401_, _11400_);
  and (_11403_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_11404_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_11405_, _11404_, _11403_);
  and (_11406_, _11405_, _11402_);
  and (_11407_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_11408_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor (_11409_, _11408_, _11407_);
  and (_11410_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_11411_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_11412_, _11411_, _11410_);
  and (_11413_, _11412_, _11409_);
  and (_11414_, _11413_, _11406_);
  nor (_11415_, _11414_, _07437_);
  and (_11416_, _07437_, _06307_);
  nor (_11418_, _11416_, _11415_);
  not (_11419_, _11418_);
  and (_11420_, _11419_, _11197_);
  not (_11421_, _11311_);
  and (_11422_, _11374_, _11421_);
  nor (_11423_, _11422_, _11420_);
  nor (_11424_, _11290_, _11287_);
  nor (_11425_, _11424_, _11291_);
  nor (_11426_, _11425_, _05936_);
  nor (_11427_, _11426_, _05993_);
  nor (_11428_, _11427_, _11224_);
  nor (_11429_, _11428_, _11289_);
  not (_11430_, _11429_);
  and (_11431_, _11430_, _11222_);
  nor (_11432_, _05547_, _06074_);
  nor (_11433_, _05616_, _05748_);
  nor (_11434_, _05631_, _05743_);
  nor (_11436_, _11434_, _11433_);
  and (_11437_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_11439_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_11440_, _11439_, _11437_);
  not (_11441_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_11442_, _05613_, _11441_);
  and (_11443_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_11444_, _11443_, _11442_);
  and (_11445_, _11444_, _11440_);
  and (_11446_, _11445_, _11436_);
  nor (_11447_, _11446_, _09039_);
  nor (_11448_, _11447_, _11432_);
  not (_11449_, _11448_);
  and (_11450_, _11449_, _11260_);
  nor (_11451_, _11450_, _11431_);
  and (_11452_, _11451_, _11423_);
  nor (_11453_, _11452_, _06764_);
  and (_11454_, _11452_, _06764_);
  nor (_11455_, _11454_, _11453_);
  nor (_11456_, _05547_, _06143_);
  and (_11457_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_11458_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_11459_, _11458_, _11457_);
  and (_11460_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_11461_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_11462_, _11461_, _11460_);
  nor (_11463_, _05613_, _11061_);
  and (_11464_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_11465_, _11464_, _11463_);
  and (_11466_, _11465_, _11462_);
  and (_11467_, _11466_, _11459_);
  nor (_11468_, _11467_, _09039_);
  nor (_11469_, _11468_, _11456_);
  not (_11470_, _11469_);
  and (_11471_, _11470_, _11260_);
  and (_11472_, _11256_, _07391_);
  nor (_11473_, _11472_, _11471_);
  and (_11474_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_11475_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_11476_, _11475_, _11474_);
  and (_11477_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_11478_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_11479_, _11478_, _11477_);
  and (_11480_, _11479_, _11476_);
  and (_11481_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_11482_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_11483_, _11482_, _11481_);
  and (_11484_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_11485_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_11486_, _11485_, _11484_);
  and (_11487_, _11486_, _11483_);
  and (_11488_, _11487_, _11480_);
  nor (_11489_, _11488_, _07437_);
  not (_11490_, _07388_);
  and (_11491_, _07437_, _11490_);
  nor (_11492_, _11491_, _11489_);
  not (_11493_, _11492_);
  and (_11494_, _11493_, _11197_);
  not (_11495_, _11494_);
  nor (_11496_, _11286_, _11244_);
  nor (_11497_, _11496_, _11287_);
  nor (_11499_, _11497_, _05936_);
  nor (_11500_, _11499_, _05976_);
  nor (_11501_, _11500_, _11224_);
  nor (_11502_, _11501_, _11285_);
  not (_11503_, _11502_);
  and (_11505_, _11503_, _11222_);
  and (_11506_, _11330_, _11141_);
  nor (_11507_, _11506_, _11505_);
  and (_11508_, _11507_, _11495_);
  and (_11509_, _11508_, _11473_);
  nor (_11510_, _11509_, _06527_);
  and (_11511_, _11509_, _06527_);
  nor (_11512_, _11511_, _11510_);
  and (_11513_, _11512_, _11455_);
  and (_11514_, _11513_, _11399_);
  and (_11515_, _11514_, _11282_);
  nor (_11516_, _06771_, _06967_);
  and (_11518_, _11516_, _11515_);
  and (_11519_, _11518_, _11082_);
  not (_11520_, _11519_);
  not (_11521_, _07224_);
  not (_11522_, _11131_);
  nor (_11523_, _06668_, _06628_);
  and (_11524_, _06668_, _06628_);
  nor (_11525_, _11524_, _11523_);
  nor (_11526_, _07680_, _06654_);
  nand (_11527_, _11526_, _08117_);
  nor (_11528_, _11527_, _11071_);
  and (_11529_, _11528_, _07462_);
  not (_11530_, _11529_);
  nor (_11531_, _11530_, _11525_);
  and (_11532_, _11531_, _07614_);
  and (_11533_, _11532_, _11522_);
  and (_11534_, _11533_, _07528_);
  and (_11535_, _11534_, _11521_);
  and (_11536_, _11082_, _06140_);
  and (_11537_, _11079_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_11538_, _11081_, _11072_);
  nor (_11539_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_11540_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_11541_, _11540_, _11539_);
  nor (_11542_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_11543_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_11544_, _11543_, _11542_);
  and (_11545_, _11544_, _11541_);
  and (_11546_, _11545_, _11538_);
  or (_11547_, _11546_, _11537_);
  or (_11548_, _11547_, _11536_);
  nor (_11549_, _11548_, _11535_);
  and (_11550_, _10938_, _05814_);
  not (_11552_, _11550_);
  nand (_11553_, _05846_, _05716_);
  nand (_11555_, _05828_, _05716_);
  and (_11556_, _11555_, _10923_);
  and (_11557_, _11556_, _11553_);
  and (_11558_, _11557_, _11552_);
  and (_11559_, _10938_, _05827_);
  not (_11560_, _11559_);
  and (_11561_, _11560_, _11109_);
  or (_11562_, _05877_, _10917_);
  nand (_11563_, _11562_, _05850_);
  and (_11564_, _11563_, _11561_);
  nand (_11565_, _11564_, _11558_);
  nor (_11566_, _11565_, _11124_);
  not (_11567_, _11566_);
  and (_11568_, _11567_, _11549_);
  not (_11569_, _11568_);
  and (_11570_, _05857_, _05850_);
  nor (_11571_, _11570_, _10918_);
  not (_11572_, _11122_);
  or (_11573_, _11572_, _05887_);
  nor (_11574_, _11134_, _05737_);
  nor (_11575_, _11574_, _11573_);
  or (_11576_, _11575_, _11549_);
  and (_11577_, _11576_, _11571_);
  and (_11578_, _11577_, _11569_);
  nor (_11579_, _11578_, _11132_);
  not (_11580_, _11101_);
  and (_11581_, _05823_, _05809_);
  nor (_11582_, _05869_, _11581_);
  nor (_11583_, _11085_, _11582_);
  nor (_11584_, _11583_, _11580_);
  not (_11585_, _11584_);
  nor (_11586_, _11585_, _11579_);
  not (_11587_, _08935_);
  and (_11589_, _11538_, _11587_);
  nor (_11590_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_11591_, _11590_);
  nor (_11592_, _11591_, _08009_);
  and (_11593_, _11592_, _06532_);
  not (_11594_, _11593_);
  and (_11595_, _11594_, _11079_);
  nor (_11596_, _11595_, _11589_);
  not (_11597_, _11596_);
  nor (_11598_, _11597_, _11586_);
  and (_11599_, _11196_, _11330_);
  not (_11600_, _11599_);
  and (_11601_, _11256_, _05819_);
  nor (_11602_, _05547_, _06228_);
  nor (_11603_, _05616_, _05611_);
  nor (_11604_, _05631_, _05615_);
  nor (_11605_, _11604_, _11603_);
  and (_11606_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_11607_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_11608_, _11607_, _11606_);
  not (_11609_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_11610_, _05613_, _11609_);
  and (_11611_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_11612_, _11611_, _11610_);
  and (_11613_, _11612_, _11608_);
  and (_11614_, _11613_, _11605_);
  nor (_11615_, _11614_, _09039_);
  nor (_11616_, _11615_, _11602_);
  not (_11617_, _11616_);
  and (_11618_, _11617_, _11260_);
  nor (_11619_, _11618_, _11601_);
  and (_11620_, _11619_, _11600_);
  nor (_11621_, _11241_, _11236_);
  nor (_11622_, _11621_, _11242_);
  nor (_11623_, _11622_, _05936_);
  nor (_11624_, _11623_, _06034_);
  nor (_11625_, _11624_, _11224_);
  nor (_11626_, _11625_, _11235_);
  not (_11627_, _11626_);
  and (_11628_, _11627_, _11222_);
  and (_11629_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_11630_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_11631_, _11630_, _11629_);
  and (_11632_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_11633_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_11634_, _11633_, _11632_);
  and (_11635_, _11634_, _11631_);
  and (_11636_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_11637_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_11638_, _11637_, _11636_);
  and (_11639_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_11640_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_11641_, _11640_, _11639_);
  and (_11642_, _11641_, _11638_);
  and (_11643_, _11642_, _11635_);
  nor (_11644_, _11643_, _07437_);
  and (_11645_, _11234_, _07437_);
  nor (_11646_, _11645_, _11644_);
  not (_11647_, _11646_);
  and (_11648_, _11647_, _11197_);
  nor (_11649_, _11648_, _11628_);
  and (_11650_, _11649_, _11620_);
  nor (_11651_, _11650_, _06043_);
  and (_11652_, _11650_, _06043_);
  nor (_11653_, _11652_, _11651_);
  and (_11654_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_11655_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_11656_, _11655_, _11654_);
  and (_11657_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_11658_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_11660_, _11658_, _11657_);
  and (_11661_, _11660_, _11656_);
  and (_11662_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_11663_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_11664_, _11663_, _11662_);
  and (_11665_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_11666_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_11667_, _11666_, _11665_);
  and (_11668_, _11667_, _11664_);
  and (_11669_, _11668_, _11661_);
  nor (_11670_, _11669_, _07437_);
  and (_11671_, _11238_, _07437_);
  nor (_11672_, _11671_, _11670_);
  not (_11673_, _11672_);
  and (_11674_, _11673_, _11197_);
  nor (_11675_, _05547_, _06186_);
  nor (_11676_, _05616_, _05656_);
  and (_11677_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_11678_, _11677_, _11676_);
  and (_11679_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_11680_, _05624_, _05652_);
  nor (_11682_, _11680_, _11679_);
  and (_11683_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_11684_, _05613_, _11006_);
  nor (_11686_, _11684_, _11683_);
  and (_11687_, _11686_, _11682_);
  and (_11688_, _11687_, _11678_);
  nor (_11689_, _11688_, _09039_);
  nor (_11690_, _11689_, _11675_);
  not (_11691_, _11690_);
  and (_11692_, _11691_, _11260_);
  nor (_11693_, _11692_, _11674_);
  nor (_11694_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_11695_, _11694_, _11241_);
  nor (_11696_, _11695_, _05936_);
  nor (_11697_, _11696_, _06026_);
  nor (_11698_, _11697_, _11224_);
  nor (_11699_, _11698_, _11239_);
  not (_11700_, _11699_);
  and (_11701_, _11700_, _11222_);
  and (_11702_, _11256_, _05669_);
  nor (_11703_, _11702_, _11701_);
  and (_11704_, _11703_, _11693_);
  and (_11705_, _11704_, _06031_);
  nor (_11706_, _11704_, _06031_);
  or (_11707_, _11706_, _11705_);
  nor (_11708_, _11707_, _11653_);
  and (_11709_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_11710_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_11711_, _11710_, _11709_);
  and (_11712_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_11713_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_11714_, _11713_, _11712_);
  and (_11715_, _11714_, _11711_);
  and (_11716_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_11717_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_11718_, _11717_, _11716_);
  and (_11719_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_11721_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_11722_, _11721_, _11719_);
  and (_11723_, _11722_, _11718_);
  and (_11724_, _11723_, _11715_);
  nor (_11725_, _11724_, _07437_);
  not (_11726_, _08041_);
  and (_11727_, _11726_, _07437_);
  nor (_11728_, _11727_, _11725_);
  not (_11729_, _11728_);
  and (_11730_, _11729_, _11197_);
  nor (_11731_, _05547_, _06209_);
  nor (_11732_, _05616_, _05677_);
  and (_11733_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11734_, _11733_, _11732_);
  and (_11735_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_11736_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_11737_, _11736_, _11735_);
  and (_11738_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not (_11739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_11740_, _05613_, _11739_);
  nor (_11742_, _11740_, _11738_);
  and (_11743_, _11742_, _11737_);
  and (_11744_, _11743_, _11734_);
  nor (_11745_, _11744_, _09039_);
  nor (_11746_, _11745_, _11731_);
  not (_11747_, _11746_);
  and (_11749_, _11747_, _11260_);
  nor (_11750_, _11749_, _11730_);
  nor (_11751_, _11242_, _11232_);
  nor (_11752_, _11751_, _11243_);
  nor (_11753_, _11752_, _05936_);
  nor (_11754_, _11753_, _06046_);
  nor (_11756_, _11754_, _11224_);
  nor (_11757_, _11756_, _11231_);
  not (_11759_, _11757_);
  and (_11760_, _11759_, _11222_);
  and (_11761_, _11256_, _05693_);
  nor (_11762_, _11761_, _11760_);
  and (_11763_, _11762_, _11750_);
  nor (_11764_, _11763_, _06054_);
  and (_11765_, _11763_, _06054_);
  nor (_11766_, _11765_, _11764_);
  nor (_11767_, _11766_, _06816_);
  and (_11768_, _11767_, _11708_);
  and (_11769_, _11768_, _11515_);
  nor (_11770_, _05971_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_11771_, _11770_, _11769_);
  not (_11772_, _11771_);
  and (_11773_, _11772_, _11598_);
  and (_11774_, _11773_, _11520_);
  and (_11775_, _11557_, _11126_);
  nand (_11776_, _11775_, _11561_);
  nand (_11777_, _11776_, _05886_);
  and (_11778_, _10905_, _11084_);
  and (_11779_, _11778_, _05850_);
  and (_11780_, _11084_, _11581_);
  nor (_11781_, _11780_, _11779_);
  and (_11782_, _11781_, _11102_);
  nand (_11783_, _11782_, _11777_);
  and (_11784_, _10918_, _05886_);
  nor (_11785_, _11784_, _11583_);
  nor (_11786_, _11785_, _11783_);
  not (_11787_, _11786_);
  nor (_11788_, _11550_, _11070_);
  nand (_11789_, _11788_, _11571_);
  nand (_11790_, _11789_, _05886_);
  nand (_11791_, _11790_, _11777_);
  nor (_11792_, _11791_, _11787_);
  and (_11793_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_11794_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_11795_, _11794_, _11793_);
  and (_11796_, \oc8051_top_1.oc8051_memory_interface1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_11797_, _11796_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_11799_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_11800_, _11799_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_11801_, _11800_, _11797_);
  and (_11802_, _11801_, _11795_);
  and (_11803_, _11802_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_11804_, _11803_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_11805_, _11804_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_11806_, _11805_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_11807_, _11806_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_11808_, _11806_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_11809_, _11808_, _11807_);
  and (_11810_, _11809_, _11792_);
  not (_11811_, _11102_);
  and (_11812_, _11811_, _07255_);
  and (_11813_, _11784_, _07360_);
  and (_11814_, _11780_, _11328_);
  and (_11815_, _11782_, _11777_);
  nand (_11816_, _11785_, _11815_);
  nor (_11817_, _11816_, _11791_);
  and (_11818_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_11819_, _11818_, _11814_);
  or (_11820_, _11819_, _11813_);
  or (_11821_, _11820_, _11812_);
  nor (_11822_, _11821_, _11810_);
  nand (_11824_, _11822_, _11774_);
  and (_11825_, _11783_, _07758_);
  and (_11827_, _11815_, _11327_);
  nor (_11828_, _11827_, _11825_);
  nor (_11829_, _11828_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_11830_, _11828_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_11831_, _05547_, _06482_);
  and (_11832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11833_, _05616_, _11383_);
  nor (_11834_, _05624_, _05791_);
  or (_11835_, _11834_, _11833_);
  nor (_11836_, _05613_, _05907_);
  nor (_11837_, _05631_, _05786_);
  or (_11838_, _11837_, _11836_);
  or (_11839_, _11838_, _11835_);
  and (_11840_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_11842_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_11843_, _11842_, _11840_);
  or (_11844_, _11843_, _11839_);
  and (_11845_, _11844_, _05671_);
  or (_11846_, _11845_, _11832_);
  and (_11847_, _11846_, _05547_);
  nor (_11848_, _11847_, _11831_);
  and (_11849_, _11848_, _11783_);
  and (_11850_, _11815_, _11390_);
  nor (_11851_, _11850_, _11849_);
  and (_11852_, _11851_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_11853_, _11851_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_11854_, _11853_, _11852_);
  nor (_11855_, _05547_, _06079_);
  and (_11856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11857_, _05613_, _11057_);
  nor (_11858_, _05624_, _05743_);
  nor (_11859_, _11858_, _11857_);
  and (_11860_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_11861_, _05631_, _05748_);
  nor (_11862_, _11861_, _11860_);
  and (_11863_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_11864_, _05616_, _11441_);
  nor (_11865_, _11864_, _11863_);
  and (_11866_, _11865_, _11862_);
  and (_11867_, _11866_, _11859_);
  nor (_11868_, _11867_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11870_, _11868_, _11856_);
  nor (_11871_, _11870_, _05548_);
  nor (_11872_, _11871_, _11855_);
  and (_11873_, _11872_, _11783_);
  and (_11874_, _11815_, _11448_);
  nor (_11875_, _11874_, _11873_);
  nor (_11876_, _11875_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_11877_, _11875_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_11878_, _05547_, _06145_);
  and (_11879_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11881_, _05616_, _11061_);
  and (_11883_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_11884_, _11883_, _11881_);
  nor (_11886_, _05613_, _10995_);
  and (_11887_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_11889_, _11887_, _11886_);
  or (_11890_, _11889_, _11884_);
  and (_11891_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_11892_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_11893_, _11892_, _11891_);
  or (_11895_, _11893_, _11890_);
  and (_11896_, _11895_, _05671_);
  or (_11898_, _11896_, _11879_);
  and (_11899_, _11898_, _05547_);
  nor (_11900_, _11899_, _11878_);
  and (_11901_, _11900_, _11783_);
  and (_11902_, _11815_, _11469_);
  nor (_11903_, _11902_, _11901_);
  nand (_11904_, _11903_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_11905_, _05547_, _06167_);
  and (_11906_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11907_, _05616_, _11002_);
  and (_11908_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_11909_, _11908_, _11907_);
  and (_11910_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_11911_, _05631_, _05699_);
  or (_11912_, _11911_, _11910_);
  or (_11913_, _11912_, _11909_);
  and (_11914_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_11915_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_11916_, _11915_, _11914_);
  or (_11917_, _11916_, _11913_);
  and (_11918_, _11917_, _05671_);
  or (_11919_, _11918_, _11906_);
  and (_11920_, _11919_, _05547_);
  nor (_11921_, _11920_, _11905_);
  and (_11922_, _11921_, _11783_);
  and (_11923_, _11815_, _11274_);
  nor (_11924_, _11923_, _11922_);
  nor (_11925_, _11924_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_11926_, _11924_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_11927_, _05547_, _06207_);
  and (_11928_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_11929_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_11930_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11931_, _11930_, _11929_);
  nor (_11932_, _05616_, _11739_);
  and (_11933_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_11934_, _11933_, _11932_);
  nor (_11935_, _05613_, _08689_);
  nor (_11936_, _05631_, _05677_);
  nor (_11937_, _11936_, _11935_);
  and (_11938_, _11937_, _11934_);
  and (_11939_, _11938_, _11931_);
  nor (_11940_, _11939_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11941_, _11940_, _11928_);
  nor (_11942_, _11941_, _05548_);
  nor (_11943_, _11942_, _11927_);
  not (_11944_, _11943_);
  or (_11945_, _11944_, _11815_);
  or (_11946_, _11783_, _11747_);
  nand (_11947_, _11946_, _11945_);
  or (_11948_, _11947_, _06217_);
  not (_11949_, _11948_);
  nor (_11950_, _05547_, _06230_);
  and (_11951_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11952_, _05613_, _05553_);
  nor (_11953_, _05624_, _05615_);
  nor (_11954_, _11953_, _11952_);
  and (_11955_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor (_11956_, _05631_, _05611_);
  nor (_11957_, _11956_, _11955_);
  and (_11958_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_11959_, _05616_, _11609_);
  nor (_11960_, _11959_, _11958_);
  and (_11961_, _11960_, _11957_);
  and (_11962_, _11961_, _11954_);
  nor (_11964_, _11962_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11965_, _11964_, _11951_);
  nor (_11966_, _11965_, _05548_);
  nor (_11967_, _11966_, _11950_);
  not (_11968_, _11967_);
  or (_11969_, _11968_, _11815_);
  or (_11970_, _11783_, _11617_);
  and (_11971_, _11970_, _11969_);
  nand (_11972_, _11971_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_11973_, _05547_, _06188_);
  and (_11975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11976_, _05616_, _11006_);
  and (_11977_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_11978_, _11977_, _11976_);
  and (_11979_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_11980_, _05631_, _05656_);
  or (_11982_, _11980_, _11979_);
  or (_11983_, _11982_, _11978_);
  and (_11985_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_11986_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_11987_, _11986_, _11985_);
  or (_11988_, _11987_, _11983_);
  and (_11989_, _11988_, _05671_);
  or (_11990_, _11989_, _11975_);
  and (_11991_, _11990_, _05547_);
  nor (_11993_, _11991_, _11973_);
  not (_11994_, _11993_);
  or (_11995_, _11994_, _11815_);
  or (_11996_, _11783_, _11691_);
  and (_11997_, _11996_, _11995_);
  and (_11998_, _11997_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_11999_, _11971_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_12000_, _11999_, _11972_);
  and (_12001_, _12000_, _11998_);
  not (_12002_, _12001_);
  nand (_12004_, _12002_, _11972_);
  nand (_12005_, _11947_, _06217_);
  and (_12006_, _12005_, _11948_);
  and (_12007_, _12006_, _12004_);
  or (_12008_, _12007_, _11949_);
  nor (_12009_, _12008_, _11926_);
  nor (_12010_, _12009_, _11925_);
  or (_12012_, _11903_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12013_, _12012_, _11904_);
  nand (_12014_, _12013_, _12010_);
  nand (_12015_, _12014_, _11904_);
  nor (_12016_, _12015_, _11877_);
  nor (_12017_, _12016_, _11876_);
  and (_12018_, _12017_, _11854_);
  or (_12019_, _12018_, _11852_);
  nor (_12020_, _12019_, _11830_);
  nor (_12021_, _12020_, _11829_);
  or (_12022_, _12021_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_12024_, _12022_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_12025_, _12024_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_12027_, _12025_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_12028_, _12027_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_12029_, _12028_, _06085_);
  nand (_12030_, _12029_, _06487_);
  nand (_12031_, _12030_, _11828_);
  not (_12032_, _11828_);
  and (_12034_, _12021_, _11797_);
  nand (_12035_, _12034_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_12036_, _12035_, _06148_);
  nor (_12037_, _12036_, _06085_);
  nand (_12038_, _12037_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_12039_, _12038_, _12032_);
  nand (_12040_, _12039_, _12031_);
  nand (_12041_, _12040_, _06590_);
  or (_12043_, _12040_, _06590_);
  and (_12044_, _12043_, _12041_);
  and (_12045_, _11084_, _05850_);
  and (_12046_, _12045_, _10905_);
  and (_12047_, _11561_, _11134_);
  and (_12048_, _12047_, _11126_);
  and (_12050_, _11571_, _11558_);
  and (_12051_, _12050_, _12048_);
  nor (_12052_, _12051_, _11132_);
  nor (_12053_, _12052_, _12046_);
  nor (_12054_, _12053_, _11786_);
  and (_12056_, _12054_, _12044_);
  or (_12057_, _12056_, _11824_);
  and (_12059_, _08238_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_12060_, _12059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12061_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12062_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_12063_, _12062_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12064_, _12063_, _12061_);
  and (_12066_, _12064_, _12060_);
  and (_12068_, _12066_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_12069_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_12071_, _12069_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_12072_, _12071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_12073_, _12072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_12074_, _12072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_12075_, _12074_, _12073_);
  or (_12076_, _12075_, _11774_);
  and (_12077_, _12076_, _05552_);
  and (_10889_, _12077_, _12057_);
  and (_12080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _05556_);
  and (_12081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_12082_, _12081_, _12080_);
  and (_10900_, _12082_, _05552_);
  or (_12083_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_12085_, _05550_, _05743_);
  and (_12086_, _12085_, _05552_);
  and (_10903_, _12086_, _12083_);
  and (_12088_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_12089_, _05550_, _11441_);
  or (_12090_, _12089_, _12088_);
  and (_10916_, _12090_, _05552_);
  and (_12091_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_12092_, _05550_, _05656_);
  or (_12093_, _12092_, _12091_);
  and (_10928_, _12093_, _05552_);
  and (_10951_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not (_12094_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_12095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not (_12096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_12097_, _10874_, _12096_);
  not (_12098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_12099_, _12098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_12100_, _12099_, _12097_);
  nor (_12101_, _12100_, _12095_);
  nand (_12103_, _12101_, _12094_);
  nor (_12104_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_12106_, _12104_, _12101_);
  nand (_12107_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_12108_, _12107_, _12106_);
  and (_12109_, _12108_, _05552_);
  and (_10954_, _12109_, _12103_);
  and (_12111_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_12112_, _05550_, _11383_);
  or (_12114_, _12112_, _12111_);
  and (_10985_, _12114_, _05552_);
  nor (_12116_, _09136_, _09133_);
  nor (_12117_, _12116_, _09137_);
  or (_12118_, _12117_, _09039_);
  or (_12119_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_12120_, _12119_, _05605_);
  and (_12121_, _12120_, _12118_);
  and (_12122_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_12123_, _12122_, _12121_);
  and (_11013_, _12123_, _05552_);
  and (_12124_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07768_);
  and (_12125_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_12126_, _12125_, _12124_);
  and (_11034_, _12126_, _05552_);
  nor (_11044_, _11921_, rst);
  nor (_11047_, _11746_, rst);
  nand (_12127_, _07483_, _06973_);
  and (_12128_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_12129_, _10632_, _08048_);
  nor (_12130_, _10632_, _06179_);
  nor (_12131_, _12130_, _12129_);
  nor (_12132_, _12131_, _08924_);
  nor (_12133_, _12132_, _12128_);
  and (_12134_, _12133_, _07261_);
  and (_12136_, _12134_, _12127_);
  and (_12137_, _07515_, _07260_);
  nor (_12138_, _12137_, _12136_);
  and (_11049_, _12138_, _05552_);
  and (_12139_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not (_12140_, _05550_);
  and (_12141_, _12140_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_12142_, _12141_, _12139_);
  and (_11055_, _12142_, _05552_);
  nor (_12143_, _09151_, _09091_);
  nor (_12144_, _12143_, _09152_);
  or (_12145_, _12144_, _09039_);
  or (_12146_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_12147_, _12146_, _07933_);
  and (_12148_, _12147_, _12145_);
  and (_12149_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_12150_, _12149_, _05552_);
  or (_11096_, _12150_, _12148_);
  and (_12152_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_12153_, _05550_, _05699_);
  or (_12154_, _12153_, _12152_);
  and (_11104_, _12154_, _05552_);
  nand (_12155_, _12027_, _11828_);
  nand (_12156_, _12035_, _12032_);
  and (_12157_, _12156_, _12155_);
  nand (_12159_, _12157_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_12160_, _11791_, _11779_);
  nor (_12161_, _12160_, _11786_);
  or (_12162_, _12157_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_12163_, _12162_, _12161_);
  and (_12164_, _12163_, _12159_);
  or (_12165_, _07178_, _07176_);
  and (_12166_, _12165_, _07603_);
  or (_12167_, _12166_, _07446_);
  or (_12168_, _07200_, _07130_);
  and (_12169_, _12168_, _12167_);
  and (_12170_, _12169_, _06314_);
  and (_12171_, _06908_, _07211_);
  and (_12172_, _11525_, _06581_);
  or (_12173_, _06698_, _06628_);
  nor (_12174_, _06699_, _06678_);
  and (_12175_, _12174_, _12173_);
  nor (_12176_, _07467_, _06118_);
  nor (_12177_, _12176_, _06164_);
  and (_12178_, _06718_, _06164_);
  and (_12179_, _06128_, _06111_);
  and (_12180_, _06184_, _06131_);
  or (_12181_, _12180_, _12179_);
  nor (_12182_, _12181_, _12178_);
  nand (_12183_, _12182_, _07386_);
  nor (_12184_, _12183_, _12177_);
  nand (_12185_, _12184_, _07375_);
  or (_12186_, _12185_, _12175_);
  or (_12187_, _12186_, _12172_);
  or (_12188_, _12187_, _12171_);
  or (_12189_, _12188_, _12170_);
  and (_12190_, _12189_, _11811_);
  or (_12192_, _07299_, _07296_);
  nor (_12193_, _07300_, _06678_);
  and (_12194_, _12193_, _12192_);
  and (_12195_, _07719_, _07211_);
  nor (_12196_, _07322_, _06142_);
  nor (_12197_, _07330_, _06253_);
  or (_12198_, _12197_, _12196_);
  nand (_12199_, _12198_, _06379_);
  or (_12200_, _12198_, _06379_);
  and (_12201_, _12200_, _06266_);
  and (_12202_, _12201_, _12199_);
  or (_12203_, _06162_, _06253_);
  or (_12204_, _06625_, _06142_);
  and (_12205_, _12204_, _06295_);
  and (_12206_, _12205_, _12203_);
  and (_12207_, _06368_, _06746_);
  and (_12208_, _06625_, _06118_);
  and (_12209_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_12210_, _12209_, _12208_);
  or (_12211_, _12210_, _12207_);
  or (_12212_, _12211_, _12206_);
  or (_12213_, _12212_, _12202_);
  or (_12214_, _12213_, _12195_);
  or (_12215_, _12214_, _12194_);
  and (_12216_, _12215_, _11784_);
  nor (_12217_, _11803_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_12218_, _12217_, _11804_);
  and (_12219_, _12218_, _11792_);
  and (_12220_, _11780_, _11470_);
  or (_12221_, _12220_, _12219_);
  and (_12222_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_12223_, _12222_, _12221_);
  nor (_12224_, _12223_, _12216_);
  nand (_12225_, _12224_, _11774_);
  or (_12226_, _12225_, _12190_);
  or (_12227_, _12226_, _12164_);
  nor (_12228_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_12229_, _12228_, _12069_);
  or (_12230_, _12229_, _11774_);
  and (_12231_, _12230_, _05552_);
  and (_11110_, _12231_, _12227_);
  nor (_11143_, _11690_, rst);
  or (_12232_, _09130_, _09127_);
  and (_12233_, _12232_, _09131_);
  or (_12234_, _12233_, _09039_);
  or (_12235_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_12236_, _12235_, _05605_);
  and (_12237_, _12236_, _12234_);
  and (_12238_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_12239_, _12238_, _12237_);
  and (_11146_, _12239_, _05552_);
  nor (_11156_, _11728_, rst);
  or (_12240_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  nand (_12241_, _05550_, _10991_);
  and (_12242_, _12241_, _05552_);
  and (_11162_, _12242_, _12240_);
  or (_12243_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_12244_, _05550_, _05762_);
  and (_12245_, _12244_, _05552_);
  and (_11165_, _12245_, _12243_);
  or (_12246_, _09126_, _09123_);
  nor (_12247_, _09039_, _09127_);
  and (_12248_, _12247_, _12246_);
  and (_12249_, _09039_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_12250_, _12249_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_12251_, _12250_, _12248_);
  or (_12252_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _05605_);
  and (_12253_, _12252_, _05552_);
  and (_11168_, _12253_, _12251_);
  and (_11184_, _05693_, _05552_);
  nor (_12254_, _06306_, _06953_);
  and (_12255_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_12256_, _12255_, _06955_);
  or (_12257_, _12256_, _12254_);
  or (_12258_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_12259_, _12258_, _05552_);
  and (_11191_, _12259_, _12257_);
  and (_12260_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_12261_, _05550_, _05762_);
  or (_12262_, _12261_, _12260_);
  and (_11215_, _12262_, _05552_);
  not (_12263_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_12264_, _09504_, _06068_);
  nor (_12265_, _12264_, _12263_);
  and (_12266_, _09504_, _07976_);
  or (_12267_, _12266_, _12265_);
  and (_11229_, _12267_, _05552_);
  nor (_11259_, _11335_, rst);
  nand (_12268_, _11161_, _11089_);
  or (_12269_, _11028_, _05861_);
  or (_12270_, _12269_, _11153_);
  and (_12271_, _06567_, _05809_);
  and (_12272_, _12271_, _05737_);
  or (_12273_, _12272_, _12270_);
  or (_12274_, _12273_, _12268_);
  or (_12276_, _05860_, _05814_);
  and (_12277_, _12276_, _10843_);
  or (_12278_, _11150_, _11016_);
  or (_12279_, _12278_, _12277_);
  and (_12280_, _10898_, _05830_);
  and (_12282_, _05894_, _05846_);
  nor (_12283_, _05737_, _05714_);
  and (_12284_, _12283_, _05813_);
  or (_12285_, _12284_, _12282_);
  or (_12287_, _12285_, _12280_);
  or (_12288_, _11103_, _10908_);
  or (_12289_, _12288_, _12287_);
  or (_12290_, _12289_, _12279_);
  and (_12291_, _11123_, _06567_);
  or (_12292_, _11025_, _12291_);
  or (_12293_, _12292_, _12290_);
  or (_12295_, _12293_, _12274_);
  and (_12296_, _12295_, _06576_);
  nor (_12297_, _11084_, rst);
  and (_12298_, _12297_, _05896_);
  and (_12299_, _05552_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_12300_, _12299_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_12301_, _12300_, _12298_);
  or (_11293_, _12301_, _12296_);
  and (_12302_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_12303_, _12302_, _10957_);
  and (_12304_, _12303_, _05552_);
  not (_12305_, _11112_);
  or (_12306_, _12305_, _10899_);
  not (_12307_, _11561_);
  and (_12308_, _12283_, _05814_);
  or (_12309_, _12308_, _10939_);
  or (_12310_, _12309_, _12307_);
  or (_12311_, _12310_, _12306_);
  nand (_12312_, _10905_, _06567_);
  and (_12313_, _10938_, _05859_);
  nor (_12314_, _12313_, _10937_);
  and (_12315_, _12314_, _11108_);
  nand (_12316_, _12315_, _12312_);
  or (_12317_, _12316_, _12311_);
  not (_12318_, _11022_);
  and (_12319_, _11161_, _12318_);
  not (_12320_, _12319_);
  or (_12321_, _12320_, _10930_);
  or (_12322_, _12321_, _12317_);
  and (_12324_, _10898_, _05824_);
  or (_12325_, _10931_, _05817_);
  or (_12327_, _12325_, _12324_);
  and (_12328_, _06567_, _05828_);
  or (_12329_, _12328_, _05829_);
  and (_12330_, _05810_, _05820_);
  and (_12331_, _10932_, _05820_);
  or (_12332_, _12331_, _12330_);
  or (_12333_, _12280_, _11154_);
  or (_12334_, _12333_, _12332_);
  or (_12335_, _12334_, _12329_);
  or (_12336_, _12335_, _12327_);
  or (_12337_, _12336_, _12322_);
  and (_12338_, _12337_, _06576_);
  or (_11295_, _12338_, _12304_);
  nor (_12339_, _07939_, _06560_);
  and (_12340_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or (_12341_, _12340_, _12339_);
  and (_11298_, _12341_, _05552_);
  nor (_12342_, _07939_, _06306_);
  and (_12344_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or (_12345_, _12344_, _12342_);
  and (_11302_, _12345_, _05552_);
  and (_12347_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07768_);
  and (_12348_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_12349_, _12348_, _12347_);
  and (_11314_, _12349_, _05552_);
  nor (_11319_, _11274_, rst);
  nor (_11350_, _11616_, rst);
  or (_12350_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand (_12351_, _05550_, _11006_);
  and (_12352_, _12351_, _05552_);
  and (_11355_, _12352_, _12350_);
  or (_12353_, _07731_, _05565_);
  or (_12354_, _07736_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_12355_, _12354_, _05552_);
  and (_11357_, _12355_, _12353_);
  nor (_12357_, _09143_, _09112_);
  nor (_12359_, _12357_, _09144_);
  or (_12360_, _12359_, _09039_);
  or (_12362_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12363_, _12362_, _07933_);
  and (_12364_, _12363_, _12360_);
  and (_12365_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12366_, _12365_, _05552_);
  or (_11369_, _12366_, _12364_);
  nor (_11375_, _07390_, rst);
  or (_12367_, _09149_, _09098_);
  nor (_12368_, _09039_, _09150_);
  and (_12369_, _12368_, _12367_);
  nor (_12371_, _09038_, _06235_);
  or (_12372_, _12371_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_12373_, _12372_, _12369_);
  or (_12374_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_12375_, _12374_, _05552_);
  and (_11417_, _12375_, _12373_);
  and (_12376_, _08362_, word_in[0]);
  or (_12377_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  or (_12378_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_12379_, _12378_, _12377_);
  and (_12380_, _12379_, _08279_);
  or (_12381_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  or (_12382_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_12384_, _12382_, _12381_);
  and (_12385_, _12384_, _08260_);
  or (_12387_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  or (_12388_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_12389_, _12388_, _12387_);
  and (_12390_, _12389_, _08257_);
  or (_12391_, _12390_, _12385_);
  or (_12392_, _12391_, _12380_);
  or (_12393_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  or (_12394_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_12395_, _12394_, _12393_);
  and (_12396_, _12395_, _08267_);
  or (_12397_, _12396_, _08286_);
  or (_12398_, _12397_, _12392_);
  or (_12399_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or (_12400_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_12401_, _12400_, _12399_);
  and (_12402_, _12401_, _08279_);
  or (_12403_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  or (_12404_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_12405_, _12404_, _12403_);
  and (_12406_, _12405_, _08260_);
  or (_12407_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or (_12408_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_12409_, _12408_, _12407_);
  and (_12410_, _12409_, _08257_);
  or (_12411_, _12410_, _12406_);
  or (_12412_, _12411_, _12402_);
  or (_12413_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  or (_12414_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_12415_, _12414_, _12413_);
  and (_12416_, _12415_, _08267_);
  or (_12417_, _12416_, _08243_);
  or (_12418_, _12417_, _12412_);
  and (_12419_, _12418_, _12398_);
  and (_12420_, _12419_, _08311_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _12420_, _12376_);
  and (_12421_, _08362_, word_in[1]);
  or (_12422_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  or (_12423_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_12424_, _12423_, _12422_);
  and (_12425_, _12424_, _08279_);
  or (_12426_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  or (_12427_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_12428_, _12427_, _12426_);
  and (_12429_, _12428_, _08260_);
  or (_12430_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  or (_12431_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_12432_, _12431_, _12430_);
  and (_12433_, _12432_, _08257_);
  or (_12434_, _12433_, _12429_);
  or (_12435_, _12434_, _12425_);
  or (_12436_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  or (_12437_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_12438_, _12437_, _12436_);
  and (_12439_, _12438_, _08267_);
  or (_12441_, _12439_, _08286_);
  or (_12442_, _12441_, _12435_);
  or (_12443_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  or (_12444_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_12445_, _12444_, _12443_);
  and (_12446_, _12445_, _08279_);
  or (_12447_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  or (_12448_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_12449_, _12448_, _12447_);
  and (_12450_, _12449_, _08260_);
  or (_12451_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  or (_12452_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_12453_, _12452_, _12451_);
  and (_12454_, _12453_, _08257_);
  or (_12456_, _12454_, _12450_);
  or (_12457_, _12456_, _12446_);
  or (_12458_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  or (_12459_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_12460_, _12459_, _12458_);
  and (_12461_, _12460_, _08267_);
  or (_12462_, _12461_, _08243_);
  or (_12463_, _12462_, _12457_);
  and (_12464_, _12463_, _12442_);
  and (_12465_, _12464_, _08311_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _12465_, _12421_);
  and (_12466_, _08362_, word_in[2]);
  or (_12468_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  or (_12469_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_12470_, _12469_, _12468_);
  and (_12471_, _12470_, _08279_);
  or (_12472_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  or (_12473_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_12474_, _12473_, _12472_);
  and (_12475_, _12474_, _08260_);
  or (_12476_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  or (_12477_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_12478_, _12477_, _12476_);
  and (_12479_, _12478_, _08257_);
  or (_12480_, _12479_, _12475_);
  or (_12481_, _12480_, _12471_);
  or (_12482_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  or (_12483_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_12484_, _12483_, _12482_);
  and (_12485_, _12484_, _08267_);
  or (_12486_, _12485_, _08286_);
  or (_12487_, _12486_, _12481_);
  or (_12488_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  or (_12489_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_12490_, _12489_, _12488_);
  and (_12491_, _12490_, _08279_);
  or (_12492_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  or (_12493_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_12494_, _12493_, _12492_);
  and (_12495_, _12494_, _08260_);
  or (_12496_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  or (_12497_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_12498_, _12497_, _12496_);
  and (_12499_, _12498_, _08257_);
  or (_12500_, _12499_, _12495_);
  or (_12501_, _12500_, _12491_);
  or (_12502_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  or (_12503_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_12504_, _12503_, _12502_);
  and (_12505_, _12504_, _08267_);
  or (_12506_, _12505_, _08243_);
  or (_12507_, _12506_, _12501_);
  and (_12508_, _12507_, _12487_);
  and (_12509_, _12508_, _08311_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _12509_, _12466_);
  and (_12510_, _08362_, word_in[3]);
  or (_12511_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  or (_12512_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_12513_, _12512_, _12511_);
  and (_12514_, _12513_, _08279_);
  or (_12515_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  or (_12516_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_12517_, _12516_, _12515_);
  and (_12518_, _12517_, _08260_);
  or (_12519_, _12518_, _12514_);
  or (_12521_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  or (_12522_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_12524_, _12522_, _12521_);
  and (_12525_, _12524_, _08267_);
  or (_12526_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  or (_12527_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_12528_, _12527_, _12526_);
  and (_12529_, _12528_, _08257_);
  or (_12530_, _12529_, _12525_);
  or (_12531_, _12530_, _12519_);
  and (_12532_, _12531_, _08243_);
  or (_12533_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  or (_12534_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_12535_, _12534_, _12533_);
  and (_12536_, _12535_, _08260_);
  or (_12537_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  or (_12538_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_12539_, _12538_, _12537_);
  and (_12540_, _12539_, _08279_);
  or (_12541_, _12540_, _12536_);
  or (_12542_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  or (_12543_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_12544_, _12543_, _12542_);
  and (_12545_, _12544_, _08267_);
  or (_12546_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  or (_12547_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_12548_, _12547_, _12546_);
  and (_12549_, _12548_, _08257_);
  or (_12550_, _12549_, _12545_);
  or (_12551_, _12550_, _12541_);
  and (_12552_, _12551_, _08286_);
  or (_12553_, _12552_, _12532_);
  and (_12554_, _12553_, _08311_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _12554_, _12510_);
  and (_12555_, _08362_, word_in[4]);
  or (_12556_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or (_12557_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_12558_, _12557_, _12556_);
  and (_12559_, _12558_, _08279_);
  or (_12560_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or (_12561_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_12562_, _12561_, _12560_);
  and (_12563_, _12562_, _08257_);
  or (_12564_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  or (_12565_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_12566_, _12565_, _12564_);
  and (_12567_, _12566_, _08260_);
  or (_12568_, _12567_, _12563_);
  or (_12569_, _12568_, _12559_);
  or (_12570_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  or (_12571_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_12572_, _12571_, _12570_);
  and (_12573_, _12572_, _08267_);
  or (_12574_, _12573_, _08286_);
  or (_12575_, _12574_, _12569_);
  or (_12576_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or (_12577_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_12578_, _12577_, _12576_);
  and (_12579_, _12578_, _08279_);
  or (_12580_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  or (_12581_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_12582_, _12581_, _12580_);
  and (_12583_, _12582_, _08260_);
  or (_12584_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  or (_12585_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_12586_, _12585_, _12584_);
  and (_12587_, _12586_, _08257_);
  or (_12588_, _12587_, _12583_);
  or (_12589_, _12588_, _12579_);
  or (_12590_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  or (_12591_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_12592_, _12591_, _12590_);
  and (_12593_, _12592_, _08267_);
  or (_12594_, _12593_, _08243_);
  or (_12595_, _12594_, _12589_);
  and (_12596_, _12595_, _12575_);
  and (_12597_, _12596_, _08311_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _12597_, _12555_);
  and (_12599_, _08362_, word_in[5]);
  or (_12600_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  or (_12601_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_12602_, _12601_, _12600_);
  and (_12603_, _12602_, _08279_);
  or (_12604_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  or (_12605_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_12606_, _12605_, _12604_);
  and (_12607_, _12606_, _08260_);
  or (_12608_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  or (_12609_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_12610_, _12609_, _12608_);
  and (_12611_, _12610_, _08257_);
  or (_12612_, _12611_, _12607_);
  or (_12613_, _12612_, _12603_);
  or (_12614_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  or (_12615_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_12616_, _12615_, _12614_);
  and (_12617_, _12616_, _08267_);
  or (_12618_, _12617_, _08286_);
  or (_12619_, _12618_, _12613_);
  or (_12620_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or (_12621_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_12622_, _12621_, _12620_);
  and (_12623_, _12622_, _08279_);
  or (_12624_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  or (_12625_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_12626_, _12625_, _12624_);
  and (_12627_, _12626_, _08260_);
  or (_12628_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or (_12629_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_12630_, _12629_, _12628_);
  and (_12631_, _12630_, _08257_);
  or (_12632_, _12631_, _12627_);
  or (_12633_, _12632_, _12623_);
  or (_12634_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  or (_12635_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_12636_, _12635_, _12634_);
  and (_12637_, _12636_, _08267_);
  or (_12638_, _12637_, _08243_);
  or (_12639_, _12638_, _12633_);
  and (_12640_, _12639_, _12619_);
  and (_12641_, _12640_, _08311_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _12641_, _12599_);
  and (_12642_, _08362_, word_in[6]);
  or (_12643_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  or (_12644_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_12645_, _12644_, _12643_);
  and (_12646_, _12645_, _08260_);
  or (_12647_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  or (_12648_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_12649_, _12648_, _12647_);
  and (_12650_, _12649_, _08257_);
  or (_12651_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or (_12652_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_12653_, _12652_, _12651_);
  and (_12654_, _12653_, _08279_);
  or (_12655_, _12654_, _12650_);
  or (_12656_, _12655_, _12646_);
  or (_12657_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  or (_12658_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_12659_, _12658_, _12657_);
  and (_12660_, _12659_, _08267_);
  or (_12661_, _12660_, _08286_);
  or (_12662_, _12661_, _12656_);
  or (_12663_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  or (_12664_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_12665_, _12664_, _12663_);
  and (_12666_, _12665_, _08260_);
  or (_12667_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or (_12668_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_12669_, _12668_, _12667_);
  and (_12670_, _12669_, _08279_);
  or (_12671_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or (_12672_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_12673_, _12672_, _12671_);
  and (_12674_, _12673_, _08257_);
  or (_12675_, _12674_, _12670_);
  or (_12676_, _12675_, _12666_);
  or (_12677_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  or (_12678_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_12679_, _12678_, _12677_);
  and (_12680_, _12679_, _08267_);
  or (_12681_, _12680_, _08243_);
  or (_12682_, _12681_, _12676_);
  and (_12683_, _12682_, _12662_);
  and (_12684_, _12683_, _08311_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _12684_, _12642_);
  nor (_12685_, _09148_, _09146_);
  nor (_12686_, _12685_, _09149_);
  or (_12687_, _12686_, _09039_);
  or (_12688_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_12689_, _12688_, _05605_);
  and (_12690_, _12689_, _12687_);
  and (_12691_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_12692_, _12691_, _12690_);
  and (_11435_, _12692_, _05552_);
  or (_12693_, _09145_, _09102_);
  nor (_12694_, _09039_, _09146_);
  and (_12695_, _12694_, _12693_);
  nor (_12696_, _09038_, _06588_);
  or (_12697_, _12696_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_12698_, _12697_, _12695_);
  or (_12699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _05605_);
  and (_12700_, _12699_, _05552_);
  and (_11438_, _12700_, _12698_);
  and (_12701_, _08439_, word_in[8]);
  or (_12702_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  or (_12703_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_12704_, _12703_, _12702_);
  and (_12705_, _12704_, _08441_);
  or (_12706_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or (_12707_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_12708_, _12707_, _12706_);
  and (_12709_, _12708_, _08440_);
  or (_12710_, _12709_, _12705_);
  and (_12711_, _12710_, _08402_);
  or (_12712_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  or (_12713_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_12714_, _12713_, _12712_);
  and (_12715_, _12714_, _08441_);
  or (_12716_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  or (_12717_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_12718_, _12717_, _12716_);
  and (_12719_, _12718_, _08440_);
  nor (_12720_, _12719_, _12715_);
  nor (_12721_, _12720_, _08406_);
  or (_12722_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  or (_12723_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_12724_, _12723_, _12722_);
  and (_12725_, _12724_, _08441_);
  or (_12726_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  or (_12727_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_12728_, _12727_, _12726_);
  and (_12729_, _12728_, _08440_);
  or (_12730_, _12729_, _12725_);
  and (_12731_, _12730_, _08467_);
  or (_12732_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  or (_12733_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_12734_, _12733_, _12732_);
  and (_12735_, _12734_, _08441_);
  or (_12736_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or (_12737_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_12738_, _12737_, _12736_);
  and (_12739_, _12738_, _08440_);
  or (_12740_, _12739_, _12735_);
  and (_12741_, _12740_, _08480_);
  or (_12742_, _12741_, _12731_);
  or (_12743_, _12742_, _12721_);
  nor (_12744_, _12743_, _12711_);
  nor (_12745_, _12744_, _08439_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _12745_, _12701_);
  and (_12746_, _08439_, word_in[9]);
  or (_12747_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  or (_12748_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_12749_, _12748_, _12747_);
  and (_12750_, _12749_, _08441_);
  or (_12751_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  or (_12752_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_12753_, _12752_, _12751_);
  and (_12754_, _12753_, _08440_);
  or (_12755_, _12754_, _12750_);
  and (_12756_, _12755_, _08402_);
  or (_12757_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  or (_12758_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_12759_, _12758_, _12757_);
  and (_12760_, _12759_, _08441_);
  or (_12761_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or (_12762_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_12763_, _12762_, _12761_);
  and (_12764_, _12763_, _08440_);
  nor (_12765_, _12764_, _12760_);
  nor (_12766_, _12765_, _08406_);
  or (_12767_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  or (_12768_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_12769_, _12768_, _12767_);
  and (_12770_, _12769_, _08441_);
  or (_12771_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  or (_12773_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_12774_, _12773_, _12771_);
  and (_12775_, _12774_, _08440_);
  or (_12776_, _12775_, _12770_);
  and (_12777_, _12776_, _08467_);
  or (_12778_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  or (_12779_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_12780_, _12779_, _12778_);
  and (_12781_, _12780_, _08441_);
  or (_12782_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  or (_12783_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_12784_, _12783_, _12782_);
  and (_12785_, _12784_, _08440_);
  or (_12786_, _12785_, _12781_);
  and (_12787_, _12786_, _08480_);
  or (_12788_, _12787_, _12777_);
  or (_12789_, _12788_, _12766_);
  nor (_12790_, _12789_, _12756_);
  nor (_12791_, _12790_, _08439_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _12791_, _12746_);
  and (_12792_, _08439_, word_in[10]);
  or (_12793_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  or (_12794_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_12795_, _12794_, _12793_);
  and (_12796_, _12795_, _08441_);
  or (_12797_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  or (_12798_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_12799_, _12798_, _12797_);
  and (_12800_, _12799_, _08440_);
  or (_12801_, _12800_, _12796_);
  and (_12802_, _12801_, _08402_);
  or (_12803_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  or (_12804_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_12805_, _12804_, _12803_);
  and (_12806_, _12805_, _08441_);
  or (_12808_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  or (_12809_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_12810_, _12809_, _12808_);
  and (_12811_, _12810_, _08440_);
  nor (_12812_, _12811_, _12806_);
  nor (_12813_, _12812_, _08406_);
  or (_12814_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  or (_12815_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_12816_, _12815_, _12814_);
  and (_12817_, _12816_, _08441_);
  or (_12818_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  or (_12819_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_12820_, _12819_, _12818_);
  and (_12821_, _12820_, _08440_);
  or (_12822_, _12821_, _12817_);
  and (_12823_, _12822_, _08467_);
  or (_12824_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  or (_12825_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_12826_, _12825_, _12824_);
  and (_12827_, _12826_, _08441_);
  or (_12828_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  or (_12829_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_12830_, _12829_, _12828_);
  and (_12831_, _12830_, _08440_);
  or (_12832_, _12831_, _12827_);
  and (_12833_, _12832_, _08480_);
  or (_12834_, _12833_, _12823_);
  or (_12835_, _12834_, _12813_);
  nor (_12836_, _12835_, _12802_);
  nor (_12837_, _12836_, _08439_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _12837_, _12792_);
  and (_12838_, _08439_, word_in[11]);
  or (_12839_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  or (_12840_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_12841_, _12840_, _12839_);
  and (_12842_, _12841_, _08441_);
  or (_12843_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  or (_12844_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_12845_, _12844_, _12843_);
  and (_12846_, _12845_, _08440_);
  or (_12847_, _12846_, _12842_);
  and (_12848_, _12847_, _08402_);
  or (_12849_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  or (_12850_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_12851_, _12850_, _12849_);
  and (_12852_, _12851_, _08441_);
  or (_12853_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  or (_12854_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_12855_, _12854_, _12853_);
  and (_12856_, _12855_, _08440_);
  nor (_12857_, _12856_, _12852_);
  nor (_12858_, _12857_, _08406_);
  or (_12859_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  or (_12860_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_12861_, _12860_, _12859_);
  and (_12862_, _12861_, _08441_);
  or (_12863_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  or (_12864_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_12865_, _12864_, _12863_);
  and (_12866_, _12865_, _08440_);
  or (_12867_, _12866_, _12862_);
  and (_12868_, _12867_, _08467_);
  or (_12869_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  or (_12870_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_12871_, _12870_, _12869_);
  and (_12872_, _12871_, _08441_);
  or (_12873_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  or (_12874_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_12875_, _12874_, _12873_);
  and (_12876_, _12875_, _08440_);
  or (_12877_, _12876_, _12872_);
  and (_12878_, _12877_, _08480_);
  or (_12879_, _12878_, _12868_);
  or (_12880_, _12879_, _12858_);
  nor (_12881_, _12880_, _12848_);
  nor (_12882_, _12881_, _08439_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _12882_, _12838_);
  and (_12883_, _08439_, word_in[12]);
  or (_12884_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  or (_12885_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_12886_, _12885_, _12884_);
  and (_12887_, _12886_, _08441_);
  or (_12888_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or (_12889_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_12890_, _12889_, _12888_);
  and (_12891_, _12890_, _08440_);
  or (_12892_, _12891_, _12887_);
  and (_12893_, _12892_, _08402_);
  or (_12894_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  or (_12895_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_12896_, _12895_, _12894_);
  and (_12897_, _12896_, _08441_);
  or (_12898_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  or (_12899_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_12900_, _12899_, _12898_);
  and (_12901_, _12900_, _08440_);
  nor (_12902_, _12901_, _12897_);
  nor (_12903_, _12902_, _08406_);
  or (_12904_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  or (_12905_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_12906_, _12905_, _12904_);
  and (_12907_, _12906_, _08441_);
  or (_12908_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or (_12909_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_12910_, _12909_, _12908_);
  and (_12911_, _12910_, _08440_);
  or (_12912_, _12911_, _12907_);
  and (_12913_, _12912_, _08467_);
  or (_12914_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  or (_12915_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_12916_, _12915_, _12914_);
  and (_12917_, _12916_, _08441_);
  or (_12918_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or (_12919_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_12920_, _12919_, _12918_);
  and (_12921_, _12920_, _08440_);
  or (_12922_, _12921_, _12917_);
  and (_12923_, _12922_, _08480_);
  or (_12924_, _12923_, _12913_);
  or (_12925_, _12924_, _12903_);
  nor (_12926_, _12925_, _12893_);
  nor (_12927_, _12926_, _08439_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _12927_, _12883_);
  and (_12928_, _08439_, word_in[13]);
  or (_12929_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  or (_12930_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_12931_, _12930_, _12929_);
  and (_12932_, _12931_, _08441_);
  or (_12933_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  or (_12934_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_12935_, _12934_, _12933_);
  and (_12936_, _12935_, _08440_);
  or (_12937_, _12936_, _12932_);
  and (_12938_, _12937_, _08402_);
  or (_12939_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or (_12940_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_12941_, _12940_, _12939_);
  and (_12942_, _12941_, _08441_);
  or (_12943_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  or (_12944_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_12945_, _12944_, _12943_);
  and (_12946_, _12945_, _08440_);
  nor (_12947_, _12946_, _12942_);
  nor (_12948_, _12947_, _08406_);
  or (_12949_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  or (_12950_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_12951_, _12950_, _12949_);
  and (_12952_, _12951_, _08441_);
  or (_12953_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  or (_12954_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_12955_, _12954_, _12953_);
  and (_12956_, _12955_, _08440_);
  or (_12957_, _12956_, _12952_);
  and (_12958_, _12957_, _08467_);
  or (_12959_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  or (_12960_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_12961_, _12960_, _12959_);
  and (_12962_, _12961_, _08441_);
  or (_12963_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  or (_12964_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_12965_, _12964_, _12963_);
  and (_12966_, _12965_, _08440_);
  or (_12967_, _12966_, _12962_);
  and (_12968_, _12967_, _08480_);
  or (_12969_, _12968_, _12958_);
  or (_12970_, _12969_, _12948_);
  nor (_12971_, _12970_, _12938_);
  nor (_12972_, _12971_, _08439_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _12972_, _12928_);
  and (_12973_, _08439_, word_in[14]);
  or (_12974_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or (_12975_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_12976_, _12975_, _12974_);
  and (_12977_, _12976_, _08441_);
  or (_12978_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or (_12979_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_12980_, _12979_, _12978_);
  and (_12981_, _12980_, _08440_);
  or (_12982_, _12981_, _12977_);
  and (_12983_, _12982_, _08402_);
  or (_12984_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  or (_12985_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_12986_, _12985_, _12984_);
  and (_12987_, _12986_, _08441_);
  or (_12988_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or (_12989_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_12990_, _12989_, _12988_);
  and (_12991_, _12990_, _08440_);
  nor (_12992_, _12991_, _12987_);
  nor (_12993_, _12992_, _08406_);
  or (_12994_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or (_12995_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_12996_, _12995_, _12994_);
  and (_12997_, _12996_, _08441_);
  or (_12998_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or (_12999_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_13000_, _12999_, _12998_);
  and (_13001_, _13000_, _08440_);
  or (_13002_, _13001_, _12997_);
  and (_13003_, _13002_, _08467_);
  or (_13004_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or (_13005_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_13006_, _13005_, _13004_);
  and (_13007_, _13006_, _08441_);
  or (_13008_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or (_13009_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_13010_, _13009_, _13008_);
  and (_13011_, _13010_, _08440_);
  or (_13012_, _13011_, _13007_);
  and (_13013_, _13012_, _08480_);
  or (_13014_, _13013_, _13003_);
  or (_13015_, _13014_, _12993_);
  nor (_13016_, _13015_, _12983_);
  nor (_13017_, _13016_, _08439_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13017_, _12973_);
  and (_13018_, _08533_, word_in[16]);
  and (_13019_, _12395_, _08257_);
  and (_13020_, _12389_, _08260_);
  or (_13021_, _13020_, _13019_);
  and (_13022_, _12384_, _08279_);
  and (_13023_, _12379_, _08267_);
  or (_13024_, _13023_, _13022_);
  or (_13025_, _13024_, _13021_);
  or (_13026_, _13025_, _08502_);
  and (_13027_, _12409_, _08260_);
  and (_13028_, _12401_, _08267_);
  or (_13029_, _13028_, _13027_);
  and (_13030_, _12415_, _08257_);
  and (_13031_, _12405_, _08279_);
  or (_13032_, _13031_, _13030_);
  nor (_13033_, _13032_, _13029_);
  nand (_13034_, _13033_, _08502_);
  nand (_13035_, _13034_, _13026_);
  nor (_13036_, _13035_, _08533_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13036_, _13018_);
  and (_13037_, _08533_, word_in[17]);
  and (_13038_, _12428_, _08279_);
  and (_13039_, _12424_, _08267_);
  or (_13040_, _13039_, _13038_);
  and (_13041_, _12438_, _08257_);
  and (_13042_, _12432_, _08260_);
  or (_13043_, _13042_, _13041_);
  or (_13044_, _13043_, _13040_);
  or (_13045_, _13044_, _08502_);
  and (_13046_, _12460_, _08257_);
  and (_13047_, _12449_, _08279_);
  or (_13048_, _13047_, _13046_);
  and (_13049_, _12453_, _08260_);
  and (_13050_, _12445_, _08267_);
  or (_13051_, _13050_, _13049_);
  nor (_13052_, _13051_, _13048_);
  nand (_13053_, _13052_, _08502_);
  nand (_13054_, _13053_, _13045_);
  nor (_13055_, _13054_, _08533_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13055_, _13037_);
  and (_13056_, _08533_, word_in[18]);
  and (_13057_, _12484_, _08257_);
  and (_13058_, _12478_, _08260_);
  or (_13059_, _13058_, _13057_);
  and (_13060_, _12474_, _08279_);
  and (_13061_, _12470_, _08267_);
  or (_13062_, _13061_, _13060_);
  nor (_13063_, _13062_, _13059_);
  nor (_13064_, _13063_, _08502_);
  and (_13065_, _12504_, _08257_);
  and (_13066_, _12498_, _08260_);
  or (_13067_, _13066_, _13065_);
  and (_13068_, _12494_, _08279_);
  and (_13069_, _12490_, _08267_);
  or (_13070_, _13069_, _13068_);
  or (_13071_, _13070_, _13067_);
  and (_13072_, _13071_, _08502_);
  nor (_13073_, _13072_, _13064_);
  nor (_13074_, _13073_, _08533_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13074_, _13056_);
  and (_13075_, _08533_, word_in[19]);
  and (_13076_, _12524_, _08257_);
  and (_13077_, _12517_, _08279_);
  or (_13078_, _13077_, _13076_);
  and (_13079_, _12528_, _08260_);
  and (_13080_, _12513_, _08267_);
  or (_13081_, _13080_, _13079_);
  or (_13082_, _13081_, _13078_);
  or (_13083_, _13082_, _08502_);
  and (_13084_, _12535_, _08279_);
  and (_13085_, _12539_, _08267_);
  or (_13086_, _13085_, _13084_);
  and (_13087_, _12544_, _08257_);
  and (_13088_, _12548_, _08260_);
  or (_13089_, _13088_, _13087_);
  nor (_13090_, _13089_, _13086_);
  nand (_13091_, _13090_, _08502_);
  nand (_13092_, _13091_, _13083_);
  nor (_13093_, _13092_, _08533_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13093_, _13075_);
  and (_13094_, _08533_, word_in[20]);
  and (_13095_, _12572_, _08257_);
  and (_13096_, _12566_, _08279_);
  or (_13097_, _13096_, _13095_);
  and (_13098_, _12562_, _08260_);
  and (_13099_, _12558_, _08267_);
  or (_13100_, _13099_, _13098_);
  or (_13101_, _13100_, _13097_);
  or (_13102_, _13101_, _08502_);
  and (_13103_, _12582_, _08279_);
  and (_13104_, _12578_, _08267_);
  or (_13105_, _13104_, _13103_);
  and (_13107_, _12592_, _08257_);
  and (_13108_, _12586_, _08260_);
  or (_13110_, _13108_, _13107_);
  nor (_13111_, _13110_, _13105_);
  nand (_13112_, _13111_, _08502_);
  nand (_13113_, _13112_, _13102_);
  nor (_13114_, _13113_, _08533_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13114_, _13094_);
  and (_13115_, _08533_, word_in[21]);
  and (_13116_, _12610_, _08260_);
  and (_13117_, _12616_, _08257_);
  or (_13118_, _13117_, _13116_);
  and (_13119_, _12606_, _08279_);
  and (_13120_, _12602_, _08286_);
  or (_13121_, _13120_, _13119_);
  or (_13122_, _13121_, _13118_);
  or (_13123_, _13122_, _08502_);
  and (_13124_, _12626_, _08279_);
  and (_13125_, _12622_, _08267_);
  or (_13126_, _13125_, _13124_);
  and (_13127_, _12636_, _08257_);
  and (_13128_, _12630_, _08260_);
  or (_13130_, _13128_, _13127_);
  nor (_13131_, _13130_, _13126_);
  nand (_13133_, _13131_, _08502_);
  nand (_13134_, _13133_, _13123_);
  nor (_13136_, _13134_, _08533_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13136_, _13115_);
  and (_13137_, _08533_, word_in[22]);
  and (_13138_, _12659_, _08257_);
  and (_13140_, _12645_, _08279_);
  or (_13141_, _13140_, _13138_);
  and (_13143_, _12649_, _08260_);
  and (_13144_, _12653_, _08267_);
  or (_13145_, _13144_, _13143_);
  or (_13146_, _13145_, _13141_);
  or (_13147_, _13146_, _08502_);
  and (_13148_, _12679_, _08257_);
  and (_13149_, _12665_, _08279_);
  or (_13151_, _13149_, _13148_);
  and (_13152_, _12673_, _08260_);
  and (_13153_, _12669_, _08267_);
  or (_13155_, _13153_, _13152_);
  nor (_13156_, _13155_, _13151_);
  nand (_13158_, _13156_, _08502_);
  nand (_13159_, _13158_, _13147_);
  nor (_13160_, _13159_, _08533_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13160_, _13137_);
  and (_13161_, _08595_, word_in[24]);
  and (_13162_, _12708_, _08441_);
  and (_13164_, _12704_, _08440_);
  or (_13165_, _13164_, _13162_);
  and (_13166_, _13165_, _08567_);
  and (_13168_, _12718_, _08441_);
  and (_13169_, _12714_, _08440_);
  or (_13170_, _13169_, _13168_);
  and (_13171_, _13170_, _08572_);
  and (_13172_, _12728_, _08441_);
  and (_13173_, _12724_, _08440_);
  or (_13174_, _13173_, _13172_);
  and (_13176_, _13174_, _08607_);
  and (_13177_, _12738_, _08441_);
  and (_13178_, _12734_, _08440_);
  or (_13179_, _13178_, _13177_);
  and (_13180_, _13179_, _08613_);
  or (_13181_, _13180_, _13176_);
  or (_13182_, _13181_, _13171_);
  nor (_13183_, _13182_, _13166_);
  nor (_13184_, _13183_, _08595_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13184_, _13161_);
  and (_13185_, _08595_, word_in[25]);
  and (_13186_, _12753_, _08441_);
  and (_13187_, _12749_, _08440_);
  or (_13188_, _13187_, _13186_);
  and (_13189_, _13188_, _08567_);
  and (_13190_, _12763_, _08441_);
  and (_13192_, _12759_, _08440_);
  or (_13193_, _13192_, _13190_);
  and (_13195_, _13193_, _08572_);
  and (_13196_, _12774_, _08441_);
  and (_13198_, _12769_, _08440_);
  or (_13199_, _13198_, _13196_);
  and (_13200_, _13199_, _08607_);
  and (_13201_, _12784_, _08441_);
  and (_13202_, _12780_, _08440_);
  or (_13204_, _13202_, _13201_);
  and (_13205_, _13204_, _08613_);
  or (_13207_, _13205_, _13200_);
  or (_13208_, _13207_, _13195_);
  nor (_13210_, _13208_, _13189_);
  nor (_13211_, _13210_, _08595_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13211_, _13185_);
  and (_13213_, _08595_, word_in[26]);
  and (_13214_, _12799_, _08441_);
  and (_13216_, _12795_, _08440_);
  or (_13217_, _13216_, _13214_);
  and (_13218_, _13217_, _08567_);
  and (_13220_, _12810_, _08441_);
  and (_13221_, _12805_, _08440_);
  or (_13223_, _13221_, _13220_);
  and (_13224_, _13223_, _08572_);
  and (_13225_, _12820_, _08441_);
  and (_13226_, _12816_, _08440_);
  or (_13227_, _13226_, _13225_);
  and (_13228_, _13227_, _08607_);
  and (_13229_, _12830_, _08441_);
  and (_13230_, _12826_, _08440_);
  or (_13231_, _13230_, _13229_);
  and (_13232_, _13231_, _08613_);
  or (_13233_, _13232_, _13228_);
  or (_13234_, _13233_, _13224_);
  nor (_13235_, _13234_, _13218_);
  nor (_13236_, _13235_, _08595_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13236_, _13213_);
  and (_13238_, _08595_, word_in[27]);
  and (_13239_, _12855_, _08441_);
  and (_13240_, _12851_, _08440_);
  or (_13241_, _13240_, _13239_);
  and (_13243_, _13241_, _08572_);
  and (_13244_, _12845_, _08441_);
  and (_13246_, _12841_, _08440_);
  or (_13247_, _13246_, _13244_);
  and (_13248_, _13247_, _08567_);
  and (_13249_, _12865_, _08441_);
  and (_13251_, _12861_, _08440_);
  or (_13252_, _13251_, _13249_);
  and (_13253_, _13252_, _08607_);
  and (_13254_, _12875_, _08441_);
  and (_13255_, _12871_, _08440_);
  or (_13256_, _13255_, _13254_);
  and (_13257_, _13256_, _08613_);
  or (_13258_, _13257_, _13253_);
  or (_13259_, _13258_, _13248_);
  nor (_13260_, _13259_, _13243_);
  nor (_13261_, _13260_, _08595_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13261_, _13238_);
  and (_13263_, _08595_, word_in[28]);
  and (_13264_, _12890_, _08441_);
  and (_13265_, _12886_, _08440_);
  or (_13266_, _13265_, _13264_);
  and (_13267_, _13266_, _08567_);
  and (_13268_, _12900_, _08441_);
  and (_13269_, _12896_, _08440_);
  or (_13270_, _13269_, _13268_);
  and (_13272_, _13270_, _08572_);
  and (_13273_, _12910_, _08441_);
  and (_13274_, _12906_, _08440_);
  or (_13275_, _13274_, _13273_);
  and (_13277_, _13275_, _08607_);
  and (_13278_, _12920_, _08441_);
  and (_13280_, _12916_, _08440_);
  or (_13281_, _13280_, _13278_);
  and (_13283_, _13281_, _08613_);
  or (_13284_, _13283_, _13277_);
  or (_13285_, _13284_, _13272_);
  nor (_13286_, _13285_, _13267_);
  nor (_13287_, _13286_, _08595_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13287_, _13263_);
  and (_13288_, _08595_, word_in[29]);
  and (_13289_, _12945_, _08441_);
  and (_13290_, _12941_, _08440_);
  or (_13291_, _13290_, _13289_);
  and (_13292_, _13291_, _08572_);
  and (_13294_, _12935_, _08441_);
  and (_13295_, _12931_, _08440_);
  or (_13297_, _13295_, _13294_);
  and (_13298_, _13297_, _08567_);
  and (_13299_, _12955_, _08441_);
  and (_13300_, _12951_, _08440_);
  or (_13302_, _13300_, _13299_);
  and (_13303_, _13302_, _08607_);
  and (_13304_, _12965_, _08441_);
  and (_13305_, _12961_, _08440_);
  or (_13306_, _13305_, _13304_);
  and (_13307_, _13306_, _08613_);
  or (_13308_, _13307_, _13303_);
  or (_13309_, _13308_, _13298_);
  nor (_13310_, _13309_, _13292_);
  nor (_13311_, _13310_, _08595_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13311_, _13288_);
  and (_13312_, _08595_, word_in[30]);
  and (_13313_, _12980_, _08441_);
  and (_13314_, _12976_, _08440_);
  or (_13315_, _13314_, _13313_);
  and (_13316_, _13315_, _08567_);
  and (_13317_, _12990_, _08441_);
  and (_13318_, _12986_, _08440_);
  or (_13319_, _13318_, _13317_);
  and (_13320_, _13319_, _08572_);
  and (_13321_, _13000_, _08441_);
  and (_13322_, _12996_, _08440_);
  or (_13323_, _13322_, _13321_);
  and (_13324_, _13323_, _08607_);
  and (_13325_, _13010_, _08441_);
  and (_13326_, _13006_, _08440_);
  or (_13327_, _13326_, _13325_);
  and (_13328_, _13327_, _08613_);
  or (_13329_, _13328_, _13324_);
  or (_13331_, _13329_, _13320_);
  nor (_13332_, _13331_, _13316_);
  nor (_13333_, _13332_, _08595_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13333_, _13312_);
  and (_13334_, _05552_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_11498_, _13334_, _05671_);
  and (_11504_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _05552_);
  nor (_11517_, _11469_, rst);
  or (_13335_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand (_13336_, _05550_, _11609_);
  and (_13337_, _13336_, _05552_);
  and (_11551_, _13337_, _13335_);
  or (_13339_, _09144_, _09105_);
  nor (_13341_, _09039_, _09145_);
  and (_13342_, _13341_, _13339_);
  nor (_13343_, _09038_, _06489_);
  or (_13344_, _13343_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_13345_, _13344_, _13342_);
  or (_13346_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_13347_, _13346_, _05552_);
  and (_11554_, _13347_, _13345_);
  nor (_13349_, _09142_, _09139_);
  nor (_13350_, _13349_, _09143_);
  or (_13352_, _13350_, _09039_);
  or (_13353_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_13354_, _13353_, _07933_);
  and (_13355_, _13354_, _13352_);
  and (_13356_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_13357_, _13356_, _05552_);
  or (_11588_, _13357_, _13355_);
  nand (_13358_, _07711_, _06973_);
  and (_13359_, _08048_, _06060_);
  nor (_13360_, _06060_, _06201_);
  nor (_13361_, _13360_, _13359_);
  or (_13362_, _13361_, _08924_);
  and (_13363_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_13365_, _13363_, _07260_);
  and (_13366_, _13365_, _13362_);
  nand (_13367_, _13366_, _13358_);
  or (_13368_, _08228_, _07261_);
  and (_13369_, _13368_, _13367_);
  and (_11659_, _13369_, _05552_);
  nand (_13371_, _06949_, _06560_);
  or (_13372_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_13373_, _13372_, _05552_);
  and (_11681_, _13373_, _13371_);
  nor (_13374_, _07211_, _06330_);
  and (_13375_, _07211_, _06330_);
  or (_13377_, _13375_, _13374_);
  and (_11685_, _13377_, _05552_);
  and (_13379_, _12299_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_13380_, _10898_, _05820_);
  and (_13381_, _13380_, _10905_);
  or (_13382_, _13381_, _10941_);
  or (_13383_, _10943_, _10899_);
  or (_13384_, _13383_, _13382_);
  or (_13385_, _11174_, _12282_);
  and (_13386_, _06567_, _05830_);
  or (_13387_, _13386_, _12307_);
  or (_13389_, _13387_, _13385_);
  or (_13390_, _13389_, _10927_);
  or (_13391_, _13390_, _13384_);
  or (_13392_, _11160_, _11151_);
  and (_13394_, _06567_, _05846_);
  or (_13395_, _13394_, _12272_);
  or (_13397_, _13395_, _13392_);
  or (_13398_, _12328_, _11155_);
  or (_13399_, _13398_, _12291_);
  or (_13400_, _13399_, _13397_);
  or (_13401_, _13400_, _13391_);
  and (_13402_, _13401_, _06576_);
  or (_11720_, _13402_, _13379_);
  and (_11741_, _07646_, _05552_);
  nor (_13404_, _07939_, _07388_);
  and (_13405_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or (_13407_, _13405_, _13404_);
  and (_11748_, _13407_, _05552_);
  and (_13408_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_13409_, _07976_, _07937_);
  or (_13410_, _13409_, _13408_);
  and (_11755_, _13410_, _05552_);
  and (_13411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _05556_);
  and (_13412_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_13413_, _13412_, _13411_);
  and (_11758_, _13413_, _05552_);
  not (_13414_, _11774_);
  or (_13415_, _12037_, _11828_);
  or (_13416_, _12029_, _12032_);
  and (_13417_, _13416_, _13415_);
  nor (_13418_, _13417_, _06487_);
  and (_13419_, _13417_, _06487_);
  or (_13420_, _13419_, _13418_);
  and (_13421_, _13420_, _12161_);
  and (_13422_, _11811_, _07574_);
  and (_13423_, _11784_, _07600_);
  nor (_13424_, _11805_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_13425_, _13424_, _11806_);
  and (_13426_, _13425_, _11792_);
  and (_13427_, _11780_, _11391_);
  and (_13428_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_13429_, _13428_, _13427_);
  or (_13430_, _13429_, _13426_);
  or (_13431_, _13430_, _13423_);
  or (_13432_, _13431_, _13422_);
  or (_13433_, _13432_, _13421_);
  or (_13434_, _13433_, _13414_);
  nor (_13435_, _12071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_13436_, _13435_, _12072_);
  or (_13437_, _13436_, _11774_);
  and (_13438_, _13437_, _05552_);
  and (_11798_, _13438_, _13434_);
  nand (_13439_, _12028_, _11828_);
  or (_13440_, _12036_, _11828_);
  and (_13441_, _13440_, _13439_);
  nand (_13442_, _13441_, _06085_);
  or (_13443_, _13441_, _06085_);
  and (_13444_, _13443_, _12161_);
  and (_13445_, _13444_, _13442_);
  and (_13446_, _11811_, _07635_);
  and (_13447_, _11784_, _07663_);
  nor (_13448_, _11804_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_13449_, _13448_, _11805_);
  and (_13450_, _13449_, _11792_);
  and (_13451_, _11780_, _11449_);
  and (_13452_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_13453_, _13452_, _13451_);
  or (_13454_, _13453_, _13450_);
  nor (_13455_, _13454_, _13447_);
  nand (_13456_, _13455_, _11774_);
  or (_13457_, _13456_, _13446_);
  or (_13458_, _13457_, _13445_);
  nor (_13459_, _12069_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_13460_, _13459_, _12071_);
  or (_13461_, _13460_, _11774_);
  and (_13462_, _13461_, _05552_);
  and (_11826_, _13462_, _13458_);
  not (_13463_, _11650_);
  and (_13464_, _11704_, _13463_);
  not (_13465_, _11509_);
  not (_13466_, _11452_);
  not (_13467_, _11335_);
  nand (_13468_, _11395_, _13467_);
  or (_13469_, _13468_, _13466_);
  or (_13471_, _13469_, _13465_);
  not (_13472_, _13471_);
  and (_13473_, _11763_, _11279_);
  and (_13474_, _13473_, _13472_);
  and (_13475_, _13474_, _13464_);
  and (_13476_, _13475_, _07485_);
  nor (_13477_, _13476_, rst);
  and (_13478_, _07711_, _05552_);
  or (_13479_, _13478_, _13477_);
  and (_13480_, _11704_, _11650_);
  not (_13481_, _11763_);
  nor (_13482_, _13481_, _11279_);
  and (_13484_, _13482_, _13480_);
  nor (_13485_, _11395_, _13466_);
  and (_13486_, _11509_, _13467_);
  and (_13487_, _13486_, _13485_);
  and (_13488_, _13487_, _13484_);
  nand (_13489_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor (_13491_, _11763_, _11279_);
  and (_13492_, _13491_, _13480_);
  and (_13494_, _13487_, _13492_);
  nand (_13495_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_13496_, _13495_, _13489_);
  nor (_13497_, _11704_, _13463_);
  and (_13498_, _13491_, _13497_);
  and (_13499_, _13487_, _13498_);
  nand (_13500_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_13501_, _13482_, _13464_);
  and (_13502_, _13487_, _13501_);
  nand (_13503_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_13504_, _13503_, _13500_);
  and (_13505_, _13504_, _13496_);
  and (_13507_, _13484_, _13472_);
  nand (_13508_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nor (_13509_, _11704_, _11650_);
  and (_13510_, _13482_, _13509_);
  and (_13511_, _13487_, _13510_);
  nand (_13512_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_13513_, _13512_, _13508_);
  nor (_13514_, _13468_, _11452_);
  and (_13515_, _13514_, _11509_);
  and (_13516_, _13515_, _13484_);
  nand (_13517_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_13518_, _13514_, _13465_);
  and (_13519_, _13509_, _13481_);
  and (_13520_, _13519_, _11279_);
  and (_13521_, _13520_, _13518_);
  nand (_13522_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_13523_, _13522_, _13517_);
  and (_13524_, _13523_, _13513_);
  and (_13525_, _13524_, _13505_);
  not (_13526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_13527_, _13497_, _13482_);
  nand (_13528_, _13527_, _13472_);
  or (_13529_, _13528_, _13526_);
  not (_13530_, _13510_);
  nor (_13531_, _13530_, _13471_);
  nand (_13532_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_13533_, _13532_, _13529_);
  and (_13534_, _13501_, _13472_);
  nand (_13535_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_13536_, _13498_, _13472_);
  nand (_13537_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_13538_, _13537_, _13535_);
  and (_13539_, _13538_, _13533_);
  nor (_13540_, _13469_, _11509_);
  and (_13541_, _13540_, _13527_);
  nand (_13542_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_13544_, _13484_, _13540_);
  nand (_13545_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_13546_, _13545_, _13542_);
  and (_13547_, _13492_, _13472_);
  nand (_13548_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_13549_, _13520_, _13472_);
  nand (_13550_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_13551_, _13550_, _13548_);
  and (_13552_, _13551_, _13546_);
  and (_13553_, _13552_, _13539_);
  and (_13554_, _13553_, _13525_);
  and (_13555_, _13497_, _13474_);
  nand (_13556_, _13555_, _11700_);
  and (_13557_, _13480_, _13473_);
  and (_13559_, _13557_, _13465_);
  nor (_13560_, _11395_, _11452_);
  and (_13561_, _13560_, _13467_);
  and (_13562_, _13561_, _13559_);
  nand (_13563_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_13565_, _13563_, _13556_);
  nand (_13566_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_13567_, _13509_, _13473_);
  nor (_13568_, _13567_, _13471_);
  nand (_13570_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_13571_, _13570_, _13566_);
  and (_13572_, _13571_, _13565_);
  not (_13573_, _13557_);
  nor (_13574_, _13573_, _13471_);
  and (_13575_, _12283_, _05852_);
  or (_13576_, _13575_, _05855_);
  nor (_13577_, _13576_, _11169_);
  and (_13578_, _10898_, _05854_);
  and (_13579_, _13578_, _05669_);
  nor (_13581_, _12331_, _13579_);
  and (_13582_, _13581_, _13577_);
  and (_13583_, _10909_, _10843_);
  or (_13584_, _12330_, _05811_);
  nor (_13585_, _13584_, _13583_);
  and (_13586_, _13585_, _12315_);
  and (_13588_, _13586_, _13582_);
  and (_13589_, _13588_, _12319_);
  and (_13591_, _13589_, _11159_);
  nor (_13592_, _13591_, _11085_);
  nor (_13593_, _13592_, p0_in[0]);
  not (_13594_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_13595_, _13592_, _13594_);
  nor (_13596_, _13595_, _13593_);
  nand (_13597_, _13596_, _13574_);
  and (_13598_, _13540_, _13557_);
  nor (_13599_, _13592_, p1_in[0]);
  not (_13600_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_13601_, _13592_, _13600_);
  nor (_13602_, _13601_, _13599_);
  nand (_13603_, _13602_, _13598_);
  and (_13604_, _13603_, _13597_);
  and (_13605_, _13518_, _13557_);
  nor (_13606_, _13592_, p3_in[0]);
  not (_13607_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_13608_, _13592_, _13607_);
  nor (_13609_, _13608_, _13606_);
  nand (_13610_, _13609_, _13605_);
  and (_13611_, _13515_, _13557_);
  nor (_13612_, _13592_, p2_in[0]);
  not (_13613_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_13614_, _13592_, _13613_);
  nor (_13615_, _13614_, _13612_);
  nand (_13616_, _13615_, _13611_);
  and (_13617_, _13616_, _13610_);
  and (_13618_, _13617_, _13604_);
  and (_13619_, _13618_, _13572_);
  nor (_13620_, _11509_, _11335_);
  and (_13621_, _13620_, _13485_);
  and (_13622_, _13621_, _13557_);
  nand (_13623_, _07362_, _07275_);
  nand (_13624_, _08920_, _13623_);
  or (_13625_, _08920_, _13623_);
  nand (_13626_, _13625_, _13624_);
  and (_13627_, _12189_, _06973_);
  nor (_13628_, _08057_, _06157_);
  or (_13629_, _13628_, _08062_);
  and (_13630_, _13629_, _08923_);
  and (_13631_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_13632_, _13631_, _07260_);
  or (_13633_, _13632_, _13630_);
  or (_13634_, _13633_, _13627_);
  or (_13635_, _12215_, _07261_);
  and (_13636_, _13635_, _13634_);
  and (_13637_, _07635_, _06973_);
  nand (_13638_, _08635_, _06763_);
  or (_13639_, _08635_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_13640_, _13639_, _08923_);
  and (_13641_, _13640_, _13638_);
  and (_13642_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_13643_, _13642_, _07260_);
  or (_13644_, _13643_, _13641_);
  or (_13645_, _13644_, _13637_);
  or (_13646_, _07663_, _07261_);
  and (_13647_, _13646_, _13645_);
  or (_13648_, _13647_, _13636_);
  nand (_13649_, _13647_, _13636_);
  and (_13650_, _13649_, _13648_);
  nand (_13651_, _13650_, _13626_);
  or (_13652_, _13650_, _13626_);
  nand (_13653_, _13652_, _13651_);
  nand (_13654_, _13368_, _13367_);
  nand (_13655_, _13654_, _08942_);
  or (_13656_, _13654_, _08942_);
  nand (_13657_, _13656_, _13655_);
  or (_13658_, _12137_, _12136_);
  nand (_13659_, _08144_, _06973_);
  and (_13660_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_13661_, _08013_, _06213_);
  nor (_13662_, _13661_, _08015_);
  nor (_13663_, _13662_, _08924_);
  nor (_13664_, _13663_, _13660_);
  and (_13665_, _13664_, _07261_);
  and (_13666_, _13665_, _13659_);
  and (_13667_, _08200_, _07260_);
  nor (_13668_, _13667_, _13666_);
  nand (_13669_, _13668_, _13658_);
  or (_13670_, _13668_, _13658_);
  and (_13671_, _13670_, _13669_);
  nand (_13672_, _13671_, _13657_);
  or (_13673_, _13671_, _13657_);
  nand (_13674_, _13673_, _13672_);
  nand (_13675_, _13674_, _13653_);
  or (_13676_, _13674_, _13653_);
  nand (_13677_, _13676_, _13675_);
  nand (_13678_, _13677_, _13622_);
  and (_13679_, _13557_, _11509_);
  and (_13681_, _13561_, _13679_);
  nand (_13683_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_13684_, _13683_, _13678_);
  and (_13685_, _13684_, _13619_);
  and (_13686_, _13685_, _13554_);
  and (_13687_, _13622_, _11591_);
  and (_13688_, _13509_, _13474_);
  and (_13689_, _13688_, _07485_);
  nor (_13690_, _13689_, _13687_);
  nor (_13691_, _13690_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_13692_, _13691_);
  nor (_13693_, _10859_, _05971_);
  not (_13694_, _13519_);
  and (_13695_, _13694_, _13693_);
  and (_13696_, _13695_, _11515_);
  or (_13697_, _07260_, _06965_);
  and (_13698_, _13681_, _13697_);
  nor (_13699_, _13698_, _13696_);
  and (_13700_, _13699_, _11772_);
  and (_13701_, _13700_, _13692_);
  not (_13702_, _13701_);
  nor (_13703_, _13702_, _13686_);
  not (_13704_, _13476_);
  nor (_13705_, _13494_, _13488_);
  nor (_13706_, _13502_, _13499_);
  and (_13707_, _13706_, _13705_);
  nor (_13708_, _13511_, _13507_);
  nor (_13710_, _13521_, _13516_);
  and (_13711_, _13710_, _13708_);
  and (_13712_, _13711_, _13707_);
  not (_13713_, _13528_);
  nor (_13715_, _13531_, _13713_);
  nor (_13716_, _13536_, _13534_);
  and (_13718_, _13716_, _13715_);
  nor (_13719_, _13544_, _13541_);
  nor (_13721_, _13549_, _13547_);
  and (_13722_, _13721_, _13719_);
  and (_13723_, _13722_, _13718_);
  and (_13724_, _13723_, _13712_);
  nor (_13725_, _13681_, _13622_);
  not (_13727_, _13468_);
  nand (_13728_, _13557_, _13727_);
  nor (_13729_, _13568_, _13475_);
  nor (_13730_, _13562_, _13555_);
  and (_13731_, _13730_, _13729_);
  and (_13732_, _13731_, _13728_);
  and (_13733_, _13732_, _13725_);
  nand (_13734_, _13733_, _13724_);
  nand (_13735_, _13734_, _13701_);
  nand (_13736_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_13737_, _13736_, _13704_);
  or (_13738_, _13737_, _13703_);
  and (_11841_, _13738_, _13479_);
  or (_13739_, _06948_, _06063_);
  or (_13740_, _09508_, _13739_);
  not (_13741_, _09503_);
  or (_13742_, _13741_, _06309_);
  and (_13743_, _13742_, _06068_);
  or (_13744_, _13743_, _13740_);
  and (_13745_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_13746_, _12264_, _06307_);
  or (_13747_, _13746_, _13745_);
  and (_11869_, _13747_, _05552_);
  and (_13748_, _09505_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_13749_, _09505_, _06560_);
  or (_13750_, _13749_, _13748_);
  or (_13751_, _13750_, _06955_);
  or (_13752_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_13753_, _13752_, _05552_);
  and (_11880_, _13753_, _13751_);
  and (_13754_, _07951_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_13755_, _07946_, _07949_);
  or (_13756_, _13755_, _13754_);
  and (_11882_, _13756_, _05552_);
  nand (_13757_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_13758_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand (_13759_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_13760_, _13759_, _13758_);
  nand (_13762_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand (_13763_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_13764_, _13763_, _13762_);
  and (_13765_, _13764_, _13760_);
  nand (_13766_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand (_13767_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_13768_, _13767_, _13766_);
  nand (_13769_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_13770_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_13771_, _13770_, _13769_);
  and (_13772_, _13771_, _13768_);
  and (_13773_, _13772_, _13765_);
  nand (_13774_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  not (_13775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or (_13776_, _13528_, _13775_);
  and (_13777_, _13776_, _13774_);
  nand (_13778_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_13779_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_13780_, _13779_, _13778_);
  and (_13781_, _13780_, _13777_);
  nand (_13782_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand (_13783_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_13784_, _13783_, _13782_);
  nand (_13785_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_13786_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_13787_, _13786_, _13785_);
  and (_13788_, _13787_, _13784_);
  and (_13789_, _13788_, _13781_);
  and (_13790_, _13789_, _13773_);
  nand (_13791_, _13555_, _11503_);
  nand (_13792_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_13793_, _13792_, _13791_);
  nand (_13794_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_13795_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_13796_, _13795_, _13794_);
  and (_13797_, _13796_, _13793_);
  nor (_13798_, _13592_, p2_in[4]);
  not (_13799_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_13800_, _13592_, _13799_);
  nor (_13801_, _13800_, _13798_);
  nand (_13802_, _13801_, _13611_);
  nor (_13803_, _13592_, p3_in[4]);
  not (_13804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_13805_, _13592_, _13804_);
  nor (_13806_, _13805_, _13803_);
  nand (_13807_, _13806_, _13605_);
  and (_13808_, _13807_, _13802_);
  nor (_13809_, _13592_, p0_in[4]);
  not (_13810_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_13811_, _13592_, _13810_);
  nor (_13812_, _13811_, _13809_);
  nand (_13813_, _13812_, _13574_);
  nor (_13814_, _13592_, p1_in[4]);
  not (_13815_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_13816_, _13592_, _13815_);
  nor (_13817_, _13816_, _13814_);
  nand (_13818_, _13817_, _13598_);
  and (_13819_, _13818_, _13813_);
  and (_13820_, _13819_, _13808_);
  and (_13821_, _13820_, _13797_);
  nand (_13822_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_13823_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_13824_, _13823_, _13822_);
  and (_13825_, _13824_, _13821_);
  and (_13826_, _13825_, _13790_);
  or (_13827_, _13826_, _13702_);
  and (_13828_, _13827_, _13757_);
  nand (_13829_, _13828_, _13704_);
  or (_13830_, _13704_, _12189_);
  and (_13831_, _13830_, _05552_);
  and (_11885_, _13831_, _13829_);
  nand (_13832_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_13833_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nand (_13834_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_13835_, _13834_, _13833_);
  nand (_13836_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_13837_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_13838_, _13837_, _13836_);
  and (_13839_, _13838_, _13835_);
  nand (_13840_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand (_13841_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_13842_, _13841_, _13840_);
  nand (_13843_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nand (_13844_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_13845_, _13844_, _13843_);
  and (_13846_, _13845_, _13842_);
  and (_13847_, _13846_, _13839_);
  nand (_13848_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_13849_, _13713_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_13850_, _13849_, _13848_);
  nand (_13851_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand (_13852_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00002_, _13852_, _13851_);
  and (_00003_, _00002_, _13850_);
  nand (_00004_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  nand (_00005_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_00006_, _00005_, _00004_);
  nand (_00007_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_00008_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_00009_, _00008_, _00007_);
  and (_00010_, _00009_, _00006_);
  and (_00011_, _00010_, _00003_);
  and (_00012_, _00011_, _13847_);
  nand (_00013_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand (_00014_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_00015_, _00014_, _00013_);
  nand (_00016_, _13555_, _11251_);
  nand (_00017_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00018_, _00017_, _00016_);
  and (_00019_, _00018_, _00015_);
  nor (_00020_, _13592_, p0_in[3]);
  not (_00021_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_00022_, _13592_, _00021_);
  nor (_00023_, _00022_, _00020_);
  nand (_00024_, _00023_, _13574_);
  nor (_00026_, _13592_, p1_in[3]);
  not (_00027_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00028_, _13592_, _00027_);
  nor (_00029_, _00028_, _00026_);
  nand (_00030_, _00029_, _13598_);
  and (_00031_, _00030_, _00024_);
  nor (_00032_, _13592_, p3_in[3]);
  not (_00033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_00034_, _13592_, _00033_);
  nor (_00035_, _00034_, _00032_);
  nand (_00036_, _00035_, _13605_);
  nor (_00037_, _13592_, p2_in[3]);
  not (_00038_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00039_, _13592_, _00038_);
  nor (_00040_, _00039_, _00037_);
  nand (_00041_, _00040_, _13611_);
  and (_00042_, _00041_, _00036_);
  and (_00043_, _00042_, _00031_);
  and (_00044_, _00043_, _00019_);
  nand (_00045_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand (_00046_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_00047_, _00046_, _00045_);
  and (_00048_, _00047_, _00044_);
  and (_00049_, _00048_, _00012_);
  or (_00050_, _00049_, _13702_);
  and (_00051_, _00050_, _13832_);
  nand (_00052_, _00051_, _13704_);
  or (_00053_, _13704_, _07483_);
  and (_00054_, _00053_, _05552_);
  and (_11888_, _00054_, _00052_);
  and (_00055_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_00056_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_00057_, _00056_, _00055_);
  and (_00058_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_00059_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_00061_, _00059_, _00058_);
  or (_00062_, _00061_, _00057_);
  and (_00063_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_00064_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_00065_, _00064_, _00063_);
  and (_00066_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_00067_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_00068_, _00067_, _00066_);
  or (_00069_, _00068_, _00065_);
  or (_00070_, _00069_, _00062_);
  and (_00072_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  not (_00073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_00074_, _13528_, _00073_);
  or (_00075_, _00074_, _00072_);
  and (_00077_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00078_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_00079_, _00078_, _00077_);
  or (_00080_, _00079_, _00075_);
  and (_00081_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_00082_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_00083_, _00082_, _00081_);
  and (_00084_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00086_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_00087_, _00086_, _00084_);
  or (_00088_, _00087_, _00083_);
  or (_00089_, _00088_, _00080_);
  or (_00090_, _00089_, _00070_);
  and (_00091_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00092_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00093_, _00092_, _00091_);
  and (_00094_, _13555_, _11759_);
  and (_00095_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00096_, _00095_, _00094_);
  or (_00097_, _00096_, _00093_);
  or (_00098_, _13592_, p3_in[2]);
  not (_00099_, _13592_);
  or (_00100_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_00101_, _00100_, _00098_);
  and (_00102_, _00101_, _13605_);
  or (_00103_, _13592_, p2_in[2]);
  or (_00104_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_00105_, _00104_, _00103_);
  and (_00106_, _00105_, _13611_);
  or (_00107_, _00106_, _00102_);
  or (_00108_, _13592_, p1_in[2]);
  or (_00109_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_00110_, _00109_, _00108_);
  and (_00111_, _00110_, _13598_);
  or (_00112_, _13592_, p0_in[2]);
  or (_00113_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_00114_, _00113_, _00112_);
  and (_00115_, _00114_, _13574_);
  or (_00116_, _00115_, _00111_);
  or (_00117_, _00116_, _00107_);
  or (_00118_, _00117_, _00097_);
  and (_00119_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_00120_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00121_, _00120_, _00119_);
  or (_00123_, _00121_, _00118_);
  or (_00124_, _00123_, _00090_);
  and (_00125_, _00124_, _13701_);
  and (_00126_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or (_00127_, _00126_, _00125_);
  or (_00128_, _00127_, _13476_);
  or (_00129_, _13704_, _08144_);
  and (_00130_, _00129_, _05552_);
  and (_11894_, _00130_, _00128_);
  and (_00131_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_00132_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_00133_, _00132_, _00131_);
  and (_00134_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_00135_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_00136_, _00135_, _00134_);
  or (_00137_, _00136_, _00133_);
  and (_00138_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_00139_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_00140_, _00139_, _00138_);
  and (_00141_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_00142_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_00143_, _00142_, _00141_);
  or (_00144_, _00143_, _00140_);
  or (_00145_, _00144_, _00137_);
  not (_00146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_00147_, _13528_, _00146_);
  and (_00148_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_00149_, _00148_, _00147_);
  and (_00150_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00151_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_00152_, _00151_, _00150_);
  or (_00154_, _00152_, _00149_);
  and (_00155_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_00156_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_00157_, _00156_, _00155_);
  and (_00158_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00160_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_00161_, _00160_, _00158_);
  or (_00162_, _00161_, _00157_);
  or (_00163_, _00162_, _00154_);
  or (_00164_, _00163_, _00145_);
  and (_00165_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00166_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00167_, _00166_, _00165_);
  and (_00168_, _13555_, _11627_);
  and (_00169_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_00170_, _00169_, _00168_);
  or (_00171_, _00170_, _00167_);
  or (_00172_, _13592_, p2_in[1]);
  not (_00173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nand (_00174_, _13592_, _00173_);
  and (_00175_, _00174_, _00172_);
  and (_00176_, _00175_, _13611_);
  or (_00177_, _13592_, p3_in[1]);
  or (_00178_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_00179_, _00178_, _00177_);
  and (_00180_, _00179_, _13605_);
  or (_00181_, _00180_, _00176_);
  or (_00182_, _13592_, p0_in[1]);
  or (_00183_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_00184_, _00183_, _00182_);
  and (_00185_, _00184_, _13574_);
  or (_00186_, _13592_, p1_in[1]);
  or (_00187_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_00188_, _00187_, _00186_);
  and (_00189_, _00188_, _13598_);
  or (_00190_, _00189_, _00185_);
  or (_00191_, _00190_, _00181_);
  or (_00192_, _00191_, _00171_);
  and (_00193_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_00194_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00195_, _00194_, _00193_);
  or (_00196_, _00195_, _00192_);
  or (_00197_, _00196_, _00164_);
  and (_00198_, _00197_, _13701_);
  and (_00199_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_00200_, _00199_, _00198_);
  or (_00202_, _00200_, _13476_);
  or (_00203_, _13704_, _08102_);
  and (_00204_, _00203_, _05552_);
  and (_11897_, _00204_, _00202_);
  nor (_11963_, _05646_, rst);
  or (_00207_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_00208_, _05550_, _05786_);
  and (_00209_, _00208_, _05552_);
  and (_11974_, _00209_, _00207_);
  and (_00210_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00211_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or (_00212_, _00211_, _00210_);
  and (_11981_, _00212_, _05552_);
  and (_00213_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00214_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or (_00215_, _00214_, _00213_);
  and (_11984_, _00215_, _05552_);
  or (_00216_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand (_00217_, _05550_, _11052_);
  and (_00218_, _00217_, _05552_);
  and (_11992_, _00218_, _00216_);
  nor (_12003_, _11646_, rst);
  and (_00220_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00221_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_00222_, _00221_, _00220_);
  and (_12011_, _00222_, _05552_);
  nand (_00223_, _10860_, _06527_);
  nor (_00224_, _00223_, _05971_);
  and (_00225_, _00224_, _06910_);
  or (_00226_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_00227_, _00226_, _00225_);
  nand (_00228_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_00229_, _00228_, _00225_);
  or (_00230_, _00229_, _08926_);
  and (_00231_, _00230_, _00227_);
  and (_00232_, _08990_, _06927_);
  or (_00233_, _00232_, _00231_);
  nand (_00234_, _00232_, _07975_);
  and (_00236_, _00234_, _05552_);
  and (_12023_, _00236_, _00233_);
  or (_00237_, _07668_, _07255_);
  or (_00238_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00239_, _00238_, _05552_);
  and (_12026_, _00239_, _00237_);
  nor (_12033_, _11872_, rst);
  and (_00240_, _06771_, _06525_);
  and (_00241_, _00240_, _07443_);
  nand (_00242_, _00241_, _08041_);
  or (_00243_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_00244_, _00243_, _05552_);
  and (_12042_, _00244_, _00242_);
  and (_00245_, _08989_, _06056_);
  and (_00246_, _00245_, _06927_);
  and (_00248_, _00246_, _05560_);
  and (_00249_, _00248_, _11490_);
  and (_00250_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_00252_, _00250_, _05560_);
  and (_00253_, _05573_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_00254_, _00253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_00255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_00256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_00257_, _00256_, _00255_);
  and (_00258_, _00257_, _00254_);
  nor (_00259_, _00258_, _00252_);
  not (_00260_, _00259_);
  and (_00261_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_00262_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_00263_, _00262_, _00261_);
  and (_00264_, _06524_, _06308_);
  and (_00265_, _00264_, _06927_);
  nor (_00266_, _00265_, _00263_);
  and (_00267_, _00246_, _05573_);
  not (_00268_, _00267_);
  nor (_00270_, _00268_, _06560_);
  or (_00272_, _00270_, _00266_);
  or (_00273_, _00272_, _00249_);
  and (_12049_, _00273_, _05552_);
  and (_00275_, _00248_, _11234_);
  and (_00276_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_00277_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_00278_, _00277_, _00276_);
  nor (_00279_, _00278_, _00265_);
  and (_00280_, _00267_, _11238_);
  or (_00281_, _00280_, _00279_);
  or (_00282_, _00281_, _00275_);
  and (_12055_, _00282_, _05552_);
  nor (_00283_, _11802_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00284_, _00283_, _11803_);
  and (_00285_, _00284_, _11792_);
  and (_00286_, _11811_, _07483_);
  not (_00287_, _11784_);
  nor (_00288_, _00287_, _07515_);
  and (_00289_, _11780_, _11275_);
  and (_00290_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_00292_, _00290_, _00289_);
  or (_00293_, _00292_, _00288_);
  or (_00294_, _00293_, _00286_);
  nor (_00295_, _00294_, _00285_);
  nand (_00296_, _00295_, _11774_);
  and (_00297_, _12025_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_00298_, _00297_, _12155_);
  or (_00299_, _12034_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00300_, _00299_, _12035_);
  or (_00301_, _00300_, _11828_);
  and (_00302_, _00301_, _12054_);
  and (_00303_, _00302_, _00298_);
  or (_00304_, _00303_, _00296_);
  nor (_00305_, _12066_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00306_, _00305_, _12068_);
  or (_00307_, _00306_, _11774_);
  and (_00308_, _00307_, _05552_);
  and (_12058_, _00308_, _00304_);
  nor (_00309_, _12017_, _11854_);
  nor (_00310_, _00309_, _12018_);
  and (_00311_, _00310_, _12054_);
  or (_00312_, _11817_, _11784_);
  and (_00313_, _00312_, _07574_);
  nor (_00314_, _11102_, _09047_);
  not (_00315_, _11848_);
  and (_00316_, _00315_, _11780_);
  and (_00317_, _11792_, _11391_);
  or (_00318_, _00317_, _00316_);
  or (_00319_, _00318_, _00314_);
  or (_00320_, _00319_, _00313_);
  or (_00321_, _00320_, _00311_);
  and (_00322_, _00321_, _11774_);
  nor (_00323_, _12060_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_00324_, _12060_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00325_, _00324_, _00323_);
  nor (_00326_, _00325_, _11774_);
  or (_00327_, _00326_, _00322_);
  and (_12065_, _00327_, _05552_);
  and (_00329_, _00254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_00330_, _00329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_00332_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_00333_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_00334_, _00333_, _00332_);
  nor (_00335_, _00246_, rst);
  and (_12067_, _00335_, _00334_);
  and (_00337_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_00338_, _05550_, _05786_);
  or (_00339_, _00338_, _00337_);
  and (_12070_, _00339_, _05552_);
  nor (_00340_, _09150_, _09094_);
  nor (_00341_, _00340_, _09151_);
  or (_00343_, _00341_, _09039_);
  or (_00344_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00345_, _00344_, _07933_);
  and (_00346_, _00345_, _00343_);
  and (_00347_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00348_, _00347_, _05552_);
  or (_12078_, _00348_, _00346_);
  and (_00349_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_00350_, _05550_, _11739_);
  or (_00351_, _00350_, _00349_);
  and (_12079_, _00351_, _05552_);
  nor (_12084_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  nor (_00352_, _09137_, _09116_);
  nor (_00353_, _00352_, _09139_);
  or (_00354_, _00353_, _09039_);
  or (_00355_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00356_, _00355_, _05605_);
  and (_00357_, _00356_, _00354_);
  and (_00358_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00359_, _00358_, _00357_);
  and (_12087_, _00359_, _05552_);
  and (_00360_, _09123_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00361_, _07919_, _05622_);
  nand (_00362_, _07919_, _05622_);
  and (_00363_, _00362_, _00361_);
  nand (_00364_, _00363_, _00360_);
  or (_00365_, _00363_, _00360_);
  and (_00366_, _00365_, _00364_);
  or (_00367_, _00366_, _05548_);
  or (_00368_, _05547_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00369_, _00368_, _07933_);
  and (_12102_, _00369_, _00367_);
  and (_00370_, _05916_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_00371_, _00370_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_12105_, _00371_, _05552_);
  nor (_12110_, _11943_, rst);
  not (_00372_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_00373_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_00374_, _00373_, _00372_);
  and (_00375_, _00374_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor (_00376_, _00373_, _00372_);
  or (_00377_, _00376_, _00374_);
  nand (_00378_, _00377_, _05552_);
  nor (_12113_, _00378_, _00375_);
  or (_00379_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_00380_, _00373_, rst);
  and (_12115_, _00380_, _00379_);
  and (_00381_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _07768_);
  and (_00382_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00383_, _00382_, _00381_);
  and (_12135_, _00383_, _05552_);
  nor (_00384_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_00385_, _00384_, _05573_);
  and (_00386_, _00385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_00387_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_00388_, _00385_, _00387_);
  or (_00389_, _00388_, _00386_);
  or (_00390_, _00389_, _00225_);
  or (_00391_, _08013_, _00387_);
  nand (_00392_, _00391_, _00225_);
  or (_00393_, _00392_, _08015_);
  and (_00394_, _00393_, _00390_);
  or (_00396_, _00394_, _00232_);
  nand (_00397_, _00232_, _08041_);
  and (_00398_, _00397_, _05552_);
  and (_12151_, _00398_, _00396_);
  nand (_00399_, _00241_, _06560_);
  or (_00400_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_00401_, _00400_, _05552_);
  and (_12158_, _00401_, _00399_);
  and (_00402_, _00248_, _06307_);
  and (_00403_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_00404_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_00405_, _00404_, _00403_);
  nor (_00406_, _00405_, _00265_);
  nor (_00407_, _00268_, _07388_);
  or (_00408_, _00407_, _00406_);
  or (_00409_, _00408_, _00402_);
  and (_12191_, _00409_, _05552_);
  nor (_00410_, _12059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00411_, _00410_, _12060_);
  or (_00412_, _00411_, _11774_);
  and (_00413_, _00412_, _05552_);
  and (_00414_, _00312_, _07635_);
  nor (_00415_, _11102_, _09106_);
  not (_00416_, _11872_);
  and (_00417_, _00416_, _11780_);
  and (_00418_, _11792_, _11449_);
  or (_00419_, _00418_, _00417_);
  or (_00420_, _00419_, _00415_);
  or (_00421_, _00420_, _00414_);
  or (_00422_, _11876_, _11877_);
  and (_00423_, _00422_, _12015_);
  nor (_00424_, _00422_, _12015_);
  or (_00425_, _00424_, _00423_);
  nand (_00426_, _00425_, _12054_);
  nand (_00427_, _00426_, _11774_);
  or (_00428_, _00427_, _00421_);
  and (_12275_, _00428_, _00413_);
  nand (_00429_, _08386_, _06949_);
  or (_00430_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_00431_, _00430_, _05552_);
  and (_12281_, _00431_, _00429_);
  and (_00432_, _00312_, _12189_);
  and (_00433_, _11792_, _11470_);
  not (_00434_, _11900_);
  and (_00435_, _00434_, _11780_);
  or (_00436_, _00435_, _00433_);
  or (_00437_, _12013_, _12010_);
  and (_00438_, _12054_, _12014_);
  and (_00439_, _00438_, _00437_);
  or (_00440_, _00439_, _00436_);
  or (_00441_, _00440_, _00432_);
  or (_00442_, _11102_, _09107_);
  nand (_00443_, _00442_, _11774_);
  or (_00444_, _00443_, _00441_);
  nor (_00445_, _08238_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00446_, _00445_, _12059_);
  or (_00447_, _00446_, _11774_);
  and (_00448_, _00447_, _05552_);
  and (_12286_, _00448_, _00444_);
  and (_00449_, _00225_, _10632_);
  nand (_00450_, _00449_, _06763_);
  not (_00451_, _00232_);
  or (_00452_, _00449_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_00453_, _00452_, _00451_);
  and (_00454_, _00453_, _00450_);
  nor (_00455_, _00451_, _06560_);
  or (_00456_, _00455_, _00454_);
  and (_12294_, _00456_, _05552_);
  nand (_00457_, _00241_, _07388_);
  or (_00458_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_00459_, _00458_, _05552_);
  and (_12323_, _00459_, _00457_);
  and (_00460_, _00248_, _11367_);
  and (_00461_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_00462_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_00463_, _00462_, _00461_);
  nor (_00464_, _00463_, _00265_);
  nor (_00465_, _00268_, _06306_);
  or (_00466_, _00465_, _00464_);
  or (_00467_, _00466_, _00460_);
  and (_12326_, _00467_, _05552_);
  or (_00468_, _11774_, _08240_);
  and (_00469_, _00468_, _05552_);
  and (_00470_, _00312_, _07483_);
  nor (_00471_, _11102_, _09048_);
  not (_00472_, _11921_);
  and (_00473_, _00472_, _11780_);
  and (_00474_, _11792_, _11275_);
  or (_00476_, _00474_, _00473_);
  or (_00477_, _00476_, _00471_);
  or (_00478_, _00477_, _00470_);
  or (_00479_, _11925_, _11926_);
  nor (_00480_, _00479_, _12008_);
  and (_00481_, _00479_, _12008_);
  or (_00482_, _00481_, _00480_);
  nand (_00483_, _00482_, _12054_);
  nand (_00484_, _00483_, _11774_);
  or (_00485_, _00484_, _00478_);
  and (_12343_, _00485_, _00469_);
  or (_00486_, _11774_, _08253_);
  and (_00487_, _00486_, _05552_);
  and (_00488_, _00312_, _08144_);
  nor (_00489_, _11102_, _08236_);
  and (_00490_, _11944_, _11780_);
  and (_00491_, _11792_, _11747_);
  or (_00492_, _00491_, _00490_);
  or (_00493_, _00492_, _00489_);
  or (_00494_, _00493_, _00488_);
  nor (_00495_, _12006_, _12004_);
  nor (_00496_, _00495_, _12007_);
  nand (_00497_, _00496_, _12054_);
  nand (_00498_, _00497_, _11774_);
  or (_00499_, _00498_, _00494_);
  and (_12346_, _00499_, _00487_);
  and (_00500_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_00501_, _00500_, _08062_);
  and (_00502_, _00501_, _00225_);
  not (_00503_, _00225_);
  or (_00504_, _00503_, _08059_);
  and (_00505_, _00504_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_00506_, _00505_, _00232_);
  or (_00507_, _00506_, _00502_);
  nand (_00508_, _00232_, _07388_);
  and (_00509_, _00508_, _05552_);
  and (_12356_, _00509_, _00507_);
  and (_00510_, _00248_, _07439_);
  not (_00511_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor (_00512_, _00259_, _00511_);
  and (_00513_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_00515_, _00513_, _00512_);
  nor (_00516_, _00515_, _00265_);
  nor (_00517_, _00268_, _08386_);
  or (_00518_, _00517_, _00516_);
  or (_00519_, _00518_, _00510_);
  and (_12358_, _00519_, _05552_);
  and (_00520_, _00312_, _08102_);
  and (_00521_, _11811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00522_, _11968_, _11780_);
  and (_00523_, _11792_, _11617_);
  or (_00524_, _00523_, _00522_);
  or (_00525_, _00524_, _00521_);
  nor (_00526_, _12000_, _11998_);
  nor (_00527_, _00526_, _12001_);
  and (_00528_, _00527_, _12054_);
  or (_00529_, _00528_, _00525_);
  nor (_00531_, _00529_, _00520_);
  nand (_00532_, _00531_, _11774_);
  or (_00534_, _11774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00535_, _00534_, _05552_);
  and (_12361_, _00535_, _00532_);
  and (_00536_, _00312_, _07711_);
  or (_00537_, _11997_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_00538_, _11998_);
  and (_00539_, _12161_, _00538_);
  and (_00540_, _00539_, _00537_);
  and (_00541_, _11994_, _11780_);
  and (_00542_, _11792_, _11691_);
  and (_00543_, _11811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00544_, _00543_, _00542_);
  or (_00545_, _00544_, _00541_);
  or (_00546_, _00545_, _00540_);
  nor (_00547_, _00546_, _00536_);
  nand (_00548_, _00547_, _11774_);
  or (_00550_, _11774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00551_, _00550_, _05552_);
  and (_12370_, _00551_, _00548_);
  and (_00552_, _00225_, _08635_);
  nand (_00553_, _00552_, _06763_);
  or (_00554_, _00552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_00555_, _00554_, _00451_);
  and (_00556_, _00555_, _00553_);
  nor (_00557_, _00451_, _06306_);
  or (_00558_, _00557_, _00556_);
  and (_12383_, _00558_, _05552_);
  and (_00559_, _00312_, _07255_);
  and (_00560_, _11792_, _11328_);
  not (_00561_, _07758_);
  and (_00562_, _11780_, _00561_);
  or (_00563_, _00562_, _00560_);
  or (_00564_, _11830_, _11829_);
  not (_00565_, _00564_);
  nand (_00566_, _00565_, _12019_);
  or (_00567_, _00565_, _12019_);
  and (_00568_, _00567_, _12054_);
  and (_00569_, _00568_, _00566_);
  or (_00570_, _00569_, _00563_);
  or (_00571_, _00570_, _00559_);
  or (_00572_, _11102_, _09046_);
  nand (_00573_, _00572_, _11774_);
  or (_00574_, _00573_, _00571_);
  nor (_00575_, _00324_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00576_, _12061_, _12060_);
  nor (_00577_, _00576_, _00575_);
  or (_00578_, _00577_, _11774_);
  and (_00579_, _00578_, _05552_);
  and (_12440_, _00579_, _00574_);
  and (_00580_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_00581_, _00580_, _08998_);
  and (_00582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08998_);
  and (_00583_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00584_, _00583_, _00582_);
  and (_00585_, _00584_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_00586_, _00585_, _08996_);
  not (_00587_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_00588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_00589_, _00588_, _00587_);
  and (_00590_, _00589_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_00591_, _00590_);
  not (_00592_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_00593_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_00594_, _00593_, _00592_);
  nand (_00595_, _00594_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_00596_, _00595_, _00591_);
  and (_00597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_00598_, _00597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  not (_00599_, _00598_);
  and (_00600_, _00599_, _00596_);
  and (_00601_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_00602_, _00601_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  not (_00603_, _00602_);
  and (_00605_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00607_, _00605_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_00608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_00609_, _00608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_00610_, _00609_, _00607_);
  and (_00611_, _00610_, _00603_);
  and (_00612_, _00611_, _00600_);
  nor (_00613_, _00612_, _00586_);
  and (_00614_, _08996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not (_00615_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_00616_, _00589_, _00615_);
  not (_00617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_00618_, _00594_, _00617_);
  nor (_00619_, _00618_, _00616_);
  not (_00620_, _00619_);
  and (_00621_, _00620_, _00614_);
  not (_00622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_00623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_00624_, _00623_, _00622_);
  and (_00625_, _00624_, _00614_);
  or (_00626_, _00625_, _00621_);
  or (_00627_, _00626_, _00613_);
  nand (_00628_, _00613_, _00600_);
  and (_00629_, _00628_, _00627_);
  and (_00630_, _00629_, _00581_);
  or (_00631_, _00630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_00632_, _00581_);
  not (_00633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_00634_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_00635_, _00634_, _00633_);
  not (_00636_, _00635_);
  not (_00637_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_00639_, _00638_, _00637_);
  not (_00640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_00641_, _00608_, _00640_);
  nor (_00642_, _00641_, _00639_);
  and (_00643_, _00642_, _00636_);
  not (_00644_, _00624_);
  and (_00645_, _00643_, _00644_);
  nand (_00646_, _00645_, _00619_);
  nand (_00647_, _00646_, _00614_);
  nor (_00648_, _00647_, _00613_);
  not (_00649_, _00648_);
  or (_00650_, _00649_, _00643_);
  or (_00651_, _00611_, _00586_);
  and (_00652_, _00651_, _00650_);
  or (_00653_, _00652_, _00632_);
  and (_00654_, _00653_, _05552_);
  and (_12455_, _00654_, _00631_);
  and (_00655_, _12024_, _11828_);
  and (_00656_, _12021_, _11796_);
  nor (_00657_, _00656_, _11828_);
  or (_00658_, _00657_, _00655_);
  nand (_00659_, _00658_, _06219_);
  or (_00660_, _00658_, _06219_);
  and (_00661_, _00660_, _12161_);
  and (_00662_, _00661_, _00659_);
  and (_00663_, _11811_, _08144_);
  nor (_00664_, _00287_, _08200_);
  and (_00665_, _11780_, _11747_);
  and (_00666_, _11792_, _05781_);
  and (_00667_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_00668_, _00667_, _00666_);
  or (_00669_, _00668_, _00665_);
  nor (_00670_, _00669_, _00664_);
  nand (_00671_, _00670_, _11774_);
  or (_00672_, _00671_, _00663_);
  or (_00673_, _00672_, _00662_);
  and (_00674_, _00324_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00675_, _00674_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00676_, _00675_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nand (_00677_, _00676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_00678_, _00676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00679_, _00678_, _00677_);
  or (_00680_, _00679_, _11774_);
  and (_00681_, _00680_, _05552_);
  and (_12467_, _00681_, _00673_);
  and (_00683_, _12021_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_00685_, _00683_, _11828_);
  nand (_00686_, _12022_, _11828_);
  and (_00687_, _00686_, _00685_);
  and (_00688_, _00687_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_00689_, _00687_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_00690_, _00689_, _12161_);
  nor (_00691_, _00690_, _00688_);
  and (_00692_, _11811_, _08102_);
  nor (_00693_, _00287_, _08173_);
  and (_00694_, _11792_, _05803_);
  and (_00695_, _11780_, _11617_);
  and (_00696_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_00697_, _00696_, _00695_);
  or (_00698_, _00697_, _00694_);
  nor (_00699_, _00698_, _00693_);
  nand (_00700_, _00699_, _11774_);
  or (_00701_, _00700_, _00692_);
  or (_00702_, _00701_, _00691_);
  nor (_00703_, _00675_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00704_, _00703_, _00676_);
  or (_00705_, _00704_, _11774_);
  and (_00706_, _00705_, _05552_);
  and (_12520_, _00706_, _00702_);
  and (_00707_, _11811_, _07711_);
  and (_00708_, _11784_, _08228_);
  and (_00709_, _11792_, _07781_);
  and (_00710_, _11780_, _11691_);
  or (_00711_, _00710_, _00709_);
  and (_00712_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00713_, _00712_, _00711_);
  or (_00714_, _00713_, _00708_);
  or (_00715_, _00686_, _00683_);
  and (_00716_, _12021_, _06192_);
  nor (_00717_, _12021_, _06192_);
  or (_00718_, _00717_, _00716_);
  or (_00719_, _00718_, _11828_);
  and (_00720_, _00719_, _00715_);
  and (_00721_, _00720_, _12054_);
  or (_00722_, _00721_, _00714_);
  or (_00723_, _00722_, _00707_);
  or (_00724_, _00723_, _13414_);
  nor (_00725_, _00576_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00726_, _00725_, _00675_);
  or (_00727_, _00726_, _11774_);
  and (_00728_, _00727_, _05552_);
  and (_12523_, _00728_, _00724_);
  nor (_12598_, _11193_, rst);
  nor (_00729_, _08041_, _07939_);
  and (_00730_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or (_00731_, _00730_, _00729_);
  and (_12772_, _00731_, _05552_);
  and (_12807_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and (pc_log_change, _05608_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_00732_, _10861_, _08013_);
  or (_00733_, _00732_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_00734_, _00733_, _08992_);
  nand (_00735_, _00732_, _06763_);
  and (_00736_, _00735_, _00734_);
  nor (_00737_, _08992_, _08041_);
  or (_00738_, _00737_, _00736_);
  and (_13106_, _00738_, _05552_);
  and (_00739_, _10861_, _06060_);
  or (_00740_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_00741_, _00740_, _08992_);
  nand (_00742_, _00739_, _06763_);
  and (_00743_, _00742_, _00741_);
  and (_00744_, _08991_, _11238_);
  or (_00745_, _00744_, _00743_);
  and (_13109_, _00745_, _05552_);
  and (_00746_, _10633_, _07443_);
  nand (_00747_, _00746_, _06306_);
  and (_00748_, _13775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_00749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00749_);
  nor (_00751_, _00750_, _00748_);
  and (_00752_, _08989_, _08635_);
  and (_00753_, _00752_, _07443_);
  nor (_00754_, _00753_, _00751_);
  not (_00755_, _00754_);
  and (_00756_, _00755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not (_00757_, _00751_);
  not (_00758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_00759_, _00758_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not (_00760_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00761_, \oc8051_top_1.oc8051_sfr1.pres_ow , _00760_);
  not (_00762_, t1_i);
  and (_00763_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00764_, _00763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or (_00765_, _00764_, _00761_);
  and (_00766_, _00765_, _00759_);
  and (_00767_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00768_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_00769_, _00768_, _00767_);
  and (_00770_, _00769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00772_, _00770_, _00766_);
  nor (_00773_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00774_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_00775_, _00774_, _00773_);
  and (_00776_, _00775_, _00757_);
  and (_00777_, _00774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00779_, _00778_, _00748_);
  and (_00780_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_00781_, _00780_, _00776_);
  nor (_00782_, _00781_, _00753_);
  or (_00783_, _00782_, _00756_);
  or (_00784_, _00783_, _00746_);
  and (_00785_, _00784_, _05552_);
  and (_13129_, _00785_, _00747_);
  nand (_00786_, _00746_, _07388_);
  and (_00787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_00788_, _00787_, _00753_);
  not (_00789_, _00788_);
  and (_00790_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00791_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not (_00792_, _00787_);
  and (_00794_, _00769_, _00766_);
  and (_00795_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_00796_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_00797_, _00796_, _00795_);
  and (_00798_, _00797_, _00792_);
  nor (_00799_, _00798_, _00791_);
  nor (_00800_, _00799_, _00753_);
  or (_00801_, _00800_, _00790_);
  or (_00802_, _00801_, _00746_);
  and (_00803_, _00802_, _05552_);
  and (_13132_, _00803_, _00786_);
  nand (_00804_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_00805_, _00804_, _00753_);
  and (_00806_, _00766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00808_, _00806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00809_, _00808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_00810_, _00809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_00811_, _00810_, _00794_);
  and (_00812_, _00811_, _00788_);
  and (_00813_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_00814_, _00813_, _00812_);
  or (_00816_, _00814_, _00805_);
  or (_00817_, _00816_, _00746_);
  nand (_00818_, _00746_, _06560_);
  and (_00819_, _00818_, _05552_);
  and (_13135_, _00819_, _00817_);
  nand (_00820_, _00746_, _08386_);
  nand (_00821_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00822_, _00821_, _00753_);
  and (_00823_, _00755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00825_, _00824_, _00795_);
  nor (_00826_, _00774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00827_, _00826_, _00825_);
  and (_00828_, _00827_, _00754_);
  or (_00829_, _00828_, _00823_);
  or (_00830_, _00829_, _00822_);
  or (_00831_, _00830_, _00746_);
  and (_00832_, _00831_, _05552_);
  and (_13139_, _00832_, _00820_);
  nor (_00833_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_00834_, _00833_, _00648_);
  and (_00835_, _00833_, _00613_);
  or (_00836_, _00835_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_00837_, _00836_, _05552_);
  and (_13142_, _00837_, _00834_);
  not (_00838_, _00580_);
  or (_00839_, _00838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00840_, _00839_, _05552_);
  not (_00841_, _00610_);
  or (_00842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_00843_, _00842_, _00841_);
  nor (_00844_, _00595_, _08998_);
  nor (_00845_, _00844_, _00598_);
  and (_00846_, _00590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00847_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00848_, _00847_, _00610_);
  and (_00849_, _00848_, _00845_);
  or (_00850_, _00849_, _00843_);
  and (_00851_, _00850_, _00603_);
  and (_00852_, _00610_, _00598_);
  or (_00853_, _00852_, _00602_);
  and (_00854_, _00853_, _09009_);
  or (_00855_, _00854_, _00851_);
  and (_00856_, _00855_, _00613_);
  not (_00857_, _00613_);
  and (_00858_, _00842_, _00636_);
  or (_00859_, _00858_, _00643_);
  and (_00860_, _00624_, _09009_);
  not (_00861_, _00642_);
  and (_00862_, _00618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00863_, _00862_, _00624_);
  and (_00864_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00865_, _00864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00866_, _00865_, _00863_);
  or (_00867_, _00866_, _00861_);
  or (_00868_, _00867_, _00860_);
  and (_00869_, _00868_, _00859_);
  and (_00870_, _00635_, _09009_);
  or (_00871_, _00870_, _00647_);
  or (_00872_, _00871_, _00869_);
  not (_00873_, _00647_);
  or (_00874_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00875_, _00874_, _00872_);
  and (_00876_, _00875_, _00857_);
  or (_00877_, _00876_, _00856_);
  or (_00878_, _00877_, _00580_);
  and (_13150_, _00878_, _00840_);
  and (_00879_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00881_, _00824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00882_, _00881_, _00880_);
  and (_00883_, _00882_, _00769_);
  and (_00884_, _00883_, _00748_);
  nor (_00885_, _00766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_00886_, _00885_, _00806_);
  and (_00887_, _00886_, _00792_);
  nor (_00888_, _00887_, _00884_);
  nor (_00889_, _00888_, _00753_);
  or (_00890_, _00889_, _00746_);
  or (_00891_, _00890_, _00879_);
  nand (_00892_, _00746_, _07945_);
  and (_00893_, _00892_, _05552_);
  and (_13154_, _00893_, _00891_);
  nor (_00895_, _08386_, _07939_);
  and (_00896_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_00897_, _00896_, _00895_);
  and (_13157_, _00897_, _05552_);
  nand (_00898_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00899_, _00898_, _00753_);
  nor (_00900_, _00806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_00901_, _00900_, _00808_);
  and (_00902_, _00901_, _00788_);
  or (_00903_, _00902_, _00899_);
  and (_00904_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_00905_, _00904_, _00746_);
  or (_00906_, _00905_, _00903_);
  nand (_00907_, _00746_, _07975_);
  and (_00908_, _00907_, _05552_);
  and (_13163_, _00908_, _00906_);
  nor (_00909_, _00808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_00911_, _00909_, _00809_);
  nand (_00912_, _00911_, _00788_);
  or (_00913_, _00788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00914_, _00913_, _00912_);
  nand (_00915_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_00916_, _00915_, _00753_);
  or (_00918_, _00916_, _00746_);
  or (_00919_, _00918_, _00914_);
  nand (_00920_, _00746_, _08041_);
  and (_00921_, _00920_, _05552_);
  and (_13167_, _00921_, _00919_);
  nand (_00923_, _00648_, _00581_);
  and (_00924_, _00613_, _00581_);
  or (_00926_, _00924_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_00927_, _00926_, _05552_);
  and (_13175_, _00927_, _00923_);
  not (_00929_, _00746_);
  and (_00931_, _00883_, _00766_);
  or (_00932_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_00934_, _00750_);
  and (_00935_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00936_, _00935_, _00934_);
  and (_00937_, _00936_, _00932_);
  nor (_00939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_00940_, _00939_);
  and (_00942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00943_, _00942_, _00772_);
  nor (_00944_, _00943_, _00940_);
  or (_00945_, _00944_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00946_, _00880_, _00794_);
  and (_00947_, _00944_, _00946_);
  or (_00948_, _00947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00949_, _00948_, _00945_);
  nor (_00950_, _00949_, _00937_);
  nor (_00951_, _00950_, _00753_);
  not (_00952_, _00753_);
  nor (_00953_, _00952_, _07975_);
  or (_00954_, _00953_, _00951_);
  and (_00955_, _00954_, _00929_);
  and (_00956_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00957_, _00956_, _00955_);
  and (_13191_, _00957_, _05552_);
  nand (_00958_, _00753_, _08041_);
  nand (_00959_, _00943_, _00939_);
  nor (_00960_, _00959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00963_, _00961_, _00931_);
  or (_00964_, _00935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_00965_, _00964_, _00750_);
  nor (_00967_, _00965_, _00963_);
  and (_00968_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_00969_, _00968_, _00967_);
  or (_00971_, _00969_, _00960_);
  or (_00972_, _00971_, _00753_);
  and (_00973_, _00972_, _00929_);
  and (_00974_, _00973_, _00958_);
  and (_00975_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_00976_, _00975_, _00974_);
  and (_13194_, _00976_, _05552_);
  and (_00977_, _00753_, _11238_);
  not (_00978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00979_, _00939_, _00795_);
  and (_00980_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00981_, _00980_, _00750_);
  nor (_00982_, _00981_, _00979_);
  nand (_00983_, _00982_, _00978_);
  or (_00984_, _00982_, _00978_);
  nand (_00985_, _00984_, _00983_);
  nor (_00986_, _00985_, _00753_);
  or (_00987_, _00986_, _00746_);
  or (_00988_, _00987_, _00977_);
  nand (_00989_, _00746_, _00978_);
  and (_00991_, _00989_, _05552_);
  and (_13197_, _00991_, _00988_);
  nand (_00993_, _00753_, _07388_);
  or (_00994_, _00963_, _00934_);
  and (_00995_, _00961_, _00749_);
  and (_00997_, _00995_, _00946_);
  or (_00998_, _00997_, _00750_);
  and (_01000_, _00998_, _00994_);
  nand (_01001_, _01000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_01002_, _01001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_01003_, _01001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_01004_, _01003_, _01002_);
  or (_01005_, _01004_, _00753_);
  and (_01006_, _01005_, _00929_);
  and (_01007_, _01006_, _00993_);
  and (_01008_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_01009_, _01008_, _01007_);
  and (_13203_, _01009_, _05552_);
  nand (_01010_, _00753_, _08386_);
  and (_01011_, _00961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_01012_, _01011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_01013_, _01012_, _00931_);
  nor (_01014_, _01013_, _00934_);
  and (_01015_, _01012_, _00749_);
  and (_01016_, _01015_, _00946_);
  nor (_01017_, _01016_, _00750_);
  nor (_01018_, _01017_, _01014_);
  nand (_01019_, _01018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_01020_, _01019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_01021_, _01019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_01022_, _01021_, _01020_);
  or (_01023_, _01022_, _00753_);
  and (_01024_, _01023_, _00929_);
  and (_01025_, _01024_, _01010_);
  and (_01026_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_01027_, _01026_, _01025_);
  and (_13206_, _01027_, _05552_);
  nand (_01029_, _00753_, _06306_);
  or (_01030_, _01018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_01031_, _01030_, _01019_);
  or (_01032_, _01031_, _00753_);
  and (_01033_, _01032_, _00929_);
  and (_01035_, _01033_, _01029_);
  and (_01036_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_01038_, _01036_, _01035_);
  and (_13209_, _01038_, _05552_);
  nand (_01039_, _00753_, _06560_);
  or (_01040_, _01000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_01041_, _01040_, _01001_);
  or (_01043_, _01041_, _00753_);
  and (_01045_, _01043_, _00929_);
  and (_01047_, _01045_, _01039_);
  and (_01048_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_01049_, _01048_, _01047_);
  and (_13212_, _01049_, _05552_);
  not (_01050_, t0_i);
  and (_01051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01050_);
  nor (_01052_, _01051_, _00073_);
  not (_01053_, _01052_);
  not (_01054_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_01055_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_01056_, _01055_, _01054_);
  and (_01058_, _01056_, _01053_);
  and (_01059_, _01058_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_01060_, _01059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_01061_, _01059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_01063_, _01061_, _01060_);
  not (_01064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_01066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_01067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_01068_, _01067_, _01066_);
  and (_01069_, _01068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_01070_, _01069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_01071_, _01070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_01072_, _01071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13526_);
  and (_01075_, _01074_, _01058_);
  nand (_01076_, _01075_, _01072_);
  or (_01078_, _01076_, _01064_);
  and (_01079_, _01078_, _01063_);
  and (_01081_, _08989_, _08057_);
  and (_01082_, _01081_, _07443_);
  nor (_01084_, _01082_, _01079_);
  and (_01085_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_01087_, _01085_, _01084_);
  and (_01089_, _10627_, _07443_);
  not (_01091_, _01089_);
  and (_01093_, _01091_, _01087_);
  nor (_01095_, _01091_, _07975_);
  or (_01096_, _01095_, _01093_);
  and (_13215_, _01096_, _05552_);
  not (_01098_, _01058_);
  nor (_01100_, _01082_, _01098_);
  or (_01101_, _01100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_01102_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_01104_, _01102_, _01072_);
  nand (_01105_, _01104_, _01059_);
  or (_01106_, _01105_, _01082_);
  and (_01107_, _01106_, _01101_);
  or (_01108_, _01107_, _01089_);
  nand (_01109_, _01089_, _07945_);
  and (_01110_, _01109_, _05552_);
  and (_13219_, _01110_, _01108_);
  not (_01111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand (_01112_, _01082_, _01111_);
  and (_01113_, _01061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_01114_, _01061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_01115_, _01114_, _01113_);
  and (_01116_, _01071_, _01058_);
  and (_01117_, _01116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01118_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01119_, _01118_, _01117_);
  or (_01120_, _01119_, _01115_);
  or (_01121_, _01120_, _01082_);
  and (_01122_, _01121_, _01112_);
  or (_01123_, _01122_, _01089_);
  nand (_01124_, _01089_, _08041_);
  and (_01126_, _01124_, _05552_);
  and (_13237_, _01126_, _01123_);
  and (_01127_, _01068_, _01058_);
  nor (_01128_, _01127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_01129_, _01127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_01131_, _01129_, _01128_);
  and (_01132_, _01072_, _01058_);
  and (_01133_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01134_, _01133_, _01132_);
  nor (_01136_, _01134_, _01131_);
  nor (_01137_, _01136_, _01082_);
  and (_01138_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_01139_, _01138_, _01137_);
  and (_01140_, _01139_, _01091_);
  nor (_01141_, _01091_, _07388_);
  or (_01142_, _01141_, _01140_);
  and (_13242_, _01142_, _05552_);
  nor (_01144_, _01113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_01145_, _01144_, _01127_);
  and (_01146_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01147_, _01146_, _01117_);
  or (_01148_, _01147_, _01145_);
  or (_01149_, _01148_, _01082_);
  not (_01151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand (_01152_, _01082_, _01151_);
  and (_01153_, _01152_, _01091_);
  and (_01154_, _01153_, _01149_);
  nor (_01155_, _01091_, _06560_);
  or (_01156_, _01155_, _01154_);
  and (_13245_, _01156_, _05552_);
  or (_01157_, _00838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01158_, _01157_, _05552_);
  and (_01159_, _00853_, _09008_);
  or (_01160_, _08998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_01161_, _01160_, _00610_);
  and (_01162_, _01161_, _00603_);
  and (_01163_, _00590_, _08998_);
  or (_01164_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nor (_01165_, _00595_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01166_, _01165_, _00598_);
  and (_01167_, _01166_, _01164_);
  or (_01168_, _01167_, _00841_);
  and (_01170_, _01168_, _01162_);
  or (_01171_, _01170_, _01159_);
  and (_01172_, _01171_, _00613_);
  and (_01173_, _01160_, _00636_);
  or (_01174_, _01173_, _00643_);
  and (_01175_, _00624_, _09008_);
  and (_01176_, _00618_, _08998_);
  nor (_01177_, _01176_, _00624_);
  and (_01178_, _00616_, _08998_);
  or (_01179_, _01178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01180_, _01179_, _01177_);
  or (_01181_, _01180_, _00861_);
  or (_01183_, _01181_, _01175_);
  and (_01184_, _01183_, _01174_);
  and (_01185_, _00635_, _09008_);
  or (_01186_, _01185_, _00647_);
  or (_01187_, _01186_, _01184_);
  or (_01188_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01189_, _01188_, _01187_);
  and (_01190_, _01189_, _00857_);
  or (_01191_, _01190_, _01172_);
  or (_01192_, _01191_, _00580_);
  and (_13250_, _01192_, _01158_);
  or (_01194_, _08998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_01195_, _01194_, _00603_);
  not (_01196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_01197_, _01163_, _01196_);
  nand (_01198_, _01197_, _01166_);
  or (_01199_, _00599_, _08997_);
  and (_01200_, _01199_, _01198_);
  or (_01202_, _01200_, _00609_);
  not (_01203_, _00607_);
  not (_01204_, _00609_);
  or (_01205_, _01194_, _01204_);
  and (_01206_, _01205_, _01203_);
  and (_01208_, _01206_, _01202_);
  and (_01209_, _00607_, _08997_);
  or (_01210_, _01209_, _00602_);
  or (_01212_, _01210_, _01208_);
  and (_01213_, _01212_, _01195_);
  or (_01214_, _01213_, _00857_);
  or (_01215_, _01194_, _00636_);
  or (_01217_, _01178_, _01196_);
  nand (_01218_, _01217_, _01177_);
  or (_01219_, _00644_, _08997_);
  and (_01220_, _01219_, _01218_);
  or (_01221_, _01220_, _00641_);
  not (_01222_, _00639_);
  not (_01223_, _00641_);
  or (_01224_, _01194_, _01223_);
  and (_01225_, _01224_, _01222_);
  and (_01226_, _01225_, _01221_);
  and (_01227_, _00639_, _08997_);
  or (_01228_, _01227_, _00635_);
  or (_01229_, _01228_, _01226_);
  and (_01230_, _01229_, _01215_);
  or (_01231_, _01230_, _00649_);
  and (_01232_, _01231_, _01214_);
  or (_01233_, _01232_, _00580_);
  nor (_01234_, _00873_, _00613_);
  nor (_01235_, _01234_, _00580_);
  or (_01236_, _01235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_01237_, _01236_, _05552_);
  and (_13262_, _01237_, _01233_);
  and (_01238_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_13271_, _01238_, _00580_);
  or (_01239_, _00641_, _00624_);
  and (_01240_, _00619_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01241_, _01240_, _01239_);
  and (_01242_, _01241_, _01222_);
  and (_01243_, _00648_, _00636_);
  and (_01244_, _01243_, _01242_);
  or (_01245_, _00609_, _00598_);
  and (_01246_, _00596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01247_, _01246_, _01245_);
  and (_01248_, _01247_, _01203_);
  and (_01249_, _00613_, _00603_);
  and (_01250_, _01249_, _01248_);
  or (_01251_, _01250_, _00580_);
  or (_01252_, _01251_, _01244_);
  nand (_01253_, _00580_, _05910_);
  and (_01254_, _01253_, _05552_);
  and (_13276_, _01254_, _01252_);
  nor (_01255_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01256_, _01255_, _00618_);
  or (_01257_, _01256_, _00624_);
  and (_01258_, _01257_, _01223_);
  or (_01259_, _01258_, _00639_);
  and (_01260_, _01259_, _01243_);
  or (_01261_, _00590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01262_, _01261_, _00595_);
  or (_01263_, _01262_, _00598_);
  and (_01264_, _01263_, _01204_);
  or (_01266_, _01264_, _00607_);
  and (_01267_, _01266_, _01249_);
  or (_01268_, _01267_, _00580_);
  or (_01269_, _01268_, _01260_);
  or (_01270_, _00838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01271_, _01270_, _05552_);
  and (_13279_, _01271_, _01269_);
  and (_01272_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_01273_, _01272_, _01235_);
  and (_13282_, _01273_, _05552_);
  not (_01274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_01275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_01276_, _01275_);
  and (_01277_, _01276_, _01058_);
  nand (_01278_, _01277_, _01071_);
  nor (_01279_, _01278_, _01082_);
  nor (_01280_, _01279_, _01274_);
  not (_01281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_01282_, _01076_, _01281_);
  not (_01283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_01284_, _01275_, _01283_);
  and (_01285_, _01284_, _01129_);
  nand (_01286_, _01285_, _01278_);
  and (_01287_, _01286_, _01282_);
  nor (_01288_, _01287_, _01082_);
  or (_01289_, _01288_, _01280_);
  and (_01290_, _01289_, _01091_);
  nor (_01291_, _01091_, _08386_);
  or (_01292_, _01291_, _01290_);
  and (_13293_, _01292_, _05552_);
  and (_13296_, _00580_, _07727_);
  and (_01293_, _01129_, _01276_);
  and (_01294_, _01293_, _01283_);
  not (_01295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_01296_, _01076_, _01295_);
  nor (_01297_, _01296_, _01294_);
  nor (_01298_, _01297_, _01082_);
  not (_01299_, _01293_);
  or (_01300_, _01299_, _01082_);
  and (_01301_, _01300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_01302_, _01301_, _01298_);
  and (_01303_, _01302_, _01091_);
  nor (_01304_, _01091_, _06306_);
  or (_01305_, _01304_, _01303_);
  and (_13301_, _01305_, _05552_);
  nand (_01306_, _01082_, _08386_);
  and (_01307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01308_, _01307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_01310_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01311_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_01312_, _01311_, _01310_);
  and (_01313_, _01312_, _01308_);
  and (_01314_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_01315_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01316_, _01312_, _01307_);
  and (_01317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01318_, _01317_, _01316_);
  nand (_01319_, _01318_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01320_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01321_, _01320_, _01315_);
  and (_01322_, _01308_, _01310_);
  and (_01323_, _01322_, _01129_);
  nor (_01324_, _01323_, _01281_);
  and (_01325_, _01323_, _01281_);
  or (_01326_, _01325_, _01324_);
  and (_01327_, _01326_, _01275_);
  and (_01328_, _01310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01329_, _01328_, _01117_);
  nand (_01330_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_01331_, _01330_, _01295_);
  nand (_01332_, _01331_, _01281_);
  and (_01333_, _00146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_01334_, _01331_, _01281_);
  and (_01335_, _01334_, _01333_);
  and (_01336_, _01335_, _01332_);
  or (_01337_, _01336_, _01327_);
  or (_01338_, _01337_, _01321_);
  or (_01339_, _01338_, _01082_);
  and (_01340_, _01339_, _01091_);
  and (_01341_, _01340_, _01306_);
  and (_01342_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_01343_, _01342_, _01341_);
  and (_13330_, _01343_, _05552_);
  nand (_01344_, _01082_, _08041_);
  and (_01345_, _01309_, _01129_);
  or (_01346_, _01345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01347_, _01345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_01348_, _01347_, _01276_);
  and (_01349_, _01348_, _01346_);
  and (_01350_, _01309_, _01132_);
  or (_01351_, _01350_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_01353_, _01310_, _01132_);
  and (_01354_, _01353_, _01333_);
  and (_01356_, _01354_, _01351_);
  and (_01357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01358_, _01311_, _01309_);
  or (_01359_, _01358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_01360_, _01359_, _01357_);
  nor (_01361_, _01360_, _01312_);
  or (_01362_, _01361_, _01118_);
  or (_01364_, _01362_, _01356_);
  or (_01365_, _01364_, _01349_);
  or (_01367_, _01365_, _01082_);
  and (_01368_, _01367_, _01091_);
  and (_01369_, _01368_, _01344_);
  and (_01370_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_01371_, _01370_, _01369_);
  and (_13338_, _01371_, _05552_);
  nand (_01372_, _01082_, _06560_);
  or (_01373_, _01347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01374_, _01347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_01375_, _01374_, _01276_);
  and (_01376_, _01375_, _01373_);
  or (_01377_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01378_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_01379_, _01378_);
  and (_01380_, _01379_, _01357_);
  and (_01381_, _01380_, _01377_);
  and (_01382_, _01132_, _00146_);
  and (_01383_, _01382_, _01310_);
  or (_01384_, _01383_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_01385_, _01333_, _01074_);
  nand (_01386_, _01383_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01388_, _01386_, _01385_);
  and (_01389_, _01388_, _01384_);
  or (_01390_, _01389_, _01381_);
  or (_01392_, _01390_, _01376_);
  or (_01393_, _01392_, _01082_);
  and (_01394_, _01393_, _01091_);
  and (_01396_, _01394_, _01372_);
  and (_01397_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_01398_, _01397_, _01396_);
  and (_13340_, _01398_, _05552_);
  nand (_01399_, _01082_, _07388_);
  or (_01400_, _01374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01401_, _01374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_01402_, _01401_, _01276_);
  and (_01404_, _01402_, _01400_);
  and (_01405_, _01328_, _01132_);
  or (_01406_, _01405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01407_, _01330_, _01333_);
  and (_01408_, _01407_, _01406_);
  or (_01409_, _01378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_01410_, _01409_, _01357_);
  nor (_01411_, _01410_, _01316_);
  or (_01412_, _01411_, _01133_);
  or (_01413_, _01412_, _01408_);
  or (_01414_, _01413_, _01404_);
  or (_01415_, _01414_, _01082_);
  and (_01416_, _01415_, _01091_);
  and (_01417_, _01416_, _01399_);
  and (_01418_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_01419_, _01418_, _01417_);
  and (_13348_, _01419_, _05552_);
  nand (_01420_, _01082_, _06306_);
  or (_01422_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_01423_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01424_, _01423_, _01275_);
  and (_01425_, _01424_, _01422_);
  or (_01426_, _01316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_01427_, _01313_);
  and (_01428_, _01427_, _01357_);
  and (_01429_, _01428_, _01426_);
  and (_01430_, _01405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01431_, _01430_, _00146_);
  nor (_01432_, _01431_, _01295_);
  and (_01433_, _01431_, _01295_);
  or (_01434_, _01433_, _01432_);
  and (_01435_, _01434_, _01385_);
  or (_01438_, _01435_, _01429_);
  or (_01439_, _01438_, _01425_);
  or (_01440_, _01439_, _01082_);
  and (_01441_, _01440_, _01091_);
  and (_01442_, _01441_, _01420_);
  and (_01443_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_01445_, _01443_, _01442_);
  and (_13351_, _01445_, _05552_);
  nand (_01446_, _01082_, _07975_);
  nand (_01448_, _01382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_01450_, _01448_, _01064_);
  not (_01451_, _01350_);
  and (_01452_, _01451_, _01333_);
  or (_01454_, _01452_, _01074_);
  and (_01455_, _01454_, _01450_);
  and (_01456_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_01457_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_01458_, _01358_);
  and (_01460_, _01458_, _01357_);
  and (_01461_, _01460_, _01457_);
  and (_01462_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_01463_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_01464_, _01345_, _01276_);
  and (_01465_, _01464_, _01463_);
  or (_01466_, _01465_, _01461_);
  or (_01467_, _01466_, _01455_);
  or (_01468_, _01467_, _01082_);
  and (_01469_, _01468_, _01446_);
  or (_01470_, _01469_, _01089_);
  nand (_01471_, _01089_, _01064_);
  and (_01472_, _01471_, _05552_);
  and (_13364_, _01472_, _01470_);
  or (_01473_, _01382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_01474_, _01448_, _01385_);
  and (_01475_, _01474_, _01473_);
  nor (_01476_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_01477_, _01476_, _01456_);
  and (_01478_, _01477_, _01357_);
  or (_01479_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_01481_, _01462_, _01276_);
  and (_01482_, _01481_, _01479_);
  or (_01483_, _01482_, _01478_);
  or (_01484_, _01483_, _01475_);
  or (_01485_, _01484_, _01082_);
  nand (_01486_, _01082_, _07945_);
  and (_01487_, _01486_, _01485_);
  or (_01488_, _01487_, _01089_);
  or (_01489_, _01091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_01491_, _01489_, _05552_);
  and (_13370_, _01491_, _01488_);
  and (_01492_, _00245_, _07443_);
  nor (_01494_, _01492_, _13526_);
  and (_01495_, _01492_, _11238_);
  or (_01496_, _01495_, _01494_);
  and (_13376_, _01496_, _05552_);
  nor (_01497_, _01492_, _00146_);
  and (_01498_, _01492_, _11234_);
  or (_01499_, _01498_, _01497_);
  and (_13378_, _01499_, _05552_);
  or (_01500_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_01501_, _01500_, _05552_);
  nand (_01502_, _01492_, _06560_);
  and (_13388_, _01502_, _01501_);
  or (_01503_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_01504_, _01503_, _05552_);
  nand (_01505_, _01492_, _07388_);
  and (_13393_, _01505_, _01504_);
  or (_01506_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_01507_, _01506_, _05552_);
  nand (_01508_, _01492_, _08041_);
  and (_13396_, _01508_, _01507_);
  or (_01509_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_01510_, _01509_, _05552_);
  nand (_01511_, _01492_, _08386_);
  and (_13403_, _01511_, _01510_);
  or (_01512_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_01513_, _01512_, _05552_);
  nand (_01514_, _01492_, _06306_);
  and (_13406_, _01514_, _01513_);
  and (_13470_, _08073_, _05552_);
  and (_01515_, _00224_, _06765_);
  and (_01516_, _01515_, _08635_);
  nand (_01517_, _01516_, _06763_);
  nor (_01518_, _06001_, _05989_);
  and (_01519_, _01518_, _06926_);
  and (_01520_, _01519_, _00240_);
  not (_01521_, _01520_);
  or (_01522_, _01516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01523_, _01522_, _01521_);
  and (_01524_, _01523_, _01517_);
  nor (_01525_, _01521_, _06306_);
  or (_01526_, _01525_, _01524_);
  and (_13483_, _01526_, _05552_);
  and (_01527_, _06054_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01528_, _01527_, _08062_);
  and (_01529_, _01528_, _01515_);
  nor (_01530_, _06059_, _06054_);
  not (_01531_, _01515_);
  or (_01532_, _01531_, _01530_);
  and (_01533_, _01532_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01534_, _01533_, _01520_);
  or (_01535_, _01534_, _01529_);
  nand (_01536_, _01520_, _07388_);
  and (_01537_, _01536_, _05552_);
  and (_13490_, _01537_, _01535_);
  and (_01538_, _01515_, _10632_);
  nand (_01540_, _01538_, _06763_);
  or (_01541_, _01538_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_01543_, _01541_, _01521_);
  and (_01544_, _01543_, _01540_);
  nor (_01546_, _01521_, _06560_);
  or (_01548_, _01546_, _01544_);
  and (_13493_, _01548_, _05552_);
  and (_13506_, _07677_, _05552_);
  and (_01550_, _01515_, _06060_);
  nand (_01551_, _01550_, _06763_);
  or (_01552_, _01550_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01553_, _01552_, _01521_);
  and (_01554_, _01553_, _01551_);
  and (_01555_, _01520_, _11238_);
  or (_01556_, _01555_, _01554_);
  and (_13543_, _01556_, _05552_);
  and (_01557_, _08990_, _06779_);
  or (_01558_, _06770_, _06769_);
  not (_01559_, _01558_);
  and (_01560_, _10860_, _06779_);
  nand (_01561_, _01560_, _01559_);
  and (_01562_, _01561_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01563_, _01562_, _01557_);
  and (_01564_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01565_, _01564_, _08015_);
  and (_01567_, _01565_, _01560_);
  or (_01568_, _01567_, _01563_);
  nand (_01570_, _01557_, _08041_);
  and (_01572_, _01570_, _05552_);
  and (_13558_, _01572_, _01568_);
  not (_01573_, _01557_);
  and (_01574_, _06064_, _05989_);
  and (_01575_, _13693_, _01574_);
  and (_01576_, _01575_, _06765_);
  and (_01577_, _01576_, _06056_);
  or (_01578_, _01577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_01579_, _01578_, _01573_);
  nand (_01580_, _01577_, _06763_);
  and (_01581_, _01580_, _01579_);
  nor (_01582_, _01573_, _07975_);
  or (_01583_, _01582_, _01581_);
  and (_13564_, _01583_, _05552_);
  and (_01585_, _01560_, _06060_);
  or (_01586_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01588_, _01586_, _01573_);
  nand (_01589_, _01585_, _06763_);
  and (_01590_, _01589_, _01588_);
  and (_01591_, _01557_, _11238_);
  or (_01592_, _01591_, _01590_);
  and (_13569_, _01592_, _05552_);
  and (_01595_, _01560_, _08365_);
  or (_01597_, _01595_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_01598_, _01597_, _01573_);
  nand (_01599_, _01595_, _06763_);
  and (_01600_, _01599_, _01598_);
  nor (_01601_, _01573_, _08386_);
  or (_01602_, _01601_, _01600_);
  and (_13580_, _01602_, _05552_);
  and (_01603_, _01560_, _08635_);
  or (_01604_, _01603_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_01605_, _01604_, _01573_);
  nand (_01606_, _01603_, _06763_);
  and (_01607_, _01606_, _01605_);
  nor (_01608_, _01573_, _06306_);
  or (_01609_, _01608_, _01607_);
  and (_13587_, _01609_, _05552_);
  not (_01610_, _01560_);
  or (_01611_, _01610_, _08059_);
  and (_01612_, _01611_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01613_, _01612_, _01557_);
  and (_01614_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01615_, _01614_, _08062_);
  and (_01616_, _01615_, _01560_);
  or (_01617_, _01616_, _01613_);
  nand (_01618_, _01557_, _07388_);
  and (_01619_, _01618_, _05552_);
  and (_13590_, _01619_, _01617_);
  nand (_13680_, _11699_, _05552_);
  nor (_01620_, _07951_, _07388_);
  and (_01621_, _07951_, _06070_);
  or (_01622_, _01621_, _06062_);
  and (_01623_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or (_01624_, _06948_, _06309_);
  or (_01625_, _01624_, _06058_);
  and (_01626_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_01627_, _01626_, _01625_);
  or (_01628_, _01627_, _01623_);
  or (_01629_, _01628_, _01620_);
  and (_13682_, _01629_, _05552_);
  nor (_13709_, _11250_, rst);
  nor (_13714_, _11344_, rst);
  nor (_13717_, _11429_, rst);
  nor (_13720_, _11502_, rst);
  nand (_13726_, _11757_, _05552_);
  and (_01632_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_01633_, _01632_, _13739_);
  and (_01634_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_01635_, _07976_, _06309_);
  or (_01636_, _01635_, _01634_);
  or (_01637_, _01636_, _01633_);
  and (_13761_, _01637_, _05552_);
  and (_01638_, _13740_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_01639_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_01640_, _01639_, _13742_);
  and (_01641_, _09504_, _07946_);
  or (_01642_, _01641_, _01640_);
  or (_01643_, _01642_, _01638_);
  and (_00025_, _01643_, _05552_);
  and (_01644_, _06072_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_01645_, _11490_, _06310_);
  or (_01646_, _01645_, _01644_);
  and (_00060_, _01646_, _05552_);
  and (_01647_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_01648_, _05550_, _11609_);
  or (_01649_, _01648_, _01647_);
  and (_00071_, _01649_, _05552_);
  and (_01650_, _06072_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_01651_, _07439_, _06310_);
  or (_01652_, _01651_, _01650_);
  and (_00076_, _01652_, _05552_);
  and (_00085_, _07522_, _05552_);
  nor (_01653_, _09030_, _06811_);
  and (_01654_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_01655_, _01654_, _01653_);
  and (_00122_, _01655_, _05552_);
  and (_00153_, _07610_, _05552_);
  and (_01656_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_01657_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or (_01658_, _01657_, _01656_);
  and (_00159_, _01658_, _05552_);
  or (_01659_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_01660_, _05550_, _05652_);
  and (_01661_, _01660_, _05552_);
  and (_00201_, _01661_, _01659_);
  and (_00205_, _12169_, _05552_);
  and (_01662_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_01663_, _05550_, _07743_);
  or (_01665_, _01663_, _01662_);
  and (_00206_, _01665_, _05552_);
  and (_01667_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_01668_, _01667_, _13739_);
  and (_01669_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_01670_, _11726_, _06310_);
  or (_01671_, _01670_, _01669_);
  or (_01672_, _01671_, _01668_);
  and (_00219_, _01672_, _05552_);
  and (_00235_, _07454_, _05552_);
  nor (_01673_, _09505_, _06811_);
  and (_01674_, _09505_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_01675_, _01674_, _06955_);
  or (_01676_, _01675_, _01673_);
  or (_01677_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_01678_, _01677_, _05552_);
  and (_00247_, _01678_, _01676_);
  and (_01679_, _11076_, _05886_);
  or (_01681_, _11174_, _05833_);
  or (_01682_, _11155_, _11078_);
  not (_01683_, _11170_);
  or (_01684_, _13392_, _01683_);
  or (_01685_, _01684_, _01682_);
  or (_01687_, _01685_, _01681_);
  and (_01688_, _01687_, _11084_);
  or (_01689_, _01688_, _01679_);
  and (_00251_, _01689_, _05552_);
  nand (_01690_, _10861_, _06056_);
  nor (_01691_, _01690_, _06763_);
  nand (_01692_, _09001_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_01693_, _09012_, _09006_);
  or (_01694_, _01693_, _01692_);
  nand (_01695_, _01694_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_01696_, _01695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01697_, _01696_, _01690_);
  or (_01698_, _01697_, _08991_);
  or (_01699_, _01698_, _01691_);
  nand (_01700_, _08991_, _07975_);
  and (_01701_, _01700_, _05552_);
  and (_00269_, _01701_, _01699_);
  nand (_01702_, _11098_, _05552_);
  nor (_02255_, _01702_, _11141_);
  and (_00271_, _02255_, _11258_);
  nand (_01703_, _10861_, _10632_);
  nor (_01704_, _01703_, _06763_);
  and (_01705_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_01706_, _01692_, _09013_);
  and (_01707_, _01706_, _01705_);
  and (_01708_, _01707_, _01703_);
  or (_01709_, _01708_, _08991_);
  or (_01710_, _01709_, _01704_);
  nand (_01711_, _08991_, _06560_);
  and (_01712_, _01711_, _05552_);
  and (_00274_, _01712_, _01710_);
  or (_01714_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_01715_, _05550_, _05695_);
  and (_01716_, _01715_, _05552_);
  and (_00291_, _01716_, _01714_);
  and (_01717_, _06068_, _06062_);
  nand (_01718_, _01717_, _07945_);
  or (_01719_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_01720_, _01719_, _01718_);
  and (_00328_, _01720_, _05552_);
  and (_00331_, _08113_, _05552_);
  and (_01721_, _01560_, _06771_);
  or (_01722_, _01721_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_01723_, _01722_, _01573_);
  nand (_01724_, _01721_, _06763_);
  and (_01725_, _01724_, _01723_);
  nor (_01726_, _01573_, _06811_);
  or (_01727_, _01726_, _01725_);
  and (_00336_, _01727_, _05552_);
  and (_01728_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_01729_, _01728_, _05576_);
  or (_01730_, _01729_, _06320_);
  and (_01731_, _01730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nand (_01732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_01733_, _01732_, _05586_);
  or (_01734_, _01733_, _13411_);
  or (_01735_, _01734_, _01731_);
  and (_00342_, _01735_, _05552_);
  and (_00475_, _07698_, _05552_);
  or (_01736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_01738_, _10626_, _10860_);
  or (_01739_, _01738_, _01736_);
  not (_01740_, _06771_);
  nor (_01741_, _01740_, _06763_);
  nand (_01742_, _01740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_01743_, _01742_, _01738_);
  or (_01744_, _01743_, _01741_);
  and (_01745_, _01744_, _01739_);
  and (_01746_, _10626_, _08990_);
  or (_01747_, _01746_, _01745_);
  nand (_01748_, _01746_, _06811_);
  and (_01749_, _01748_, _05552_);
  and (_00514_, _01749_, _01747_);
  and (_01750_, _07262_, _06915_);
  nand (_01751_, _01750_, _06060_);
  or (_01752_, _01751_, _07635_);
  not (_01753_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_01754_, _01751_, _01753_);
  and (_01755_, _01754_, _06524_);
  and (_01756_, _01755_, _01752_);
  nor (_01757_, _06774_, _01753_);
  and (_01758_, _01750_, _08635_);
  nand (_01759_, _01758_, _06763_);
  or (_01760_, _01758_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01762_, _01760_, _06775_);
  and (_01763_, _01762_, _01759_);
  or (_01764_, _01763_, _01757_);
  or (_01765_, _01764_, _01756_);
  and (_00530_, _01765_, _05552_);
  or (_01766_, _01751_, _12189_);
  not (_01767_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_01768_, _01751_, _01767_);
  and (_01769_, _01768_, _06524_);
  and (_01770_, _01769_, _01766_);
  nor (_01771_, _06774_, _01767_);
  not (_01772_, _01750_);
  or (_01773_, _01772_, _01530_);
  and (_01774_, _01773_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01775_, _06054_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_01776_, _01775_, _08062_);
  and (_01777_, _01776_, _01750_);
  or (_01778_, _01777_, _01774_);
  and (_01779_, _01778_, _06775_);
  or (_01780_, _01779_, _01771_);
  or (_01781_, _01780_, _01770_);
  and (_00533_, _01781_, _05552_);
  or (_01782_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_01783_, _05550_, _11739_);
  and (_01784_, _01783_, _05552_);
  and (_00549_, _01784_, _01782_);
  not (_01785_, _06321_);
  and (_01786_, _09817_, _01785_);
  or (_01787_, _01729_, _06319_);
  and (_01788_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_01789_, _01788_, _01787_);
  or (_00604_, _01789_, _01786_);
  and (_01790_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01791_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_00606_, _01791_, _05552_);
  nor (_01792_, _00329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_01793_, _01792_, _00330_);
  and (_00682_, _01793_, _00335_);
  nor (_01795_, _00254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_01796_, _01795_, _00329_);
  and (_00684_, _01796_, _00335_);
  and (_01798_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01799_, _05550_, _08689_);
  or (_01800_, _01799_, _01798_);
  and (_00771_, _01800_, _05552_);
  and (_01801_, _01081_, _10626_);
  and (_01802_, _00752_, _10626_);
  nor (_01803_, _01802_, _01801_);
  and (_01804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_01805_, _01804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_01806_, _01805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_01807_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_01808_, _01807_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_01809_, _01808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_01810_, _01809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01811_, _01810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_01812_, _01811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_01813_, _01812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_01814_, _01813_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_01815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_01816_, _01815_, _01814_);
  and (_01818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_01819_, _01818_, _01816_);
  or (_01820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_01821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_01822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01821_);
  and (_01823_, _01822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_01824_, _01823_, _01820_);
  not (_01825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_01826_, _10638_, _01825_);
  and (_01827_, _01826_, _10639_);
  not (_01828_, _01827_);
  and (_01829_, _01828_, _01824_);
  and (_01830_, _01829_, _01819_);
  nand (_01831_, _01830_, _10639_);
  nand (_01832_, _01831_, _01803_);
  or (_01833_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_01834_, _01833_, _05552_);
  and (_00793_, _01834_, _01832_);
  or (_01835_, _01751_, _08144_);
  not (_01836_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_01837_, _01751_, _01836_);
  and (_01838_, _01837_, _06524_);
  and (_01839_, _01838_, _01835_);
  nor (_01840_, _06774_, _01836_);
  nand (_01841_, _01750_, _01559_);
  and (_01842_, _01841_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01843_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_01844_, _01843_, _08015_);
  and (_01845_, _01844_, _01750_);
  or (_01846_, _01845_, _01842_);
  and (_01847_, _01846_, _06775_);
  or (_01848_, _01847_, _01840_);
  or (_01849_, _01848_, _01839_);
  and (_00807_, _01849_, _05552_);
  or (_01850_, _01751_, _08102_);
  not (_01851_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_01852_, _01751_, _01851_);
  and (_01853_, _01852_, _06524_);
  and (_01854_, _01853_, _01850_);
  nor (_01855_, _06774_, _01851_);
  and (_01856_, _01750_, _06056_);
  nand (_01857_, _01856_, _06763_);
  or (_01858_, _01856_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01859_, _01858_, _06775_);
  and (_01860_, _01859_, _01857_);
  or (_01861_, _01860_, _01855_);
  or (_01862_, _01861_, _01854_);
  and (_00815_, _01862_, _05552_);
  and (_00894_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _05552_);
  and (_00910_, _07995_, _05552_);
  not (_01865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_01866_, _10638_, _01865_);
  or (_01867_, _01866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_01868_, _01867_, _01738_);
  nand (_01869_, _08366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_01870_, _01869_, _01738_);
  or (_01871_, _01870_, _08367_);
  and (_01872_, _01871_, _01868_);
  or (_01873_, _01872_, _01746_);
  nand (_01874_, _01746_, _08386_);
  and (_01875_, _01874_, _05552_);
  and (_00917_, _01875_, _01873_);
  not (_01876_, _01746_);
  and (_01877_, _01738_, _08635_);
  or (_01878_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_01879_, _01878_, _01876_);
  nand (_01880_, _01877_, _06763_);
  and (_01881_, _01880_, _01879_);
  nor (_01882_, _01876_, _06306_);
  or (_01883_, _01882_, _01881_);
  and (_00922_, _01883_, _05552_);
  or (_01885_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_01886_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_01888_, pc_log_change, _01886_);
  and (_01889_, _01888_, _05552_);
  and (_00925_, _01889_, _01885_);
  not (_01890_, _01738_);
  or (_01891_, _01890_, _08059_);
  and (_01892_, _01891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_01893_, _01892_, _01746_);
  and (_01894_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_01896_, _01894_, _08062_);
  and (_01897_, _01896_, _01738_);
  or (_01898_, _01897_, _01893_);
  nand (_01900_, _01746_, _07388_);
  and (_01901_, _01900_, _05552_);
  and (_00928_, _01901_, _01898_);
  and (_01902_, _01738_, _10632_);
  or (_01903_, _01902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_01905_, _01903_, _01876_);
  nand (_01906_, _01902_, _06763_);
  and (_01907_, _01906_, _01905_);
  nor (_01908_, _01876_, _06560_);
  or (_01909_, _01908_, _01907_);
  and (_00930_, _01909_, _05552_);
  or (_01910_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not (_01911_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01912_, pc_log_change, _01911_);
  and (_01913_, _01912_, _05552_);
  and (_00933_, _01913_, _01910_);
  or (_01914_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not (_01915_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_01916_, pc_log_change, _01915_);
  and (_01917_, _01916_, _05552_);
  and (_00938_, _01917_, _01914_);
  and (_01919_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_01920_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_01921_, pc_log_change, _01920_);
  or (_01922_, _01921_, _01919_);
  and (_00941_, _01922_, _05552_);
  and (_01923_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_01924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_01925_, pc_log_change, _01924_);
  or (_01926_, _01925_, _01923_);
  and (_00962_, _01926_, _05552_);
  nand (_01927_, _01738_, _01559_);
  and (_01928_, _01927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_01929_, _01928_, _01746_);
  and (_01930_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_01931_, _01930_, _08015_);
  and (_01933_, _01931_, _01738_);
  or (_01934_, _01933_, _01929_);
  nand (_01935_, _01746_, _08041_);
  and (_01936_, _01935_, _05552_);
  and (_00966_, _01936_, _01934_);
  and (_01937_, _01575_, _08007_);
  and (_01938_, _01937_, _06056_);
  or (_01939_, _01938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_01940_, _01939_, _01876_);
  nand (_01941_, _01938_, _06763_);
  and (_01942_, _01941_, _01940_);
  nor (_01943_, _01876_, _07975_);
  or (_01944_, _01943_, _01942_);
  and (_00970_, _01944_, _05552_);
  and (_01945_, _01738_, _06060_);
  or (_01946_, _01945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_01947_, _01946_, _01876_);
  nand (_01948_, _01945_, _06763_);
  and (_01949_, _01948_, _01947_);
  and (_01950_, _01746_, _11238_);
  or (_01951_, _01950_, _01949_);
  and (_00990_, _01951_, _05552_);
  or (_01952_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01953_, pc_log_change, _06192_);
  and (_01954_, _01953_, _05552_);
  and (_00992_, _01954_, _01952_);
  and (_01955_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_01956_, pc_log_change);
  and (_01957_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_01958_, _01957_, _01955_);
  and (_00996_, _01958_, _05552_);
  and (_01959_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_01960_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_01961_, pc_log_change, _01960_);
  or (_01962_, _01961_, _01959_);
  and (_00999_, _01962_, _05552_);
  and (_01963_, _01824_, _01816_);
  and (_01964_, _01963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_01965_, _01963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_01966_, _01965_, _01964_);
  not (_01967_, _10641_);
  and (_01968_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_01969_, _01968_, _01824_);
  and (_01970_, _01969_, _01819_);
  or (_01971_, _01970_, _01827_);
  or (_01972_, _01971_, _01966_);
  or (_01973_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_01974_, _01973_, _01803_);
  and (_01975_, _01974_, _01972_);
  and (_01976_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_01977_, _01976_, _01975_);
  not (_01978_, _01802_);
  nor (_01979_, _01978_, _08386_);
  or (_01980_, _01979_, _01977_);
  and (_01028_, _01980_, _05552_);
  and (_01981_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_01982_, _01824_, _01814_);
  and (_01983_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_01984_, _01983_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_01985_, _01984_, _01963_);
  and (_01986_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_01987_, _01986_, _01824_);
  and (_01988_, _01987_, _01819_);
  or (_01989_, _01988_, _01827_);
  or (_01990_, _01989_, _01985_);
  or (_01991_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_01992_, _01991_, _01803_);
  and (_01993_, _01992_, _01990_);
  nor (_01994_, _01978_, _06306_);
  or (_01995_, _01994_, _01993_);
  or (_01996_, _01995_, _01981_);
  and (_01034_, _01996_, _05552_);
  not (_01997_, _01801_);
  or (_01998_, _01997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_01999_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_02000_, _01983_, _01827_);
  or (_02001_, _02000_, _01801_);
  and (_02002_, _02001_, _01999_);
  and (_02003_, _01827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_02005_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_02006_, _02005_, _01830_);
  or (_02007_, _02006_, _02003_);
  or (_02008_, _02007_, _02002_);
  and (_02009_, _02008_, _01998_);
  or (_02011_, _02009_, _01802_);
  nand (_02013_, _01802_, _07388_);
  and (_02014_, _02013_, _05552_);
  and (_01037_, _02014_, _02011_);
  or (_02015_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_02016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _02016_);
  or (_02018_, _02017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_02019_, _02018_, _01132_);
  or (_02020_, _02019_, _01082_);
  and (_02021_, _02020_, _01091_);
  and (_02022_, _02021_, _02015_);
  nor (_02023_, _01091_, _06811_);
  or (_02024_, _02023_, _02022_);
  and (_01042_, _02024_, _05552_);
  nor (_02025_, _01082_, rst);
  not (_02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_02027_, _01311_, _02026_);
  and (_02028_, _01322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_02029_, _02028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02030_, _02029_, _01311_);
  or (_02031_, _02030_, _02027_);
  nand (_02032_, _02031_, _01357_);
  nor (_02033_, _02032_, _01089_);
  and (_01044_, _02033_, _02025_);
  nand (_02034_, _01082_, _06811_);
  and (_02035_, _01431_, _01317_);
  or (_02036_, _02035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_02037_, _02035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02038_, _02037_, _01385_);
  and (_02039_, _02038_, _02036_);
  nor (_02040_, _01318_, _02016_);
  and (_02041_, _01318_, _02016_);
  or (_02042_, _02041_, _02040_);
  and (_02043_, _02042_, _01357_);
  and (_02044_, _01069_, _01058_);
  and (_02045_, _02044_, _02028_);
  or (_02046_, _02045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02047_, _02044_, _02029_);
  nor (_02048_, _02047_, _01276_);
  and (_02049_, _02048_, _02046_);
  or (_02050_, _02049_, _02043_);
  or (_02051_, _02050_, _02039_);
  or (_02052_, _02051_, _01082_);
  and (_02053_, _02052_, _01091_);
  and (_02054_, _02053_, _02034_);
  and (_02055_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_02056_, _02055_, _02054_);
  and (_01046_, _02056_, _05552_);
  or (_02057_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_02058_, _02057_, _05552_);
  nand (_02059_, _01492_, _06811_);
  and (_01057_, _02059_, _02058_);
  and (_02060_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_02061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_02062_, pc_log_change, _02061_);
  or (_02063_, _02062_, _02060_);
  and (_01062_, _02063_, _05552_);
  or (_02064_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not (_02065_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_02066_, pc_log_change, _02065_);
  and (_02067_, _02066_, _05552_);
  and (_01065_, _02067_, _02064_);
  and (_02068_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02069_, pc_log_change, _01886_);
  or (_02070_, _02069_, _02068_);
  and (_01073_, _02070_, _05552_);
  and (_02071_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_02072_, pc_log_change, _01915_);
  or (_02073_, _02072_, _02071_);
  and (_01077_, _02073_, _05552_);
  and (_01080_, t0_i, _05552_);
  and (_01083_, t1_i, _05552_);
  and (_02075_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_02076_, _01824_, _01819_);
  and (_02077_, _02076_, _02075_);
  not (_02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_02079_, _01824_, _01813_);
  and (_02080_, _02079_, _02078_);
  nor (_02081_, _02080_, _01982_);
  or (_02082_, _02081_, _01827_);
  or (_02083_, _02082_, _02077_);
  nor (_02084_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_02085_, _02084_, _01801_);
  and (_02086_, _02085_, _02083_);
  and (_02087_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_02088_, _02087_, _01802_);
  or (_02090_, _02088_, _02086_);
  nand (_02091_, _01802_, _06560_);
  and (_02092_, _02091_, _05552_);
  and (_01086_, _02092_, _02090_);
  nand (_02093_, _00753_, _06811_);
  and (_02094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_02095_, _02094_, _01011_);
  and (_02096_, _02095_, _00931_);
  and (_02097_, _02096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_02098_, _02097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02099_, _02097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_02100_, _02099_, _00934_);
  and (_02101_, _02100_, _02098_);
  and (_02102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02103_, _02102_, _01012_);
  and (_02104_, _02103_, _00946_);
  or (_02105_, _02104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02106_, _02104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_02107_, _02106_, _00940_);
  and (_02108_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_02109_, _02108_, _02107_);
  and (_02110_, _02109_, _02105_);
  or (_02111_, _02110_, _02101_);
  or (_02112_, _02111_, _00753_);
  and (_02113_, _02112_, _00929_);
  and (_02114_, _02113_, _02093_);
  and (_02115_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02116_, _02115_, _02114_);
  and (_01088_, _02116_, _05552_);
  and (_02118_, _01098_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  or (_02119_, _02118_, _02047_);
  and (_02120_, _02119_, _01275_);
  or (_02121_, _02118_, _01132_);
  or (_02122_, _02118_, _02029_);
  and (_02123_, _02122_, _01333_);
  or (_02124_, _02123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_02125_, _02124_, _02121_);
  nor (_02126_, _02125_, _02120_);
  nor (_02127_, _02126_, _01089_);
  and (_01090_, _02127_, _02025_);
  not (_02128_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_02129_, _00766_, _02128_);
  or (_02130_, _02129_, _02106_);
  and (_02131_, _02130_, _00939_);
  or (_02132_, _02129_, _02099_);
  and (_02133_, _02132_, _00750_);
  and (_02134_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_02135_, _02129_, _00748_);
  or (_02136_, _02135_, _00779_);
  or (_02137_, _02136_, _02134_);
  or (_02138_, _02137_, _02133_);
  or (_02139_, _02138_, _02131_);
  nor (_02140_, _00746_, rst);
  and (_02141_, _02140_, _00952_);
  and (_01092_, _02141_, _02139_);
  nand (_02142_, _00746_, _06811_);
  and (_02143_, _00755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_02144_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_02145_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_02146_, _02145_, _00980_);
  and (_02147_, _02146_, _00757_);
  nor (_02148_, _02147_, _02144_);
  nor (_02149_, _02148_, _00753_);
  or (_02150_, _02149_, _02143_);
  or (_02151_, _02150_, _00746_);
  and (_02152_, _02151_, _05552_);
  and (_01094_, _02152_, _02142_);
  and (_02154_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_02155_, _02154_, _02076_);
  and (_02156_, _01824_, _01812_);
  or (_02157_, _02156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_02158_, _02157_, _02079_);
  or (_02159_, _02158_, _01827_);
  or (_02160_, _02159_, _02155_);
  nor (_02161_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_02162_, _02161_, _01801_);
  and (_02163_, _02162_, _02160_);
  and (_02164_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_02166_, _02164_, _01802_);
  or (_02167_, _02166_, _02163_);
  nand (_02169_, _01802_, _08041_);
  and (_02170_, _02169_, _05552_);
  and (_01097_, _02170_, _02167_);
  and (_02171_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_02172_, _02171_, _02076_);
  and (_02173_, _01824_, _01811_);
  nor (_02174_, _02173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_02175_, _02174_, _02156_);
  or (_02176_, _02175_, _01827_);
  or (_02177_, _02176_, _02172_);
  nor (_02178_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_02179_, _02178_, _01801_);
  and (_02180_, _02179_, _02177_);
  and (_02181_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_02182_, _02181_, _01802_);
  or (_02183_, _02182_, _02180_);
  nand (_02184_, _01802_, _07975_);
  and (_02185_, _02184_, _05552_);
  and (_01103_, _02185_, _02183_);
  nor (_01125_, _11139_, rst);
  or (_02186_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not (_02187_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_02188_, pc_log_change, _02187_);
  and (_02189_, _02188_, _05552_);
  and (_01130_, _02189_, _02186_);
  or (_02191_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_02192_, pc_log_change, _06085_);
  and (_02193_, _02192_, _05552_);
  and (_01135_, _02193_, _02191_);
  and (_02194_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_02195_, _02194_, _02076_);
  and (_02196_, _01824_, _01810_);
  nor (_02197_, _02196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_02198_, _02197_, _02173_);
  or (_02199_, _02198_, _01827_);
  or (_02200_, _02199_, _02195_);
  nor (_02201_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_02202_, _02201_, _01801_);
  and (_02203_, _02202_, _02200_);
  and (_02204_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_02205_, _02204_, _01802_);
  or (_02206_, _02205_, _02203_);
  nand (_02207_, _01802_, _07945_);
  and (_02208_, _02207_, _05552_);
  and (_01143_, _02208_, _02206_);
  and (_02209_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_02210_, pc_log_change, _02187_);
  or (_02211_, _02210_, _02209_);
  and (_01150_, _02211_, _05552_);
  nor (_02212_, _01997_, _08386_);
  and (_02213_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_02214_, _02213_, _02076_);
  and (_02215_, _01824_, _01808_);
  or (_02216_, _02215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_02217_, _01824_, _01809_);
  and (_02218_, _02217_, _02216_);
  or (_02219_, _02218_, _01827_);
  or (_02220_, _02219_, _02214_);
  nor (_02221_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_02222_, _02221_, _01801_);
  and (_02223_, _02222_, _02220_);
  or (_02224_, _02223_, _01802_);
  or (_02225_, _02224_, _02212_);
  or (_02226_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_02227_, _02226_, _05552_);
  and (_01169_, _02227_, _02225_);
  and (_02228_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_02229_, _02228_, _02076_);
  and (_02230_, _01824_, _01807_);
  nor (_02231_, _02230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_02232_, _02231_, _02215_);
  or (_02233_, _02232_, _01827_);
  or (_02234_, _02233_, _02229_);
  nor (_02235_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_02236_, _02235_, _01801_);
  and (_02237_, _02236_, _02234_);
  and (_02239_, _09018_, _06059_);
  and (_02240_, _02239_, _10626_);
  and (_02241_, _02240_, _06524_);
  not (_02242_, _02241_);
  nor (_02243_, _02242_, _06306_);
  or (_02244_, _02243_, _02237_);
  or (_02245_, _02244_, _01802_);
  or (_02246_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_02247_, _02246_, _05552_);
  and (_01182_, _02247_, _02245_);
  and (_02248_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02249_, _02248_, _02076_);
  nand (_02250_, _01824_, _01804_);
  and (_02251_, _02250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_02252_, _02250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_02254_, _02252_, _01827_);
  or (_02256_, _02254_, _02251_);
  or (_02257_, _02256_, _02249_);
  nor (_02258_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor (_02259_, _02258_, _01801_);
  and (_02260_, _02259_, _02257_);
  nor (_02261_, _01997_, _08041_);
  or (_02262_, _02261_, _01802_);
  or (_02263_, _02262_, _02260_);
  or (_02264_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_02265_, _02264_, _05552_);
  and (_01201_, _02265_, _02263_);
  and (_02266_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_02267_, _02266_, _02076_);
  and (_02268_, _01824_, _01806_);
  nor (_02269_, _02268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_02270_, _02269_, _02230_);
  or (_02271_, _02270_, _01827_);
  or (_02272_, _02271_, _02267_);
  nor (_02273_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_02274_, _02273_, _01801_);
  and (_02275_, _02274_, _02272_);
  nor (_02276_, _02242_, _07388_);
  or (_02277_, _02276_, _02275_);
  or (_02278_, _02277_, _01802_);
  or (_02279_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_02280_, _02279_, _05552_);
  and (_01207_, _02280_, _02278_);
  and (_02281_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_02282_, _02281_, _02076_);
  and (_02283_, _01824_, _01805_);
  nor (_02284_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_02285_, _02284_, _02268_);
  or (_02287_, _02285_, _01827_);
  or (_02288_, _02287_, _02282_);
  nor (_02289_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor (_02290_, _02289_, _01801_);
  and (_02291_, _02290_, _02288_);
  nor (_02292_, _01997_, _06560_);
  or (_02293_, _02292_, _01802_);
  or (_02294_, _02293_, _02291_);
  or (_02295_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_02296_, _02295_, _05552_);
  and (_01211_, _02296_, _02294_);
  and (_02297_, _01827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_02298_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_02299_, _02298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_02300_, _02250_, _01828_);
  and (_02301_, _02300_, _02299_);
  or (_02302_, _02301_, _02297_);
  or (_02303_, _02302_, _01801_);
  and (_02304_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_02305_, _02304_, _01830_);
  or (_02306_, _02305_, _02303_);
  nand (_02307_, _01801_, _07975_);
  and (_02308_, _02307_, _02306_);
  or (_02309_, _02308_, _01802_);
  or (_02310_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_02311_, _02310_, _05552_);
  and (_01216_, _02311_, _02309_);
  or (_02312_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_02313_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_02314_, _02313_, _01819_);
  nand (_02315_, _02314_, _02298_);
  and (_02316_, _02315_, _02312_);
  or (_02317_, _02316_, _01827_);
  nor (_02318_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_02319_, _02318_, _01801_);
  and (_02320_, _02319_, _02317_);
  and (_02321_, _01801_, _11238_);
  or (_02322_, _02321_, _01802_);
  or (_02323_, _02322_, _02320_);
  or (_02324_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_02325_, _02324_, _05552_);
  and (_01265_, _02325_, _02323_);
  or (_02326_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_02327_, _05550_, _05770_);
  and (_02329_, _02327_, _05552_);
  and (_01352_, _02329_, _02326_);
  not (_02331_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_02332_, _00258_, _02331_);
  nor (_02333_, _00258_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_02334_, _02333_, _00252_);
  or (_02335_, _02334_, _02332_);
  nor (_02336_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02337_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_02338_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_02339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02340_, _02339_, _02338_);
  and (_02341_, _02340_, _02337_);
  nor (_02342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_02343_, _02342_, _00511_);
  and (_02344_, _02343_, _02331_);
  and (_02345_, _02344_, _02341_);
  nor (_02346_, _02345_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02347_, _02346_, _02336_);
  nand (_02348_, _02347_, _00252_);
  and (_02349_, _02348_, _02335_);
  nor (_02350_, _02349_, _00265_);
  and (_02351_, _00248_, _11238_);
  or (_02352_, _02351_, _02350_);
  and (_01355_, _02352_, _05552_);
  nor (_02354_, _10629_, _10643_);
  and (_02355_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  not (_02356_, _02354_);
  and (_02357_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_02358_, _02357_, _02355_);
  or (_02359_, _02358_, _10635_);
  nand (_02360_, _10635_, _08041_);
  and (_02361_, _02360_, _05552_);
  and (_01363_, _02361_, _02359_);
  nand (_02362_, _10635_, _08386_);
  and (_02363_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_02364_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_02365_, _02364_, _02363_);
  or (_02366_, _02365_, _10635_);
  and (_02367_, _02366_, _05552_);
  and (_01366_, _02367_, _02362_);
  nand (_02368_, _10635_, _06306_);
  and (_02369_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_02370_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_02371_, _02370_, _02369_);
  or (_02372_, _02371_, _10635_);
  and (_02373_, _02372_, _05552_);
  and (_01387_, _02373_, _02368_);
  nand (_02374_, _10635_, _07388_);
  and (_02375_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_02377_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_02379_, _02377_, _02375_);
  or (_02380_, _02379_, _10635_);
  and (_02381_, _02380_, _05552_);
  and (_01391_, _02381_, _02374_);
  nand (_02383_, _10635_, _06560_);
  or (_02384_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nand (_02385_, _02354_, _02078_);
  and (_02386_, _02385_, _02384_);
  or (_02387_, _02386_, _10635_);
  and (_02388_, _02387_, _05552_);
  and (_01395_, _02388_, _02383_);
  or (_02389_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_02390_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_02391_, _02390_, _02389_);
  or (_02392_, _02391_, _10635_);
  nand (_02393_, _10635_, _07975_);
  and (_02394_, _02393_, _05552_);
  and (_01403_, _02394_, _02392_);
  or (_02395_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_02396_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_02397_, _02396_, _02395_);
  or (_02398_, _02397_, _10635_);
  nand (_02399_, _10635_, _07945_);
  and (_02400_, _02399_, _05552_);
  and (_01421_, _02400_, _02398_);
  and (_02401_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02402_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_02403_, pc_log_change, _02402_);
  or (_02404_, _02403_, _02401_);
  and (_01437_, _02404_, _05552_);
  and (_02405_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_02406_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_02407_, pc_log_change, _02406_);
  or (_02408_, _02407_, _02405_);
  and (_01444_, _02408_, _05552_);
  and (_02409_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_02410_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_02411_, pc_log_change, _02410_);
  or (_02412_, _02411_, _02409_);
  and (_01447_, _02412_, _05552_);
  and (_02414_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_02415_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_02416_, pc_log_change, _02415_);
  or (_02417_, _02416_, _02414_);
  and (_01449_, _02417_, _05552_);
  and (_02418_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_02419_, pc_log_change, _02065_);
  or (_02420_, _02419_, _02418_);
  and (_01453_, _02420_, _05552_);
  or (_02421_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_02422_, pc_log_change, _06219_);
  and (_02423_, _02422_, _05552_);
  and (_01459_, _02423_, _02421_);
  nand (_02424_, _10629_, _08386_);
  and (_02425_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_02426_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_02427_, _02426_, _02425_);
  or (_02428_, _02427_, _10629_);
  and (_02429_, _02428_, _10636_);
  and (_02430_, _02429_, _02424_);
  and (_02431_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_02432_, _02431_, _02430_);
  and (_01480_, _02432_, _05552_);
  nand (_02433_, _10629_, _06306_);
  and (_02434_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_02436_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_02437_, _02436_, _02434_);
  or (_02438_, _02437_, _10629_);
  and (_02439_, _02438_, _10636_);
  and (_02440_, _02439_, _02433_);
  and (_02441_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_02442_, _02441_, _02440_);
  and (_01490_, _02442_, _05552_);
  and (_02443_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02444_, pc_log_change, _01911_);
  or (_02445_, _02444_, _02443_);
  and (_01493_, _02445_, _05552_);
  nand (_02446_, _10629_, _07388_);
  and (_02447_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_02448_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_02449_, _02448_, _02447_);
  or (_02451_, _02449_, _10629_);
  and (_02452_, _02451_, _10636_);
  and (_02453_, _02452_, _02446_);
  and (_02454_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_02455_, _02454_, _02453_);
  and (_01539_, _02455_, _05552_);
  nand (_02457_, _10629_, _06560_);
  and (_02459_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_02460_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_02461_, _02460_, _02459_);
  or (_02462_, _02461_, _10629_);
  and (_02463_, _02462_, _10636_);
  and (_02464_, _02463_, _02457_);
  and (_02466_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_02467_, _02466_, _02464_);
  and (_01542_, _02467_, _05552_);
  nand (_02469_, _10629_, _08041_);
  and (_02470_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02472_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_02473_, _02472_, _02470_);
  or (_02475_, _02473_, _10629_);
  and (_02476_, _02475_, _10636_);
  and (_02477_, _02476_, _02469_);
  and (_02478_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_02479_, _02478_, _02477_);
  and (_01545_, _02479_, _05552_);
  nand (_02480_, _10629_, _07975_);
  or (_02481_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_02482_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_02483_, _02482_, _02481_);
  or (_02484_, _02483_, _10629_);
  and (_02485_, _02484_, _10636_);
  and (_02486_, _02485_, _02480_);
  and (_02487_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_02488_, _02487_, _02486_);
  and (_01547_, _02488_, _05552_);
  or (_02489_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_02490_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_02491_, _02490_, _02489_);
  or (_02492_, _02491_, _10629_);
  nand (_02493_, _10629_, _07945_);
  and (_02494_, _02493_, _02492_);
  or (_02495_, _02494_, _10635_);
  or (_02496_, _10636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_02497_, _02496_, _05552_);
  and (_01549_, _02497_, _02495_);
  and (_02499_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_02500_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_02501_, pc_log_change, _02500_);
  or (_02502_, _02501_, _02499_);
  and (_01566_, _02502_, _05552_);
  and (_02504_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_02505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_02506_, pc_log_change, _02505_);
  or (_02507_, _02506_, _02504_);
  and (_01569_, _02507_, _05552_);
  and (_02508_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_02509_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_02510_, _02509_, _02508_);
  and (_01571_, _02510_, _05552_);
  and (_02511_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_02512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_02513_, pc_log_change, _02512_);
  or (_02514_, _02513_, _02511_);
  and (_01584_, _02514_, _05552_);
  and (_02515_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_02516_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02517_, _02516_, _02515_);
  and (_01587_, _02517_, _05552_);
  or (_02518_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand (_02520_, pc_log_change, _02415_);
  and (_02521_, _02520_, _05552_);
  and (_01593_, _02521_, _02518_);
  and (_02522_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_02523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_02524_, pc_log_change, _02523_);
  or (_02525_, _02524_, _02522_);
  and (_01594_, _02525_, _05552_);
  and (_02526_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_02527_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02528_, _02527_, _02526_);
  and (_01596_, _02528_, _05552_);
  and (_01630_, _13647_, _05552_);
  nor (_02529_, _07388_, _06953_);
  and (_02530_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_02531_, _02530_, _06955_);
  or (_02532_, _02531_, _02529_);
  or (_02533_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_02534_, _02533_, _05552_);
  and (_01631_, _02534_, _02532_);
  and (_01761_, _10981_, _05552_);
  and (_02535_, _06691_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_01664_, _02535_, _01761_);
  or (_02538_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  nand (_02539_, _05550_, _10995_);
  and (_02541_, _02539_, _05552_);
  and (_01666_, _02541_, _02538_);
  not (_02542_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_02543_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_02544_, _02543_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not (_02546_, _02544_);
  nor (_02547_, _05560_, _05556_);
  and (_02548_, _02547_, _02546_);
  and (_02549_, _02548_, _05593_);
  nor (_02550_, _02549_, _02542_);
  and (_02551_, _02549_, rxd_i);
  or (_02552_, _02551_, rst);
  or (_01680_, _02552_, _02550_);
  and (_01686_, _12106_, _05552_);
  and (_02553_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_02554_, _02553_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_01713_, _02554_, _05552_);
  and (_01737_, _07998_, _05552_);
  nand (_02555_, _10635_, _06811_);
  and (_02556_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_02557_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_02558_, _02557_, _02556_);
  or (_02559_, _02558_, _10635_);
  and (_02560_, _02559_, _05552_);
  and (_01794_, _02560_, _02555_);
  and (_02561_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_02562_, _05550_, _05907_);
  or (_02563_, _02562_, _02561_);
  and (_01797_, _02563_, _05552_);
  and (_02564_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_02565_, _05550_, _06564_);
  or (_02566_, _02565_, _02564_);
  and (_01817_, _02566_, _05552_);
  and (_01863_, t2ex_i, _05552_);
  nand (_02567_, _05547_, _05605_);
  nand (_02568_, _02567_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_02569_, _02568_, _05917_);
  and (_01864_, _02569_, _05552_);
  and (_02570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _05552_);
  and (_02572_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _05552_);
  and (_02573_, _02572_, _05917_);
  or (_01884_, _02573_, _02570_);
  nor (_02574_, _05550_, _05548_);
  and (_02575_, _00364_, _00361_);
  nor (_02576_, _02575_, _05548_);
  and (_02577_, _02576_, _05542_);
  nor (_02578_, _02576_, _05542_);
  nor (_02579_, _02578_, _02577_);
  nor (_02580_, _02579_, _02574_);
  and (_02581_, _05623_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_02582_, _02581_, _02574_);
  and (_02583_, _02582_, _07929_);
  or (_02584_, _02583_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02585_, _02584_, _02580_);
  and (_01887_, _02585_, _05552_);
  and (_02586_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_02587_, _12264_, _11367_);
  or (_02588_, _02587_, _02586_);
  and (_01895_, _02588_, _05552_);
  nor (_01899_, _11993_, rst);
  and (_02589_, _11102_, _05552_);
  and (_01918_, _02589_, _11774_);
  nand (_02590_, _01717_, _06560_);
  or (_02591_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_02592_, _02591_, _05552_);
  and (_01932_, _02592_, _02590_);
  nor (_02593_, _09030_, _07388_);
  and (_02594_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_02595_, _02594_, _02593_);
  and (_02010_, _02595_, _05552_);
  and (_02596_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_02598_, _09030_, _06560_);
  or (_02599_, _02598_, _02596_);
  and (_02012_, _02599_, _05552_);
  nor (_02600_, t2ex_i, rst);
  and (_02074_, _02600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor (_02089_, _11967_, rst);
  or (_02601_, _12189_, _07668_);
  or (_02602_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_02603_, _02602_, _05552_);
  and (_02153_, _02603_, _02601_);
  and (_02605_, _11367_, _06310_);
  or (_02606_, _13739_, _06070_);
  and (_02607_, _02606_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_02608_, _02607_, _02605_);
  and (_02165_, _02608_, _05552_);
  and (_02610_, _12189_, _07445_);
  and (_02611_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_02613_, _02611_, _07485_);
  or (_02614_, _02613_, _02610_);
  or (_02615_, _12215_, _07579_);
  and (_02616_, _02615_, _05552_);
  and (_02168_, _02616_, _02614_);
  nor (_02617_, _08386_, _06953_);
  and (_02618_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_02619_, _02618_, _06955_);
  or (_02620_, _02619_, _02617_);
  or (_02621_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_02622_, _02621_, _05552_);
  and (_02190_, _02622_, _02620_);
  and (_02238_, _08982_, _05552_);
  not (_02623_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02624_, _02623_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_02253_, _02624_, _05552_);
  and (_02625_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_02626_, _12264_, _11490_);
  or (_02627_, _02626_, _02625_);
  and (_02286_, _02627_, _05552_);
  nand (_02628_, _01717_, _07388_);
  or (_02629_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_02630_, _02629_, _05552_);
  and (_02330_, _02630_, _02628_);
  and (_02631_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_02632_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_02633_, _02632_, _01625_);
  nor (_02634_, _08041_, _07951_);
  or (_02635_, _02634_, _02633_);
  or (_02637_, _02635_, _02631_);
  and (_02353_, _02637_, _05552_);
  nor (_02376_, _11448_, rst);
  and (_02638_, _05607_, _05545_);
  and (_02639_, _02638_, _05884_);
  and (_02640_, _07865_, _07784_);
  or (_02641_, _02640_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_02642_, _07788_, _05756_);
  and (_02643_, _07898_, _02642_);
  not (_02644_, _05733_);
  and (_02645_, _07805_, _07788_);
  and (_02646_, _07865_, _07810_);
  or (_02647_, _02646_, _02645_);
  and (_02648_, _02647_, _02644_);
  or (_02649_, _02648_, _02643_);
  or (_02650_, _02649_, _02641_);
  and (_02651_, _02650_, _02639_);
  nor (_02652_, _02638_, _05884_);
  or (_02653_, _02652_, rst);
  or (_02378_, _02653_, _02651_);
  nor (_02382_, _11390_, rst);
  nand (_02655_, _07945_, _06949_);
  or (_02656_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_02657_, _02656_, _02655_);
  and (_02413_, _02657_, _05552_);
  nor (_02658_, t2_i, rst);
  and (_02435_, _02658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and (_02659_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_02660_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or (_02661_, _02660_, _02659_);
  and (_02450_, _02661_, _05552_);
  and (_02456_, _13668_, _05552_);
  and (_02458_, _13636_, _05552_);
  and (_02662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _05556_);
  and (_02663_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02664_, _02663_, _02662_);
  and (_02465_, _02664_, _05552_);
  and (_02665_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _05556_);
  and (_02666_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02667_, _02666_, _02665_);
  and (_02468_, _02667_, _05552_);
  and (_02669_, _11214_, _06310_);
  and (_02670_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_02671_, _02670_, _13739_);
  and (_02672_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_02673_, _02672_, _02671_);
  or (_02674_, _02673_, _02669_);
  and (_02471_, _02674_, _05552_);
  and (_02675_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_02474_, _02675_, _05591_);
  and (_02498_, _02570_, _00580_);
  nand (_02676_, _01717_, _08386_);
  or (_02678_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02679_, _02678_, _05552_);
  and (_02503_, _02679_, _02676_);
  nor (_02519_, _08986_, rst);
  and (_02680_, _06068_, _06058_);
  not (_02681_, _02680_);
  and (_02682_, _02681_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_02683_, _02680_, _11234_);
  or (_02684_, _02683_, _02682_);
  and (_02536_, _02684_, _05552_);
  and (_02685_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_02686_, _02685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_02537_, _02686_, _05552_);
  and (_02687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _05556_);
  and (_02688_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02689_, _02688_, _02687_);
  and (_02540_, _02689_, _05552_);
  nand (_02690_, _01717_, _06306_);
  or (_02691_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_02692_, _02691_, _05552_);
  and (_02545_, _02692_, _02690_);
  or (_02693_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_02694_, _05550_, _05615_);
  and (_02695_, _02694_, _05552_);
  and (_02571_, _02695_, _02693_);
  and (_02597_, _05669_, _05552_);
  and (_02696_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_02697_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_02698_, pc_log_change, _02697_);
  or (_02699_, _02698_, _02696_);
  and (_02604_, _02699_, _05552_);
  nand (_02700_, _01717_, _07975_);
  or (_02701_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_02702_, _02701_, _02700_);
  and (_02609_, _02702_, _05552_);
  nand (_02703_, _01717_, _08041_);
  or (_02704_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_02705_, _02704_, _05552_);
  and (_02612_, _02705_, _02703_);
  nor (_02707_, _00613_, _00580_);
  or (_02709_, _02707_, _08998_);
  nand (_02710_, _01234_, _00833_);
  and (_02711_, _02710_, _05552_);
  and (_02636_, _02711_, _02709_);
  and (_02712_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_02713_, _02712_, _08015_);
  and (_02714_, _02713_, _01515_);
  nand (_02715_, _01515_, _01559_);
  and (_02716_, _02715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_02717_, _02716_, _01520_);
  or (_02718_, _02717_, _02714_);
  nand (_02719_, _01520_, _08041_);
  and (_02720_, _02719_, _05552_);
  and (_02654_, _02720_, _02718_);
  or (_02721_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02722_, _02721_, _00636_);
  not (_02723_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_02724_, _00864_, _02723_);
  nand (_02725_, _02724_, _00863_);
  or (_02727_, _00644_, _08999_);
  and (_02728_, _02727_, _02725_);
  or (_02729_, _02728_, _00641_);
  or (_02730_, _02721_, _01223_);
  and (_02731_, _02730_, _01222_);
  and (_02732_, _02731_, _02729_);
  and (_02733_, _00639_, _08999_);
  or (_02734_, _02733_, _00635_);
  or (_02735_, _02734_, _02732_);
  and (_02737_, _02735_, _02722_);
  or (_02738_, _02737_, _00649_);
  or (_02740_, _02721_, _00603_);
  or (_02741_, _00846_, _02723_);
  nand (_02742_, _02741_, _00845_);
  or (_02743_, _00599_, _08999_);
  and (_02744_, _02743_, _02742_);
  or (_02745_, _02744_, _00609_);
  or (_02746_, _02721_, _01204_);
  and (_02747_, _02746_, _01203_);
  and (_02748_, _02747_, _02745_);
  and (_02749_, _00607_, _08999_);
  or (_02750_, _02749_, _00602_);
  or (_02751_, _02750_, _02748_);
  and (_02752_, _02751_, _02740_);
  or (_02753_, _02752_, _00857_);
  and (_02754_, _02753_, _02738_);
  or (_02755_, _02754_, _00580_);
  or (_02756_, _01235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_02757_, _02756_, _05552_);
  and (_02668_, _02757_, _02755_);
  and (_02758_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_02759_, _02758_, _01235_);
  and (_02677_, _02759_, _05552_);
  and (_02706_, _08976_, _05552_);
  or (_02760_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_02761_, _05550_, _05791_);
  and (_02762_, _02761_, _05552_);
  and (_02708_, _02762_, _02760_);
  and (_02763_, _00225_, _06771_);
  nand (_02764_, _02763_, _06763_);
  or (_02765_, _02763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_02767_, _02765_, _00451_);
  and (_02768_, _02767_, _02764_);
  nor (_02769_, _00451_, _06811_);
  or (_02770_, _02769_, _02768_);
  and (_02726_, _02770_, _05552_);
  and (_02771_, _02336_, _00257_);
  and (_02772_, _02771_, _02343_);
  and (_02773_, _02772_, _02341_);
  not (_02774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_02775_, _00257_, _02774_);
  or (_02776_, _02775_, _02773_);
  and (_02777_, _02776_, _00254_);
  nand (_02778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_02780_, _02778_, _00253_);
  nor (_02781_, _02780_, _02777_);
  nor (_02782_, _02781_, _00252_);
  and (_02783_, _02345_, _00252_);
  or (_02784_, _02783_, _02782_);
  and (_02736_, _02784_, _00335_);
  not (_02785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_02786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_02787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_02788_, _10874_, _02787_);
  or (_02789_, _02788_, _12099_);
  nor (_02790_, _02789_, _02786_);
  nand (_02791_, _02790_, _02785_);
  nor (_02792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_02793_, _02792_, _02790_);
  nand (_02794_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_02795_, _02794_, _02793_);
  and (_02796_, _02795_, _05552_);
  and (_02739_, _02796_, _02791_);
  or (_02797_, _00333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_02798_, _00333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02799_, _02798_, _02797_);
  and (_02766_, _02799_, _00335_);
  or (_02800_, _02542_, rxd_i);
  nand (_02801_, _02800_, _05574_);
  or (_02802_, _05575_, _05561_);
  and (_02803_, _02802_, _02801_);
  or (_02804_, _05580_, _05572_);
  or (_02806_, _02804_, _05562_);
  or (_02807_, _02806_, _02803_);
  and (_02779_, _02807_, _05585_);
  and (_02808_, _01560_, _10632_);
  or (_02809_, _02808_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_02810_, _02809_, _01573_);
  nand (_02811_, _02808_, _06763_);
  and (_02812_, _02811_, _02810_);
  nor (_02813_, _01573_, _06560_);
  or (_02814_, _02813_, _02812_);
  and (_02805_, _02814_, _05552_);
  and (_02816_, _01515_, _06056_);
  nand (_02817_, _02816_, _06763_);
  or (_02819_, _02816_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_02820_, _02819_, _01521_);
  and (_02822_, _02820_, _02817_);
  nor (_02823_, _01521_, _07975_);
  or (_02824_, _02823_, _02822_);
  and (_02815_, _02824_, _05552_);
  and (_02825_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_02826_, _12264_, _11726_);
  or (_02827_, _02826_, _02825_);
  and (_02818_, _02827_, _05552_);
  and (_02828_, _01515_, _08365_);
  nand (_02829_, _02828_, _06763_);
  or (_02830_, _02828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_02832_, _02830_, _01521_);
  and (_02833_, _02832_, _02829_);
  nor (_02835_, _01521_, _08386_);
  or (_02837_, _02835_, _02833_);
  and (_02821_, _02837_, _05552_);
  and (_02831_, _02793_, _05552_);
  or (_02839_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_02840_, _02839_, _05552_);
  or (_02841_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and (_02842_, _02841_, _05568_);
  or (_02843_, _02842_, _05582_);
  nand (_02844_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nor (_02845_, _02844_, _05582_);
  or (_02846_, _02845_, rxd_i);
  and (_02847_, _02846_, _02843_);
  and (_02848_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_02849_, _02848_, _02847_);
  and (_02834_, _02849_, _02840_);
  nand (_02852_, _02773_, _00253_);
  nand (_02854_, _02852_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02855_, _02854_, _02783_);
  or (_02856_, _02855_, _00265_);
  and (_02836_, _02856_, _05552_);
  or (_02857_, _05803_, _08675_);
  or (_02858_, _05546_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_02859_, _02858_, _05552_);
  and (_02838_, _02859_, _02857_);
  nand (_02860_, _05756_, _05546_);
  or (_02861_, _05546_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_02862_, _02861_, _05552_);
  and (_02850_, _02862_, _02860_);
  nand (_02863_, _00241_, _06811_);
  or (_02864_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_02865_, _02864_, _05552_);
  and (_02851_, _02865_, _02863_);
  and (_02866_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_02868_, _02866_, _00335_);
  and (_02869_, _00246_, _05552_);
  and (_02870_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_02853_, _02870_, _02868_);
  nand (_02871_, _00645_, _00621_);
  nor (_02872_, _02871_, _00613_);
  and (_02873_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or (_02874_, _00598_, _00580_);
  nor (_02875_, _02874_, _00586_);
  not (_02876_, _00611_);
  nor (_02877_, _02876_, _00596_);
  and (_02878_, _02877_, _02875_);
  or (_02879_, _02878_, _02873_);
  or (_02880_, _02879_, _02872_);
  and (_02867_, _02880_, _05552_);
  and (_02881_, _10861_, _08057_);
  or (_02882_, _02881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_02883_, _02882_, _08992_);
  nand (_02884_, _02881_, _06763_);
  and (_02885_, _02884_, _02883_);
  nor (_02886_, _08992_, _07388_);
  or (_02887_, _02886_, _02885_);
  and (_02889_, _02887_, _05552_);
  and (_02888_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_02890_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_02891_, _02890_, _02888_);
  and (_02892_, _02891_, _00335_);
  nand (_02893_, _06560_, _05560_);
  nand (_02894_, _08041_, _05573_);
  and (_02895_, _02894_, _02869_);
  and (_02896_, _02895_, _02893_);
  or (_03014_, _02896_, _02892_);
  and (_02897_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_02898_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_02899_, _02898_, _02897_);
  and (_02900_, _02899_, _00335_);
  nand (_02901_, _08041_, _05560_);
  nand (_02902_, _07975_, _05573_);
  and (_02903_, _02902_, _02869_);
  and (_02904_, _02903_, _02901_);
  or (_03048_, _02904_, _02900_);
  and (_02905_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_02906_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_02907_, _02906_, _02905_);
  and (_02908_, _02907_, _00335_);
  or (_02909_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _12098_);
  and (_02910_, _02909_, _05552_);
  and (_02911_, _02910_, _00267_);
  or (_03075_, _02911_, _02908_);
  nand (_02912_, _01802_, _06811_);
  or (_02913_, _01964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_02914_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_02915_, _02914_, _01824_);
  nand (_02916_, _02915_, _01819_);
  and (_02917_, _02916_, _02913_);
  or (_02918_, _02917_, _01827_);
  nor (_02919_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_02920_, _02919_, _01801_);
  and (_02921_, _02920_, _02918_);
  nor (_02922_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_02923_, _02922_, _01803_);
  or (_02924_, _02923_, _02921_);
  and (_02925_, _02924_, _05552_);
  and (_03078_, _02925_, _02912_);
  and (_02926_, _01519_, _06061_);
  nand (_02927_, _02926_, _06763_);
  or (_02928_, _02926_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_02929_, _02928_, _06775_);
  and (_02930_, _02929_, _02927_);
  and (_02931_, _02926_, _11238_);
  nor (_02932_, _02926_, _13607_);
  or (_02933_, _02932_, _02931_);
  and (_02934_, _02933_, _06524_);
  nor (_02935_, _06774_, _13607_);
  or (_02936_, _02935_, rst);
  or (_02937_, _02936_, _02934_);
  or (_03126_, _02937_, _02930_);
  and (_02938_, _08365_, _06768_);
  nand (_02939_, _02938_, _06763_);
  or (_02940_, _02938_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_02941_, _02940_, _06775_);
  and (_02942_, _02941_, _02939_);
  nor (_02943_, _08386_, _06782_);
  and (_02944_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02945_, _02944_, _02943_);
  and (_02946_, _02945_, _06524_);
  and (_02947_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02948_, _02947_, rst);
  or (_02949_, _02948_, _02946_);
  or (_03128_, _02949_, _02942_);
  and (_02950_, _06916_, _08013_);
  nand (_02951_, _02950_, _06763_);
  or (_02952_, _02950_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02953_, _02952_, _06775_);
  and (_02954_, _02953_, _02951_);
  nand (_02955_, _08041_, _06928_);
  or (_02956_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02957_, _02956_, _06524_);
  and (_02958_, _02957_, _02955_);
  and (_02959_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_02960_, _02959_, rst);
  or (_02961_, _02960_, _02958_);
  or (_03132_, _02961_, _02954_);
  or (_02962_, _06781_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_02963_, _02962_, _06775_);
  nand (_02964_, _06781_, _06763_);
  and (_02965_, _02964_, _02963_);
  and (_02966_, _11238_, _06781_);
  nor (_02967_, _06781_, _13613_);
  or (_02968_, _02967_, _02966_);
  and (_02969_, _02968_, _06524_);
  nor (_02970_, _06774_, _13613_);
  or (_02971_, _02970_, rst);
  or (_02972_, _02971_, _02969_);
  or (_03134_, _02972_, _02965_);
  and (_02973_, _06910_, _06767_);
  nand (_02974_, _02973_, _06054_);
  and (_02975_, _02974_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_02976_, _01558_, _00021_);
  or (_02977_, _02976_, _12129_);
  and (_02978_, _02977_, _02973_);
  or (_02979_, _02978_, _02975_);
  and (_02980_, _02979_, _06775_);
  and (_02981_, _07443_, _06061_);
  nand (_02982_, _02981_, _06560_);
  or (_02983_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02984_, _02983_, _06524_);
  and (_02985_, _02984_, _02982_);
  nor (_02986_, _06774_, _00021_);
  or (_02987_, _02986_, rst);
  or (_02988_, _02987_, _02985_);
  or (_03136_, _02988_, _02980_);
  or (_02989_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_02990_, _02989_, _06775_);
  nand (_02991_, _02981_, _06763_);
  and (_02992_, _02991_, _02990_);
  nand (_02993_, _07945_, _02981_);
  and (_02994_, _02989_, _06524_);
  and (_02995_, _02994_, _02993_);
  nor (_02996_, _06774_, _13594_);
  or (_02997_, _02996_, rst);
  or (_02998_, _02997_, _02995_);
  or (_03138_, _02998_, _02992_);
  and (_02999_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_03000_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_03001_, _03000_, _02999_);
  or (_03002_, _03001_, _00265_);
  and (_03003_, _03002_, _05552_);
  nand (_03004_, _00267_, _06811_);
  and (_03153_, _03004_, _03003_);
  and (_03005_, _06915_, _06765_);
  and (_03006_, _03005_, _08635_);
  nand (_03007_, _03006_, _06763_);
  or (_03008_, _03006_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03009_, _03008_, _06775_);
  and (_03010_, _03009_, _03007_);
  not (_03011_, _02926_);
  nor (_03012_, _03011_, _06306_);
  and (_03013_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_03015_, _03013_, _03012_);
  and (_03016_, _03015_, _06524_);
  and (_03017_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_03018_, _03017_, rst);
  or (_03019_, _03018_, _03016_);
  or (_03158_, _03019_, _03010_);
  and (_03020_, _08635_, _06768_);
  nand (_03021_, _03020_, _06763_);
  or (_03022_, _03020_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03023_, _03022_, _06775_);
  and (_03024_, _03023_, _03021_);
  nor (_03025_, _06782_, _06306_);
  and (_03026_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_03027_, _03026_, _03025_);
  and (_03028_, _03027_, _06524_);
  and (_03029_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_03030_, _03029_, rst);
  or (_03031_, _03030_, _03028_);
  or (_03160_, _03031_, _03024_);
  and (_03032_, _06916_, _08365_);
  nand (_03033_, _03032_, _06763_);
  or (_03034_, _03032_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03035_, _03034_, _06775_);
  and (_03036_, _03035_, _03033_);
  nand (_03037_, _08386_, _06928_);
  or (_03038_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03039_, _03038_, _06524_);
  and (_03040_, _03039_, _03037_);
  and (_03041_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_03042_, _03041_, rst);
  or (_03043_, _03042_, _03040_);
  or (_03162_, _03043_, _03036_);
  and (_03044_, _06916_, _06056_);
  nand (_03045_, _03044_, _06763_);
  or (_03046_, _03044_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03047_, _03046_, _06775_);
  and (_03049_, _03047_, _03045_);
  nand (_03050_, _07975_, _06928_);
  or (_03051_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03052_, _03051_, _06524_);
  and (_03053_, _03052_, _03050_);
  and (_03054_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_03055_, _03054_, rst);
  or (_03056_, _03055_, _03053_);
  or (_03164_, _03056_, _03049_);
  and (_03057_, _06916_, _08057_);
  nand (_03058_, _03057_, _06763_);
  or (_03059_, _03057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03060_, _03059_, _06775_);
  and (_03061_, _03060_, _03058_);
  nand (_03062_, _07388_, _06928_);
  or (_03063_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03064_, _03063_, _06524_);
  and (_03065_, _03064_, _03062_);
  nor (_03066_, _06774_, _13815_);
  or (_03067_, _03066_, rst);
  or (_03068_, _03067_, _03065_);
  or (_03167_, _03068_, _03061_);
  nand (_03069_, _02973_, _01559_);
  and (_03070_, _03069_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03071_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_03072_, _03071_, _08015_);
  and (_03073_, _03072_, _02973_);
  or (_03074_, _03073_, _03070_);
  and (_03076_, _03074_, _06775_);
  nand (_03077_, _08041_, _02981_);
  or (_03079_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03080_, _03079_, _06524_);
  and (_03081_, _03080_, _03077_);
  and (_03082_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_03083_, _03082_, rst);
  or (_03084_, _03083_, _03081_);
  or (_03170_, _03084_, _03076_);
  and (_03085_, _02973_, _08635_);
  nand (_03086_, _03085_, _06763_);
  or (_03087_, _03085_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03088_, _03087_, _06775_);
  and (_03089_, _03088_, _03086_);
  nand (_03090_, _02981_, _06306_);
  or (_03091_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03092_, _03091_, _06524_);
  and (_03093_, _03092_, _03090_);
  and (_03094_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_03095_, _03094_, rst);
  or (_03096_, _03095_, _03093_);
  or (_03172_, _03096_, _03089_);
  and (_03097_, _08057_, _06768_);
  nand (_03098_, _03097_, _06763_);
  or (_03099_, _03097_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03100_, _03099_, _06775_);
  and (_03101_, _03100_, _03098_);
  nor (_03102_, _07388_, _06782_);
  nor (_03103_, _06781_, _13799_);
  or (_03104_, _03103_, _03102_);
  and (_03105_, _03104_, _06524_);
  nor (_03106_, _06774_, _13799_);
  or (_03107_, _03106_, rst);
  or (_03108_, _03107_, _03105_);
  or (_03256_, _03108_, _03101_);
  and (_03109_, _10632_, _06768_);
  nand (_03110_, _03109_, _06763_);
  or (_03111_, _03109_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03112_, _03111_, _06775_);
  and (_03113_, _03112_, _03110_);
  nor (_03114_, _06782_, _06560_);
  nor (_03115_, _06781_, _00038_);
  or (_03116_, _03115_, _03114_);
  and (_03117_, _03116_, _06524_);
  nor (_03118_, _06774_, _00038_);
  or (_03119_, _03118_, rst);
  or (_03120_, _03119_, _03117_);
  or (_03257_, _03120_, _03113_);
  nor (_03121_, _09030_, _08041_);
  and (_03122_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_03123_, _03122_, _03121_);
  and (_03270_, _03123_, _05552_);
  and (_03124_, _08013_, _06768_);
  nand (_03125_, _03124_, _06763_);
  or (_03127_, _03124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03129_, _03127_, _06775_);
  and (_03130_, _03129_, _03125_);
  nor (_03131_, _08041_, _06782_);
  and (_03133_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_03135_, _03133_, _03131_);
  and (_03137_, _03135_, _06524_);
  and (_03139_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_03140_, _03139_, rst);
  or (_03141_, _03140_, _03137_);
  or (_03281_, _03141_, _03130_);
  and (_03142_, _06916_, _06060_);
  nand (_03143_, _03142_, _06763_);
  or (_03144_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_03145_, _03144_, _06775_);
  and (_03146_, _03145_, _03143_);
  nand (_03147_, _07945_, _06928_);
  and (_03148_, _03147_, _06524_);
  and (_03149_, _03148_, _03144_);
  nor (_03150_, _06774_, _13600_);
  or (_03151_, _03150_, rst);
  or (_03152_, _03151_, _03149_);
  or (_03283_, _03152_, _03146_);
  and (_03154_, _03005_, _10632_);
  nand (_03155_, _03154_, _06763_);
  or (_03156_, _03154_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03157_, _03156_, _06775_);
  and (_03159_, _03157_, _03155_);
  nor (_03161_, _03011_, _06560_);
  nor (_03163_, _02926_, _00033_);
  or (_03165_, _03163_, _03161_);
  and (_03166_, _03165_, _06524_);
  nor (_03168_, _06774_, _00033_);
  or (_03169_, _03168_, rst);
  or (_03171_, _03169_, _03166_);
  or (_03286_, _03171_, _03159_);
  and (_03173_, _03005_, _08013_);
  nand (_03174_, _03173_, _06763_);
  or (_03175_, _03173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03176_, _03175_, _06775_);
  and (_03177_, _03176_, _03174_);
  nor (_03178_, _03011_, _08041_);
  and (_03179_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_03180_, _03179_, _03178_);
  and (_03181_, _03180_, _06524_);
  and (_03182_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_03183_, _03182_, rst);
  or (_03184_, _03183_, _03181_);
  or (_03287_, _03184_, _03177_);
  nand (_03185_, _11223_, _06763_);
  or (_03186_, _11223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03187_, _03186_, _06775_);
  and (_03188_, _03187_, _03185_);
  nand (_03189_, _07975_, _02981_);
  or (_03190_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03191_, _03190_, _06524_);
  and (_03192_, _03191_, _03189_);
  and (_03193_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_03194_, _03193_, rst);
  or (_03195_, _03194_, _03192_);
  or (_03305_, _03195_, _03188_);
  and (_03196_, _02973_, _08365_);
  nand (_03197_, _03196_, _06763_);
  or (_03198_, _03196_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03199_, _03198_, _06775_);
  and (_03200_, _03199_, _03197_);
  nand (_03201_, _08386_, _02981_);
  or (_03202_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03203_, _03202_, _06524_);
  and (_03204_, _03203_, _03201_);
  and (_03205_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_03206_, _03205_, rst);
  or (_03207_, _03206_, _03204_);
  or (_03307_, _03207_, _03200_);
  and (_03208_, _02973_, _08057_);
  nand (_03209_, _03208_, _06763_);
  or (_03210_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03211_, _03210_, _06775_);
  and (_03212_, _03211_, _03209_);
  nand (_03213_, _07388_, _02981_);
  or (_03214_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03215_, _03214_, _06524_);
  and (_03216_, _03215_, _03213_);
  nor (_03217_, _06774_, _13810_);
  or (_03218_, _03217_, rst);
  or (_03219_, _03218_, _03216_);
  or (_03309_, _03219_, _03212_);
  nand (_03220_, _06768_, _06056_);
  nand (_03221_, _03220_, _00173_);
  and (_03222_, _03221_, _06775_);
  or (_03223_, _03220_, _08048_);
  and (_03224_, _03223_, _03222_);
  nor (_03225_, _07975_, _06782_);
  nor (_03226_, _06781_, _00173_);
  or (_03227_, _03226_, _03225_);
  and (_03228_, _03227_, _06524_);
  nor (_03229_, _06774_, _00173_);
  or (_03230_, _03229_, rst);
  or (_03231_, _03230_, _03228_);
  or (_03311_, _03231_, _03224_);
  and (_03232_, _06916_, _08635_);
  nand (_03233_, _03232_, _06763_);
  or (_03234_, _03232_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03235_, _03234_, _06775_);
  and (_03236_, _03235_, _03233_);
  nand (_03237_, _06928_, _06306_);
  or (_03238_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03239_, _03238_, _06524_);
  and (_03240_, _03239_, _03237_);
  and (_03241_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_03242_, _03241_, rst);
  or (_03243_, _03242_, _03240_);
  or (_03312_, _03243_, _03236_);
  and (_03244_, _06916_, _10632_);
  nand (_03245_, _03244_, _06763_);
  or (_03246_, _03244_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03247_, _03246_, _06775_);
  and (_03248_, _03247_, _03245_);
  nand (_03249_, _06928_, _06560_);
  or (_03250_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03251_, _03250_, _06524_);
  and (_03252_, _03251_, _03249_);
  nor (_03253_, _06774_, _00027_);
  or (_03254_, _03253_, rst);
  or (_03255_, _03254_, _03252_);
  or (_03314_, _03255_, _03248_);
  and (_03258_, _03005_, _06056_);
  nand (_03259_, _03258_, _06763_);
  or (_03260_, _03258_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03261_, _03260_, _06775_);
  and (_03262_, _03261_, _03259_);
  nor (_03263_, _03011_, _07975_);
  and (_03264_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_03265_, _03264_, _03263_);
  and (_03266_, _03265_, _06524_);
  and (_03267_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_03268_, _03267_, rst);
  or (_03269_, _03268_, _03266_);
  or (_03317_, _03269_, _03262_);
  and (_03271_, _03005_, _08365_);
  nand (_03272_, _03271_, _06763_);
  or (_03273_, _03271_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03274_, _03273_, _06775_);
  and (_03275_, _03274_, _03272_);
  nor (_03277_, _03011_, _08386_);
  and (_03278_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_03279_, _03278_, _03277_);
  and (_03280_, _03279_, _06524_);
  and (_03282_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_03284_, _03282_, rst);
  or (_03285_, _03284_, _03280_);
  or (_03320_, _03285_, _03275_);
  and (_03288_, _03005_, _08057_);
  nand (_03289_, _03288_, _06763_);
  or (_03290_, _03288_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03291_, _03290_, _06775_);
  and (_03292_, _03291_, _03289_);
  nor (_03293_, _03011_, _07388_);
  nor (_03294_, _02926_, _13804_);
  or (_03295_, _03294_, _03293_);
  and (_03296_, _03295_, _06524_);
  nor (_03297_, _06774_, _13804_);
  or (_03298_, _03297_, rst);
  or (_03299_, _03298_, _03296_);
  or (_03322_, _03299_, _03292_);
  nand (_03300_, _01717_, _06811_);
  or (_03301_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_03302_, _03301_, _05552_);
  and (_03324_, _03302_, _03300_);
  not (_03303_, _00833_);
  or (_03304_, _03303_, _00652_);
  and (_03306_, _00833_, _00629_);
  or (_03308_, _03306_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_03310_, _03308_, _05552_);
  and (_03329_, _03310_, _03304_);
  nor (_03313_, _06811_, _06953_);
  and (_03315_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03316_, _03315_, _06955_);
  or (_03318_, _03316_, _03313_);
  or (_03319_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03321_, _03319_, _05552_);
  and (_03332_, _03321_, _03318_);
  or (_03323_, _05586_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_03325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_03326_, _03325_, _05560_);
  or (_03327_, _03326_, _05562_);
  nand (_03328_, _03327_, _03323_);
  nand (_03346_, _03328_, _05585_);
  or (_03330_, _05710_, _08675_);
  or (_03331_, _05546_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_03333_, _03331_, _05552_);
  and (_03347_, _03333_, _03330_);
  and (_03334_, _07485_, _07360_);
  or (_03335_, _07445_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_03336_, _03335_, _07579_);
  or (_03337_, _07486_, _07255_);
  and (_03338_, _03337_, _03336_);
  or (_03339_, _03338_, _03334_);
  and (_03398_, _03339_, _05552_);
  or (_03340_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_03341_, _05550_, _05768_);
  and (_03342_, _03341_, _05552_);
  and (_03415_, _03342_, _03340_);
  nor (_03424_, _11327_, rst);
  and (_03343_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_03344_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_03345_, _03344_, _03343_);
  and (_03428_, _03345_, _05552_);
  nor (_03433_, _11370_, rst);
  nor (_03436_, _11418_, rst);
  nor (_03439_, _11492_, rst);
  nor (_03441_, _11217_, rst);
  nand (_03348_, _06949_, _06811_);
  or (_03349_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_03350_, _03349_, _05552_);
  and (_03446_, _03350_, _03348_);
  or (_03351_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_03352_, _05550_, _05656_);
  and (_03353_, _03352_, _05552_);
  and (_03454_, _03353_, _03351_);
  nor (_03467_, _11848_, rst);
  nor (_03354_, _01997_, _06811_);
  and (_03355_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_03356_, _03355_, _02076_);
  not (_03357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_03358_, _02217_, _03357_);
  nor (_03359_, _03358_, _02196_);
  or (_03360_, _03359_, _01827_);
  or (_03361_, _03360_, _03356_);
  nor (_03362_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_03363_, _03362_, _01801_);
  and (_03364_, _03363_, _03361_);
  or (_03365_, _03364_, _01802_);
  or (_03366_, _03365_, _03354_);
  nand (_03367_, _01802_, _03357_);
  and (_03368_, _03367_, _05552_);
  and (_03493_, _03368_, _03366_);
  and (_03495_, t2_i, _05552_);
  nand (_03369_, _00241_, _07975_);
  or (_03370_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_03371_, _03370_, _05552_);
  and (_03522_, _03371_, _03369_);
  and (_03372_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_03373_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_03374_, _03373_, _03372_);
  and (_03375_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_03376_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03377_, _03376_, _03375_);
  or (_03378_, _03377_, _03374_);
  and (_03379_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03380_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_03381_, _03380_, _03379_);
  and (_03382_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03383_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_03384_, _03383_, _03382_);
  or (_03385_, _03384_, _03381_);
  or (_03386_, _03385_, _03378_);
  nor (_03387_, _13528_, _00760_);
  and (_03388_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_03389_, _03388_, _03387_);
  and (_03390_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_03391_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_03392_, _03391_, _03390_);
  or (_03393_, _03392_, _03389_);
  and (_03394_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_03395_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_03396_, _03395_, _03394_);
  and (_03397_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_03399_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_03400_, _03399_, _03397_);
  or (_03401_, _03400_, _03396_);
  or (_03402_, _03401_, _03393_);
  or (_03403_, _03402_, _03386_);
  and (_03404_, _13555_, _11345_);
  and (_03405_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_03406_, _03405_, _03404_);
  and (_03407_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_03408_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_03409_, _03408_, _03407_);
  or (_03410_, _03409_, _03406_);
  or (_03411_, _13592_, p0_in[6]);
  or (_03412_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03413_, _03412_, _03411_);
  and (_03414_, _03413_, _13574_);
  or (_03416_, _13592_, p1_in[6]);
  or (_03417_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03418_, _03417_, _03416_);
  and (_03419_, _03418_, _13598_);
  or (_03420_, _03419_, _03414_);
  or (_03421_, _13592_, p3_in[6]);
  or (_03422_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03423_, _03422_, _03421_);
  and (_03425_, _03423_, _13605_);
  or (_03426_, _13592_, p2_in[6]);
  or (_03427_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03429_, _03427_, _03426_);
  and (_03430_, _03429_, _13611_);
  or (_03431_, _03430_, _03425_);
  or (_03432_, _03431_, _03420_);
  or (_03434_, _03432_, _03410_);
  and (_03435_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_03437_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03438_, _03437_, _03435_);
  or (_03440_, _03438_, _03434_);
  or (_03442_, _03440_, _03403_);
  and (_03443_, _03442_, _13701_);
  and (_03444_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_03445_, _03444_, _13476_);
  or (_03447_, _03445_, _03443_);
  or (_03448_, _13704_, _07574_);
  and (_03449_, _03448_, _05552_);
  and (_03526_, _03449_, _03447_);
  and (_03450_, _05894_, _10917_);
  or (_03451_, _13578_, _10937_);
  or (_03452_, _03451_, _03450_);
  or (_03453_, _03452_, _10901_);
  or (_03455_, _03453_, _10934_);
  or (_03456_, _11149_, _10913_);
  or (_03457_, _03456_, _10941_);
  or (_03458_, _11115_, _11088_);
  or (_03459_, _03458_, _03457_);
  or (_03460_, _11022_, _10943_);
  or (_03461_, _11178_, _11015_);
  or (_03462_, _03461_, _03460_);
  and (_03463_, _12283_, _05837_);
  or (_03464_, _03463_, _13575_);
  or (_03465_, _03464_, _10929_);
  or (_03466_, _03465_, _10908_);
  or (_03468_, _03466_, _03462_);
  or (_03469_, _03468_, _03459_);
  or (_03470_, _03469_, _03455_);
  and (_03471_, _03470_, _05547_);
  and (_03472_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03473_, _03472_, _10956_);
  or (_03474_, _03473_, _03471_);
  and (_03548_, _03474_, _05552_);
  or (_03475_, _12332_, _12329_);
  or (_03476_, _10933_, _05842_);
  or (_03477_, _03476_, _13392_);
  or (_03478_, _03477_, _03475_);
  or (_03479_, _10851_, _05878_);
  and (_03480_, _10929_, _05737_);
  or (_03481_, _03480_, _12271_);
  or (_03482_, _03481_, _03479_);
  or (_03483_, _12308_, _05845_);
  nor (_03484_, _03483_, _11022_);
  nand (_03485_, _03484_, _12315_);
  or (_03486_, _03485_, _03482_);
  or (_03487_, _03486_, _12325_);
  or (_03488_, _03487_, _03478_);
  and (_03489_, _03488_, _05547_);
  and (_03490_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03491_, _03490_, _10958_);
  or (_03492_, _03491_, _03489_);
  and (_03558_, _03492_, _05552_);
  nor (_03494_, _09030_, _08386_);
  and (_03496_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_03497_, _03496_, _03494_);
  and (_03566_, _03497_, _05552_);
  or (_03498_, _01751_, _07483_);
  not (_03499_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_03500_, _01751_, _03499_);
  and (_03501_, _03500_, _06524_);
  and (_03502_, _03501_, _03498_);
  nor (_03503_, _06774_, _03499_);
  and (_03504_, _01750_, _10632_);
  nand (_03505_, _03504_, _06763_);
  or (_03506_, _03504_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_03507_, _03506_, _06775_);
  and (_03508_, _03507_, _03505_);
  or (_03509_, _03508_, _03503_);
  or (_03510_, _03509_, _03502_);
  and (_03593_, _03510_, _05552_);
  or (_03511_, _05689_, _08675_);
  or (_03512_, _05546_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_03513_, _03512_, _05552_);
  and (_03600_, _03513_, _03511_);
  or (_03514_, _01751_, _07711_);
  not (_03515_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_03516_, _01751_, _03515_);
  and (_03517_, _03516_, _06524_);
  and (_03518_, _03517_, _03514_);
  nor (_03519_, _06774_, _03515_);
  or (_03520_, _01751_, _08048_);
  and (_03521_, _03516_, _06775_);
  and (_03523_, _03521_, _03520_);
  or (_03524_, _03523_, _03519_);
  or (_03525_, _03524_, _03518_);
  and (_03603_, _03525_, _05552_);
  or (_03527_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_03528_, _06315_, rst);
  and (_03614_, _03528_, _03527_);
  and (_03529_, _02973_, _06771_);
  nand (_03530_, _03529_, _06763_);
  or (_03531_, _03529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03532_, _03531_, _06775_);
  and (_03533_, _03532_, _03530_);
  nand (_03534_, _02981_, _06811_);
  or (_03535_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03536_, _03535_, _06524_);
  and (_03537_, _03536_, _03534_);
  and (_03538_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_03539_, _03538_, rst);
  or (_03540_, _03539_, _03537_);
  or (_03623_, _03540_, _03533_);
  and (_03541_, _07951_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_03542_, _08386_, _07951_);
  or (_03543_, _03542_, _03541_);
  and (_03636_, _03543_, _05552_);
  or (_03544_, _01751_, _07574_);
  not (_03545_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_03546_, _01751_, _03545_);
  and (_03547_, _03546_, _06524_);
  and (_03549_, _03547_, _03544_);
  nor (_03550_, _06774_, _03545_);
  and (_03551_, _01750_, _08365_);
  nand (_03552_, _03551_, _06763_);
  or (_03553_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03554_, _03553_, _06775_);
  and (_03555_, _03554_, _03552_);
  or (_03556_, _03555_, _03550_);
  or (_03557_, _03556_, _03549_);
  and (_03638_, _03557_, _05552_);
  and (_03651_, _11308_, _05552_);
  and (_03559_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _07768_);
  and (_03560_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_03561_, _03560_, _03559_);
  and (_03660_, _03561_, _05552_);
  and (_03562_, _07635_, _05552_);
  or (_03563_, _03562_, _13477_);
  and (_03564_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_03565_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_03567_, _03565_, _03564_);
  and (_03568_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_03569_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_03570_, _03569_, _03568_);
  or (_03571_, _03570_, _03567_);
  and (_03572_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_03573_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or (_03574_, _03573_, _03572_);
  and (_03575_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_03576_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_03577_, _03576_, _03575_);
  or (_03578_, _03577_, _03574_);
  or (_03579_, _03578_, _03571_);
  nor (_03580_, _13528_, _00749_);
  and (_03581_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_03582_, _03581_, _03580_);
  and (_03583_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_03584_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_03585_, _03584_, _03583_);
  or (_03586_, _03585_, _03582_);
  and (_03587_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_03588_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_03589_, _03588_, _03587_);
  and (_03590_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_03591_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_03592_, _03591_, _03590_);
  or (_03594_, _03592_, _03589_);
  or (_03595_, _03594_, _03586_);
  or (_03596_, _03595_, _03579_);
  and (_03597_, _13555_, _11430_);
  and (_03598_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_03599_, _03598_, _03597_);
  and (_03601_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_03602_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_03604_, _03602_, _03601_);
  or (_03605_, _03604_, _03599_);
  or (_03606_, _13592_, p0_in[5]);
  or (_03607_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03608_, _03607_, _03606_);
  and (_03609_, _03608_, _13574_);
  or (_03610_, _13592_, p1_in[5]);
  or (_03611_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03612_, _03611_, _03610_);
  and (_03613_, _03612_, _13598_);
  or (_03615_, _03613_, _03609_);
  or (_03616_, _13592_, p2_in[5]);
  or (_03617_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03618_, _03617_, _03616_);
  and (_03619_, _03618_, _13611_);
  or (_03620_, _13592_, p3_in[5]);
  or (_03621_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03622_, _03621_, _03620_);
  and (_03624_, _03622_, _13605_);
  or (_03625_, _03624_, _03619_);
  or (_03626_, _03625_, _03615_);
  or (_03627_, _03626_, _03605_);
  and (_03628_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03629_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_03630_, _03629_, _03628_);
  or (_03631_, _03630_, _03627_);
  or (_03632_, _03631_, _03596_);
  and (_03633_, _03632_, _13701_);
  and (_03634_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_03635_, _03634_, _13476_);
  or (_03637_, _03635_, _03633_);
  and (_03665_, _03637_, _03563_);
  and (_03639_, _12299_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_03640_, _10945_, _10905_);
  or (_03641_, _11088_, _05816_);
  or (_03642_, _03641_, _03476_);
  or (_03643_, _03642_, _03640_);
  or (_03644_, _12331_, _12309_);
  or (_03646_, _05830_, _05824_);
  and (_03647_, _03646_, _10843_);
  or (_03648_, _03647_, _13383_);
  or (_03649_, _03648_, _03644_);
  or (_03650_, _11020_, _05841_);
  or (_03652_, _03650_, _05848_);
  or (_03653_, _03652_, _03649_);
  or (_03654_, _03653_, _03643_);
  or (_03655_, _03654_, _13400_);
  and (_03656_, _03655_, _06576_);
  or (_03671_, _03656_, _03639_);
  nand (_03657_, _08041_, _06949_);
  or (_03658_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_03659_, _03658_, _05552_);
  and (_03673_, _03659_, _03657_);
  nand (_03675_, _11626_, _05552_);
  and (_03661_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _07768_);
  and (_03662_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_03663_, _03662_, _03661_);
  and (_03679_, _03663_, _05552_);
  nand (_03664_, _00647_, _08996_);
  or (_03666_, _03664_, _00613_);
  nor (_03667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _08998_);
  nand (_03668_, _03667_, _00580_);
  and (_03669_, _03668_, _05552_);
  and (_03681_, _03669_, _03666_);
  or (_03670_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  nand (_03672_, _05550_, _11057_);
  and (_03674_, _03672_, _05552_);
  and (_03688_, _03674_, _03670_);
  nor (_03705_, _11900_, rst);
  and (_03676_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07768_);
  and (_03677_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_03678_, _03677_, _03676_);
  and (_03712_, _03678_, _05552_);
  nand (_03680_, _00241_, _07945_);
  or (_03682_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_03683_, _03682_, _05552_);
  and (_03714_, _03683_, _03680_);
  nand (_03684_, _00241_, _08386_);
  or (_03685_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_03686_, _03685_, _05552_);
  and (_03718_, _03686_, _03684_);
  nor (_03687_, _08041_, _06953_);
  and (_03689_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03690_, _03689_, _06955_);
  or (_03691_, _03690_, _03687_);
  or (_03692_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03693_, _03692_, _05552_);
  and (_03720_, _03693_, _03691_);
  nor (_03750_, _11672_, rst);
  and (_03694_, _03005_, _06771_);
  nand (_03695_, _03694_, _06763_);
  or (_03696_, _03694_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03697_, _03696_, _06775_);
  and (_03698_, _03697_, _03695_);
  nor (_03699_, _03011_, _06811_);
  and (_03700_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_03701_, _03700_, _03699_);
  and (_03702_, _03701_, _06524_);
  and (_03703_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_03704_, _03703_, rst);
  or (_03706_, _03704_, _03702_);
  or (_03760_, _03706_, _03698_);
  and (_03707_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_03708_, _07951_, _06560_);
  and (_03709_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03710_, _03709_, _01625_);
  or (_03711_, _03710_, _03708_);
  or (_03713_, _03711_, _03707_);
  and (_03769_, _03713_, _05552_);
  and (_03715_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07768_);
  and (_03716_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_03717_, _03716_, _03715_);
  and (_03771_, _03717_, _05552_);
  or (_03719_, _10982_, _08102_);
  or (_03721_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_03722_, _03721_, _05552_);
  and (_03775_, _03722_, _03719_);
  and (_03723_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_03724_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or (_03725_, _03724_, _03723_);
  and (_03784_, _03725_, _05552_);
  or (_03726_, _10982_, _07711_);
  or (_03727_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_03728_, _03727_, _05552_);
  and (_03814_, _03728_, _03726_);
  and (_03729_, _12299_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nand (_03730_, _06568_, _05738_);
  nor (_03731_, _05854_, _05840_);
  nand (_03732_, _03731_, _10906_);
  nand (_03733_, _03732_, _05894_);
  and (_03734_, _03733_, _11166_);
  and (_03735_, _03734_, _03730_);
  nand (_03736_, _05861_, _05818_);
  or (_03737_, _13583_, _10851_);
  and (_03738_, _05855_, _05818_);
  nor (_03739_, _03738_, _03737_);
  and (_03740_, _03739_, _03736_);
  nand (_03741_, _10929_, _05738_);
  or (_03743_, _13575_, _12284_);
  nor (_03744_, _03743_, _10924_);
  and (_03745_, _03744_, _03741_);
  nor (_03746_, _03456_, _12307_);
  and (_03747_, _03746_, _03745_);
  and (_03748_, _03747_, _03740_);
  nand (_03749_, _03748_, _03735_);
  and (_03751_, _03749_, _06576_);
  or (_03824_, _03751_, _03729_);
  nand (_03752_, _00241_, _06306_);
  or (_03753_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_03754_, _03753_, _05552_);
  and (_03844_, _03754_, _03752_);
  and (_03846_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_03755_, _07951_, _06811_);
  and (_03756_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_03757_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_03758_, _03757_, _01625_);
  or (_03759_, _03758_, _03756_);
  or (_03761_, _03759_, _03755_);
  and (_03850_, _03761_, _05552_);
  or (_03762_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_03763_, _05550_, _05748_);
  and (_03764_, _03763_, _05552_);
  and (_03873_, _03764_, _03762_);
  and (_03765_, _08874_, rxd_i);
  not (_03766_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nor (_03767_, _08874_, _03766_);
  or (_03768_, _03767_, _03765_);
  and (_03881_, _03768_, _05552_);
  and (_03883_, _07209_, _05552_);
  and (_03770_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_03772_, _07939_, _06811_);
  or (_03773_, _03772_, _03770_);
  and (_03888_, _03773_, _05552_);
  or (_03774_, _01751_, _07255_);
  not (_03776_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_03777_, _01751_, _03776_);
  and (_03778_, _03777_, _06524_);
  and (_03779_, _03778_, _03774_);
  nor (_03780_, _06774_, _03776_);
  and (_03781_, _01750_, _06771_);
  nand (_03782_, _03781_, _06763_);
  or (_03783_, _03781_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03785_, _03783_, _06775_);
  and (_03786_, _03785_, _03782_);
  or (_03787_, _03786_, _03780_);
  or (_03788_, _03787_, _03779_);
  and (_03895_, _03788_, _05552_);
  and (_03789_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_03790_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_03791_, _03790_, _03789_);
  and (_03902_, _03791_, _05552_);
  and (_03792_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_03793_, _03792_, _13739_);
  and (_03794_, _07946_, _06309_);
  and (_03795_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_03796_, _03795_, _03794_);
  or (_03797_, _03796_, _03793_);
  and (_03914_, _03797_, _05552_);
  or (_03798_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand (_03799_, _05550_, _05699_);
  and (_03800_, _03799_, _05552_);
  and (_03936_, _03800_, _03798_);
  not (_03801_, _01819_);
  not (_03802_, _10639_);
  and (_03803_, _01824_, _03802_);
  and (_03804_, _03803_, _01803_);
  nand (_03805_, _03804_, _03801_);
  or (_03806_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_03807_, _03806_, _05552_);
  and (_03966_, _03807_, _03805_);
  not (_03808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_03809_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_03810_, _03809_, _05560_);
  and (_03811_, _03810_, _00384_);
  or (_03812_, _03811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_03813_, _03812_, _00225_);
  or (_03815_, _06060_, _05570_);
  nand (_03816_, _03815_, _00225_);
  or (_03817_, _03816_, _13359_);
  and (_03818_, _03817_, _03813_);
  or (_03819_, _03818_, _00232_);
  nand (_03820_, _00232_, _07945_);
  and (_03821_, _03820_, _05552_);
  and (_03974_, _03821_, _03819_);
  or (_03822_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_03823_, _05550_, _11002_);
  and (_03825_, _03823_, _05552_);
  and (_04015_, _03825_, _03822_);
  or (_03826_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_03827_, _05550_, _07743_);
  and (_03828_, _03827_, _05552_);
  and (_04017_, _03828_, _03826_);
  and (_03829_, _00225_, _08365_);
  nand (_03830_, _03829_, _06763_);
  or (_03831_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03832_, _03831_, _00451_);
  and (_03833_, _03832_, _03830_);
  nor (_03834_, _00451_, _08386_);
  or (_03835_, _03834_, _03833_);
  and (_04020_, _03835_, _05552_);
  or (_03836_, _13701_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_03837_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03838_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_03839_, _03838_, _03837_);
  and (_03840_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_03841_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_03842_, _03841_, _03840_);
  or (_03843_, _03842_, _03839_);
  and (_03845_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03847_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_03848_, _03847_, _03845_);
  and (_03849_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03851_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03852_, _03851_, _03849_);
  or (_03853_, _03852_, _03848_);
  or (_03854_, _03853_, _03843_);
  and (_03855_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_03856_, _13528_, _00758_);
  or (_03857_, _03856_, _03855_);
  and (_03858_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_03859_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_03860_, _03859_, _03858_);
  or (_03861_, _03860_, _03857_);
  and (_03862_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03863_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03864_, _03863_, _03862_);
  and (_03865_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03866_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03867_, _03866_, _03865_);
  or (_03868_, _03867_, _03864_);
  or (_03869_, _03868_, _03861_);
  or (_03870_, _03869_, _03854_);
  and (_03871_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_03872_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_03874_, _03872_, _03871_);
  and (_03875_, _13555_, _11308_);
  and (_03876_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_03877_, _03876_, _03875_);
  or (_03878_, _03877_, _03874_);
  or (_03879_, _13592_, p3_in[7]);
  or (_03880_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03882_, _03880_, _03879_);
  and (_03884_, _03882_, _13605_);
  or (_03885_, _13592_, p2_in[7]);
  or (_03886_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03887_, _03886_, _03885_);
  and (_03889_, _03887_, _13611_);
  or (_03890_, _03889_, _03884_);
  or (_03891_, _13592_, p1_in[7]);
  or (_03892_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03893_, _03892_, _03891_);
  and (_03894_, _03893_, _13598_);
  or (_03896_, _13592_, p0_in[7]);
  or (_03897_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03898_, _03897_, _03896_);
  and (_03899_, _03898_, _13574_);
  or (_03900_, _03899_, _03894_);
  or (_03901_, _03900_, _03890_);
  or (_03903_, _03901_, _03878_);
  and (_03904_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_03905_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03906_, _03905_, _03904_);
  or (_03907_, _03906_, _03903_);
  or (_03908_, _03907_, _03870_);
  and (_03909_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_03910_, _03909_, _03908_);
  and (_03911_, _03910_, _03836_);
  or (_03912_, _03911_, _13476_);
  or (_03913_, _13704_, _07255_);
  and (_03915_, _03913_, _05552_);
  and (_04036_, _03915_, _03912_);
  nor (_03916_, _00374_, rst);
  or (_03917_, _00373_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand (_03918_, _00373_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03919_, _03918_, _03917_);
  and (_04039_, _03919_, _03916_);
  or (_03920_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_03921_, _05550_, _05677_);
  and (_03922_, _03921_, _05552_);
  and (_04044_, _03922_, _03920_);
  and (_04050_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_03923_, _07951_, _06306_);
  and (_03924_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_03925_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_03926_, _03925_, _01625_);
  or (_03927_, _03926_, _03924_);
  or (_03928_, _03927_, _03923_);
  and (_04052_, _03928_, _05552_);
  and (_04054_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_03929_, _12308_, _10851_);
  or (_03930_, _12280_, _10913_);
  or (_03931_, _03930_, _03929_);
  or (_03932_, _03931_, _11088_);
  and (_03933_, _03932_, _05547_);
  and (_03934_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03935_, _03934_, _05901_);
  or (_03937_, _03935_, _03933_);
  and (_04062_, _03937_, _05552_);
  and (_03938_, _01740_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03939_, _03938_, _01741_);
  and (_03940_, _03939_, _08009_);
  nand (_03941_, _11591_, _06763_);
  nor (_03942_, _11591_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_03943_, _03942_, _08009_);
  and (_03944_, _03943_, _03941_);
  or (_03945_, _03944_, _06531_);
  or (_03946_, _03945_, _03940_);
  nand (_03947_, _06811_, _06531_);
  and (_03948_, _03947_, _05552_);
  and (_04069_, _03948_, _03946_);
  and (_04074_, _07117_, _05552_);
  and (_03949_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_03950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _08998_);
  nor (_03951_, _03950_, _03667_);
  nor (_03952_, _03951_, _00857_);
  or (_03953_, _03952_, _00580_);
  or (_03954_, _03953_, _03949_);
  or (_03955_, _03951_, _00838_);
  and (_03956_, _03955_, _05552_);
  and (_04077_, _03956_, _03954_);
  nor (_04080_, _11095_, rst);
  or (_03957_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_03958_, _05550_, _05611_);
  and (_03959_, _03958_, _05552_);
  and (_04082_, _03959_, _03957_);
  and (_03960_, _12299_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_03961_, _06567_, _05857_);
  or (_03962_, _03961_, _05831_);
  or (_03963_, _03962_, _11133_);
  or (_03964_, _11570_, _11124_);
  and (_03965_, _06570_, _05894_);
  or (_03967_, _13386_, _03965_);
  or (_03968_, _03967_, _03964_);
  or (_03969_, _11127_, _11167_);
  or (_03970_, _03969_, _11573_);
  or (_03971_, _03970_, _03968_);
  or (_03972_, _03971_, _03963_);
  and (_03973_, _03972_, _06576_);
  or (_04091_, _03973_, _03960_);
  and (_04128_, _07200_, _05552_);
  and (_04133_, _00375_, _05552_);
  or (_04142_, _08764_, _06568_);
  and (_03975_, _05803_, _07781_);
  and (_03976_, _03975_, _05781_);
  or (_03977_, _07897_, _07775_);
  and (_03978_, _03977_, _03976_);
  and (_03979_, _07898_, _07807_);
  or (_03980_, _03979_, _02640_);
  or (_03981_, _03980_, _03978_);
  or (_03982_, _07853_, _07840_);
  and (_03983_, _07862_, _05710_);
  or (_03984_, _07923_, _03983_);
  or (_03985_, _03984_, _03982_);
  nand (_03986_, _07848_, _07815_);
  nor (_03987_, _07798_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_03988_, _03987_, _03986_);
  nand (_03989_, _03988_, _07786_);
  nand (_03990_, _07867_, _07864_);
  or (_03991_, _03990_, _03989_);
  or (_03992_, _03991_, _03985_);
  or (_03993_, _03992_, _03981_);
  or (_03994_, _03993_, _02649_);
  and (_03995_, _03994_, _05608_);
  nor (_03996_, _02639_, _05891_);
  or (_03997_, _03996_, rst);
  or (_04144_, _03997_, _03995_);
  and (_04147_, _13702_, _13477_);
  and (_03998_, _13621_, _11279_);
  or (_03999_, _13677_, _13481_);
  or (_04000_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_04001_, _04000_, _13480_);
  and (_04002_, _04001_, _03999_);
  and (_04003_, _13509_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_04004_, _13497_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_04005_, _04004_, _04003_);
  and (_04006_, _04005_, _13481_);
  and (_04007_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_04008_, _11763_, _07468_);
  or (_04009_, _04008_, _04007_);
  and (_04010_, _04009_, _13464_);
  and (_04011_, _13509_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_04012_, _13497_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_04013_, _04012_, _04011_);
  and (_04014_, _04013_, _11763_);
  or (_04016_, _04014_, _04010_);
  or (_04018_, _04016_, _04006_);
  or (_04019_, _04018_, _04002_);
  and (_04021_, _04019_, _03998_);
  not (_04022_, _11279_);
  and (_04023_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_04024_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_04025_, _04024_, _04023_);
  and (_04026_, _04025_, _13509_);
  and (_04027_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_04028_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_04029_, _04028_, _04027_);
  and (_04030_, _04029_, _13464_);
  nor (_04031_, _11763_, _00592_);
  and (_04032_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_04033_, _04032_, _04031_);
  and (_04034_, _04033_, _13480_);
  or (_04035_, _04034_, _04030_);
  nor (_04037_, _11763_, _00587_);
  and (_04038_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_04040_, _04038_, _04037_);
  and (_04041_, _04040_, _13497_);
  or (_04042_, _04041_, _04035_);
  or (_04043_, _04042_, _04026_);
  and (_04045_, _04043_, _13515_);
  and (_04046_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_04047_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_04048_, _04047_, _04046_);
  and (_04049_, _04048_, _13509_);
  and (_04051_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_04053_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_04055_, _04053_, _04051_);
  and (_04056_, _04055_, _13464_);
  nor (_04057_, _11763_, _01054_);
  and (_04058_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_04059_, _04058_, _04057_);
  and (_04060_, _04059_, _13480_);
  or (_04061_, _04060_, _04056_);
  and (_04063_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_04064_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_04065_, _04064_, _04063_);
  and (_04066_, _04065_, _13497_);
  or (_04067_, _04066_, _04061_);
  or (_04068_, _04067_, _04049_);
  and (_04070_, _04068_, _13472_);
  or (_04071_, _04070_, _04045_);
  and (_04072_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04073_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_04075_, _04073_, _04072_);
  and (_04076_, _04075_, _13464_);
  nor (_04078_, _11763_, _02787_);
  and (_04079_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_04081_, _04079_, _04078_);
  and (_04083_, _04081_, _13480_);
  or (_04084_, _04083_, _04076_);
  and (_04085_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_04086_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_04087_, _04086_, _04085_);
  and (_04088_, _04087_, _13509_);
  nor (_04089_, _11763_, _12096_);
  and (_04090_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_04092_, _04090_, _04089_);
  and (_04093_, _04092_, _13497_);
  or (_04094_, _04093_, _04088_);
  or (_04095_, _04094_, _04084_);
  and (_04096_, _04095_, _13487_);
  or (_04097_, _04096_, _04071_);
  and (_04098_, _04097_, _04022_);
  and (_04099_, _13620_, _11279_);
  and (_04100_, _04099_, _13560_);
  nor (_04101_, _04100_, _03998_);
  and (_04102_, _11509_, _11279_);
  and (_04103_, _13561_, _04102_);
  nor (_04104_, _13469_, _04022_);
  nor (_04105_, _04104_, _04103_);
  and (_04106_, _04105_, _04101_);
  nor (_04107_, _13487_, _13727_);
  or (_04108_, _04107_, _11279_);
  nand (_04109_, _13514_, _11279_);
  and (_04110_, _04109_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_04111_, _04110_, _04108_);
  and (_04112_, _04111_, _04106_);
  nor (_04113_, _13471_, _04022_);
  and (_04114_, _00114_, _11763_);
  and (_04115_, _03413_, _13481_);
  or (_04116_, _04115_, _04114_);
  and (_04117_, _04116_, _13464_);
  and (_04118_, _13812_, _13481_);
  and (_04119_, _13596_, _11763_);
  or (_04120_, _04119_, _04118_);
  and (_04121_, _04120_, _13480_);
  or (_04122_, _04121_, _04117_);
  and (_04123_, _00184_, _11763_);
  and (_04124_, _03608_, _13481_);
  or (_04125_, _04124_, _04123_);
  and (_04126_, _04125_, _13497_);
  and (_04127_, _03898_, _13481_);
  and (_04129_, _00023_, _11763_);
  or (_04130_, _04129_, _04127_);
  and (_04131_, _04130_, _13509_);
  or (_04132_, _04131_, _04126_);
  or (_04134_, _04132_, _04122_);
  and (_04135_, _04134_, _04113_);
  or (_04136_, _04135_, _04112_);
  and (_04137_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor (_04138_, _11763_, _03545_);
  or (_04139_, _04138_, _04137_);
  and (_04140_, _04139_, _13464_);
  nor (_04141_, _11763_, _01767_);
  and (_04143_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_04145_, _04143_, _04141_);
  and (_04146_, _04145_, _13480_);
  or (_04148_, _04146_, _04140_);
  and (_04149_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_04150_, _11763_, _03776_);
  or (_04151_, _04150_, _04149_);
  and (_04152_, _04151_, _13509_);
  nor (_04153_, _11763_, _01753_);
  and (_04155_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_04156_, _04155_, _04153_);
  and (_04157_, _04156_, _13497_);
  or (_04158_, _04157_, _04152_);
  or (_04159_, _04158_, _04148_);
  and (_04160_, _04159_, _04100_);
  and (_04161_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_04162_, _11763_, _06396_);
  or (_04163_, _04162_, _04161_);
  and (_04164_, _04163_, _13464_);
  nor (_04165_, _11763_, _06157_);
  and (_04167_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_04169_, _04167_, _04165_);
  and (_04170_, _04169_, _13480_);
  or (_04171_, _04170_, _04164_);
  and (_04172_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_04173_, _11763_, _06361_);
  or (_04174_, _04173_, _04172_);
  and (_04175_, _04174_, _13509_);
  nor (_04177_, _11763_, _06103_);
  and (_04178_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_04180_, _04178_, _04177_);
  and (_04182_, _04180_, _13497_);
  or (_04183_, _04182_, _04175_);
  or (_04185_, _04183_, _04171_);
  and (_04187_, _04185_, _04103_);
  or (_04189_, _04187_, _04160_);
  or (_04190_, _04189_, _04136_);
  nor (_04191_, _11763_, _03808_);
  and (_04192_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_04193_, _04192_, _04191_);
  and (_04194_, _04193_, _13497_);
  or (_04195_, _04194_, _11279_);
  and (_04196_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_04197_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04198_, _04197_, _04196_);
  and (_04199_, _04198_, _13464_);
  and (_04200_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_04201_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_04202_, _04201_, _04200_);
  and (_04203_, _04202_, _13480_);
  and (_04204_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_04205_, _11763_, _12098_);
  or (_04206_, _04205_, _04204_);
  and (_04207_, _04206_, _13509_);
  or (_04208_, _04207_, _04203_);
  or (_04209_, _04208_, _04199_);
  or (_04210_, _04209_, _04195_);
  and (_04211_, _13602_, _11763_);
  and (_04212_, _13817_, _13481_);
  or (_04213_, _04212_, _04211_);
  and (_04214_, _04213_, _13480_);
  and (_04215_, _00188_, _11763_);
  and (_04216_, _03612_, _13481_);
  or (_04217_, _04216_, _04215_);
  and (_04218_, _04217_, _13497_);
  or (_04219_, _04218_, _04022_);
  or (_04220_, _04219_, _04214_);
  and (_04222_, _00110_, _13464_);
  and (_04223_, _00029_, _13509_);
  or (_04224_, _04223_, _04222_);
  and (_04225_, _04224_, _11763_);
  and (_04226_, _03418_, _13464_);
  and (_04227_, _03893_, _13509_);
  or (_04228_, _04227_, _04226_);
  and (_04229_, _04228_, _13481_);
  or (_04230_, _04229_, _04225_);
  or (_04231_, _04230_, _04220_);
  and (_04232_, _04231_, _13540_);
  and (_04233_, _04232_, _04210_);
  and (_04234_, _13615_, _11763_);
  and (_04235_, _13801_, _13481_);
  or (_04236_, _04235_, _04234_);
  and (_04237_, _04236_, _13480_);
  and (_04238_, _00175_, _11763_);
  and (_04239_, _03618_, _13481_);
  or (_04240_, _04239_, _04238_);
  and (_04241_, _04240_, _13497_);
  or (_04242_, _04241_, _13465_);
  or (_04243_, _04242_, _04237_);
  and (_04244_, _00105_, _13464_);
  and (_04245_, _00040_, _13509_);
  or (_04246_, _04245_, _04244_);
  and (_04247_, _04246_, _11763_);
  and (_04248_, _03429_, _13464_);
  and (_04249_, _03887_, _13509_);
  or (_04250_, _04249_, _04248_);
  and (_04251_, _04250_, _13481_);
  or (_04252_, _04251_, _04247_);
  or (_04253_, _04252_, _04243_);
  and (_04254_, _13609_, _11763_);
  and (_04255_, _13806_, _13481_);
  or (_04256_, _04255_, _04254_);
  and (_04257_, _04256_, _13480_);
  and (_04258_, _00179_, _11763_);
  and (_04259_, _03622_, _13481_);
  or (_04260_, _04259_, _04258_);
  and (_04261_, _04260_, _13497_);
  or (_04262_, _04261_, _11509_);
  nor (_04263_, _04262_, _04257_);
  nand (_04264_, _00101_, _13464_);
  nand (_04265_, _00035_, _13509_);
  and (_04266_, _04265_, _04264_);
  or (_04267_, _04266_, _13481_);
  nand (_04268_, _03423_, _13464_);
  nand (_04269_, _03882_, _13509_);
  and (_04270_, _04269_, _04268_);
  or (_04271_, _04270_, _11763_);
  and (_04272_, _04271_, _04267_);
  and (_04273_, _04272_, _04263_);
  nor (_04274_, _04273_, _04109_);
  and (_04276_, _04274_, _04253_);
  and (_04277_, _13518_, _04022_);
  nor (_04278_, _11763_, _00617_);
  and (_04279_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_04280_, _04279_, _04278_);
  and (_04281_, _04280_, _13480_);
  nor (_04282_, _11763_, _00615_);
  and (_04283_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_04285_, _04283_, _04282_);
  and (_04286_, _04285_, _13497_);
  or (_04287_, _04286_, _04281_);
  and (_04288_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_04289_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_04290_, _04289_, _04288_);
  and (_04291_, _04290_, _13464_);
  and (_04292_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_04293_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_04294_, _04293_, _04292_);
  and (_04296_, _04294_, _13509_);
  or (_04297_, _04296_, _04291_);
  or (_04298_, _04297_, _04287_);
  and (_04299_, _04298_, _04277_);
  and (_04300_, _11769_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or (_04301_, _04300_, _04299_);
  or (_04302_, _04301_, _04276_);
  or (_04303_, _04302_, _04233_);
  or (_04304_, _04303_, _04190_);
  or (_04305_, _04304_, _04098_);
  or (_04306_, _04305_, _04021_);
  and (_04307_, _04103_, _06965_);
  nor (_04308_, _04307_, _11518_);
  nand (_04309_, _04300_, _06763_);
  and (_04310_, _04309_, _04308_);
  and (_04311_, _04310_, _04306_);
  and (_04312_, _11763_, _11214_);
  nor (_04313_, _11763_, _06811_);
  or (_04314_, _04313_, _04312_);
  and (_04315_, _04314_, _13509_);
  nor (_04316_, _11763_, _07388_);
  and (_04317_, _11763_, _11238_);
  or (_04318_, _04317_, _04316_);
  and (_04319_, _04318_, _13480_);
  nor (_04320_, _11763_, _08386_);
  and (_04321_, _11763_, _11726_);
  or (_04322_, _04321_, _04320_);
  and (_04323_, _04322_, _13464_);
  or (_04324_, _04323_, _04319_);
  nor (_04325_, _11763_, _06306_);
  and (_04326_, _11763_, _11234_);
  or (_04327_, _04326_, _04325_);
  and (_04328_, _04327_, _13497_);
  or (_04329_, _04328_, _04324_);
  nor (_04330_, _04329_, _04315_);
  nor (_04331_, _04330_, _04308_);
  or (_04332_, _04331_, _04311_);
  and (_04154_, _04332_, _05552_);
  and (_04333_, _02681_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_04334_, _02680_, _11238_);
  or (_04335_, _04334_, _04333_);
  and (_04166_, _04335_, _05552_);
  or (_04336_, _05781_, _08675_);
  or (_04337_, _05546_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_04338_, _04337_, _05552_);
  and (_04168_, _04338_, _04336_);
  and (_04339_, _12299_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_04340_, _11559_, _10913_);
  nand (_04341_, _05894_, _05840_);
  nand (_04342_, _10923_, _04341_);
  or (_04343_, _04342_, _04340_);
  not (_04344_, _11088_);
  nand (_04345_, _11111_, _04344_);
  or (_04346_, _04345_, _04343_);
  or (_04347_, _04346_, _12332_);
  or (_04348_, _04347_, _12327_);
  and (_04349_, _04348_, _06576_);
  or (_04176_, _04349_, _04339_);
  and (_04350_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_04351_, _05858_, _05547_);
  or (_04353_, _04351_, _04350_);
  or (_04354_, _04353_, _05901_);
  and (_04179_, _04354_, _05552_);
  or (_04355_, _03961_, _05889_);
  or (_04356_, _05890_, _05547_);
  and (_04357_, _04356_, _04355_);
  and (_04358_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04359_, _04358_, _10956_);
  or (_04360_, _04359_, _04357_);
  and (_04181_, _04360_, _05552_);
  and (_04361_, _12299_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_04362_, _11174_, _05829_);
  or (_04363_, _03647_, _12331_);
  or (_04364_, _04363_, _04362_);
  or (_04365_, _12324_, _11167_);
  or (_04366_, _04365_, _03483_);
  or (_04367_, _04366_, _03641_);
  or (_04368_, _04367_, _04364_);
  and (_04369_, _04368_, _06576_);
  or (_04184_, _04369_, _04361_);
  and (_04370_, _12299_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_04371_, _03743_, _05855_);
  or (_04372_, _13578_, _10847_);
  or (_04373_, _04372_, _04371_);
  or (_04374_, _03737_, _10897_);
  or (_04375_, _04374_, _04373_);
  or (_04376_, _12270_, _11152_);
  or (_04377_, _04376_, _12334_);
  or (_04378_, _04377_, _04375_);
  or (_04379_, _04378_, _12327_);
  and (_04380_, _04379_, _06576_);
  or (_04186_, _04380_, _04370_);
  and (_04381_, _13384_, _05547_);
  nand (_04382_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_04383_, _04382_, _10959_);
  or (_04384_, _04383_, _04381_);
  and (_04188_, _04384_, _05552_);
  or (_04385_, _12308_, _11033_);
  or (_04386_, _04385_, _05876_);
  or (_04387_, _04386_, _11180_);
  or (_04388_, _03479_, _05873_);
  or (_04389_, _04388_, _04387_);
  or (_04390_, _12332_, _10849_);
  or (_04391_, _04390_, _04389_);
  or (_04392_, _04391_, _05868_);
  and (_04393_, _04392_, _05547_);
  and (_04394_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04395_, _04394_, _05903_);
  or (_04396_, _04395_, _04393_);
  and (_04221_, _04396_, _05552_);
  or (_04397_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_04398_, _05550_, _11383_);
  and (_04399_, _04398_, _05552_);
  and (_04275_, _04399_, _04397_);
  or (_04400_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand (_04401_, _05550_, _11441_);
  and (_04402_, _04401_, _05552_);
  and (_04284_, _04402_, _04400_);
  or (_04403_, _07668_, _07635_);
  or (_04404_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_04405_, _04404_, _05552_);
  and (_04295_, _04405_, _04403_);
  or (_04406_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand (_04407_, _05550_, _11061_);
  and (_04408_, _04407_, _05552_);
  and (_04352_, _04408_, _04406_);
  and (_04409_, _01515_, _06771_);
  nand (_04410_, _04409_, _06763_);
  or (_04411_, _04409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_04412_, _04411_, _01521_);
  and (_04413_, _04412_, _04410_);
  nor (_04415_, _01521_, _06811_);
  or (_04416_, _04415_, _04413_);
  and (_04414_, _04416_, _05552_);
  and (_04417_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_04418_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_04419_, pc_log_change, _04418_);
  or (_04420_, _04419_, _04417_);
  and (_04429_, _04420_, _05552_);
  not (_04421_, cy_reg);
  and (_04422_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04423_, _04422_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04424_, _04423_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04425_, _04423_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04426_, _04425_, _04424_);
  and (_04427_, _04426_, _08302_);
  nor (_04428_, _04422_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04430_, _04428_, _04423_);
  or (_04431_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_04432_, _04431_, _04422_);
  nand (_04433_, _04432_, _04430_);
  nor (_04434_, _04433_, _04427_);
  nor (_04435_, _04426_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand (_04436_, _04426_, _08796_);
  nand (_04437_, _04436_, _04423_);
  nor (_04438_, _04437_, _04435_);
  or (_04439_, _04438_, _04434_);
  and (_04440_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02500_);
  nand (_04441_, _04426_, _08298_);
  or (_04442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_04443_, _04442_, _04430_);
  and (_04444_, _04443_, _04441_);
  not (_04445_, _04430_);
  nor (_04446_, _04426_, _08424_);
  and (_04447_, _04426_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_04448_, _04447_, _04446_);
  and (_04449_, _04448_, _04445_);
  or (_04450_, _04449_, _04444_);
  and (_04451_, _04450_, _04440_);
  or (_04452_, _04451_, _04439_);
  nor (_04453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_04454_, _04426_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_04455_, _02512_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_04456_, _04455_, _04430_);
  and (_04457_, _04456_, _04454_);
  nor (_04458_, _04426_, _08276_);
  and (_04459_, _04426_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_04460_, _04459_, _04458_);
  and (_04461_, _04460_, _04445_);
  or (_04462_, _04461_, _04457_);
  and (_04463_, _04462_, _04453_);
  and (_04464_, _02505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_04465_, _04426_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_04466_, _02512_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_04467_, _04466_, _04430_);
  and (_04468_, _04467_, _04465_);
  nor (_04469_, _04426_, _08262_);
  and (_04470_, _04426_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_04471_, _04470_, _04469_);
  and (_04472_, _04471_, _04445_);
  or (_04473_, _04472_, _04468_);
  and (_04474_, _04473_, _04464_);
  or (_04475_, _04474_, _04463_);
  or (_04476_, _04475_, _04452_);
  and (_04477_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_04478_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or (_04479_, _04478_, _04477_);
  and (_04480_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04481_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  or (_04482_, _04481_, _04480_);
  or (_04483_, _04482_, _04479_);
  or (_04484_, _04483_, _04445_);
  not (_04485_, _04426_);
  and (_04486_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04487_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  or (_04488_, _04487_, _04486_);
  and (_04489_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_04491_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  or (_04492_, _04491_, _04489_);
  or (_04493_, _04492_, _04488_);
  or (_04494_, _04493_, _04430_);
  and (_04495_, _04494_, _04485_);
  and (_04496_, _04495_, _04484_);
  and (_04497_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04498_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  or (_04499_, _04498_, _04497_);
  and (_04500_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_04501_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  or (_04502_, _04501_, _04500_);
  or (_04503_, _04502_, _04499_);
  or (_04504_, _04503_, _04430_);
  and (_04505_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04506_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  or (_04507_, _04506_, _04505_);
  and (_04508_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_04509_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  or (_04510_, _04509_, _04508_);
  or (_04511_, _04510_, _04507_);
  or (_04512_, _04511_, _04445_);
  and (_04513_, _04512_, _04426_);
  and (_04514_, _04513_, _04504_);
  or (_04515_, _04514_, _04496_);
  and (_04516_, _04515_, _04476_);
  and (_04517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04518_, _04517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04519_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_04520_, _04519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_04521_, _04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_04522_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_04523_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_04524_, _04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_04525_, _04524_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_04526_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_04527_, _04526_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_04528_, _04527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_04529_, _04528_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04530_, _04528_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04531_, _04530_, _04529_);
  and (_04532_, _04531_, _04516_);
  nor (_04533_, _04526_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04534_, _04533_, _04527_);
  and (_04535_, _04534_, _04516_);
  and (_04536_, _04535_, _02061_);
  nor (_04537_, _04527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_04538_, _04537_, _04528_);
  and (_04539_, _04538_, _04516_);
  nor (_04540_, _04538_, _04516_);
  nor (_04541_, _04540_, _04539_);
  nor (_04542_, _04524_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_04543_, _04542_, _04525_);
  and (_04544_, _04543_, _04516_);
  and (_04545_, _04544_, _02523_);
  nor (_04546_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04547_, _04546_, _04526_);
  and (_04548_, _04547_, _04516_);
  nor (_04549_, _04547_, _04516_);
  nor (_04550_, _04549_, _04548_);
  nor (_04551_, _04543_, _04516_);
  nor (_04552_, _04551_, _04544_);
  not (_04553_, _04552_);
  nor (_04554_, _04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_04555_, _04554_, _04524_);
  and (_04556_, _04555_, _04516_);
  nor (_04557_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_04558_, _04557_, _04523_);
  and (_04559_, _04558_, _04516_);
  nor (_04560_, _04555_, _04516_);
  nor (_04561_, _04560_, _04556_);
  nor (_04562_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_04563_, _04562_, _04522_);
  and (_04564_, _04563_, _04516_);
  nor (_04565_, _04563_, _04516_);
  nor (_04566_, _04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_04567_, _04566_, _04521_);
  and (_04568_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_04569_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or (_04570_, _04569_, _04568_);
  and (_04572_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_04573_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or (_04574_, _04573_, _04572_);
  or (_04575_, _04574_, _04570_);
  or (_04576_, _04575_, _04430_);
  and (_04577_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_04578_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  or (_04579_, _04578_, _04577_);
  and (_04580_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04581_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or (_04582_, _04581_, _04580_);
  or (_04583_, _04582_, _04579_);
  or (_04584_, _04583_, _04445_);
  and (_04585_, _04584_, _04576_);
  or (_04586_, _04585_, _04485_);
  and (_04587_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_04588_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or (_04589_, _04588_, _04587_);
  and (_04590_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_04591_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or (_04592_, _04591_, _04590_);
  or (_04593_, _04592_, _04589_);
  or (_04594_, _04593_, _04430_);
  and (_04595_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04596_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or (_04597_, _04596_, _04595_);
  and (_04598_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04599_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or (_04600_, _04599_, _04598_);
  or (_04601_, _04600_, _04597_);
  or (_04602_, _04601_, _04445_);
  and (_04603_, _04602_, _04594_);
  or (_04604_, _04603_, _04426_);
  and (_04605_, _04604_, _04586_);
  and (_04606_, _04605_, _04476_);
  and (_04607_, _04606_, _04567_);
  nor (_04608_, _04606_, _04567_);
  nor (_04609_, _04608_, _04607_);
  not (_04610_, _04609_);
  and (_04611_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_04612_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  or (_04613_, _04612_, _04611_);
  and (_04614_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_04615_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or (_04616_, _04615_, _04614_);
  or (_04617_, _04616_, _04613_);
  or (_04618_, _04617_, _04445_);
  and (_04619_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_04620_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  or (_04621_, _04620_, _04619_);
  and (_04622_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_04623_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or (_04624_, _04623_, _04622_);
  or (_04625_, _04624_, _04621_);
  or (_04626_, _04625_, _04430_);
  and (_04627_, _04626_, _04485_);
  and (_04628_, _04627_, _04618_);
  and (_04629_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_04630_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  or (_04631_, _04630_, _04629_);
  and (_04632_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_04633_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  or (_04634_, _04633_, _04632_);
  or (_04635_, _04634_, _04631_);
  or (_04636_, _04635_, _04430_);
  and (_04637_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_04638_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  or (_04639_, _04638_, _04637_);
  and (_04640_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_04641_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  or (_04642_, _04641_, _04640_);
  or (_04643_, _04642_, _04639_);
  or (_04644_, _04643_, _04445_);
  and (_04645_, _04644_, _04426_);
  and (_04646_, _04645_, _04636_);
  or (_04647_, _04646_, _04628_);
  and (_04648_, _04647_, _04476_);
  nor (_04649_, _04519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_04650_, _04649_, _04520_);
  and (_04651_, _04650_, _04648_);
  nor (_04652_, _04650_, _04648_);
  nor (_04653_, _04652_, _04651_);
  not (_04654_, _04653_);
  nor (_04655_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_04656_, _04655_, _04519_);
  and (_04657_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_04658_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  or (_04659_, _04658_, _04657_);
  and (_04660_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_04661_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or (_04662_, _04661_, _04660_);
  or (_04663_, _04662_, _04659_);
  or (_04664_, _04663_, _04445_);
  and (_04665_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_04666_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  or (_04667_, _04666_, _04665_);
  and (_04668_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_04669_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or (_04670_, _04669_, _04668_);
  or (_04671_, _04670_, _04667_);
  or (_04672_, _04671_, _04430_);
  and (_04673_, _04672_, _04485_);
  and (_04674_, _04673_, _04664_);
  and (_04675_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04676_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or (_04677_, _04676_, _04675_);
  and (_04678_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_04679_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or (_04680_, _04679_, _04678_);
  or (_04681_, _04680_, _04677_);
  or (_04682_, _04681_, _04430_);
  and (_04683_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04684_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or (_04685_, _04684_, _04683_);
  and (_04686_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04687_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or (_04688_, _04687_, _04686_);
  or (_04689_, _04688_, _04685_);
  or (_04690_, _04689_, _04445_);
  and (_04691_, _04690_, _04426_);
  and (_04692_, _04691_, _04682_);
  or (_04693_, _04692_, _04674_);
  and (_04694_, _04693_, _04476_);
  and (_04695_, _04694_, _04656_);
  nor (_04696_, _04517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04697_, _04696_, _04518_);
  and (_04698_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_04699_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  or (_04700_, _04699_, _04698_);
  and (_04701_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_04702_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  or (_04703_, _04702_, _04701_);
  or (_04704_, _04703_, _04700_);
  or (_04705_, _04704_, _04445_);
  and (_04706_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_04707_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  or (_04708_, _04707_, _04706_);
  and (_04709_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_04710_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  or (_04711_, _04710_, _04709_);
  or (_04712_, _04711_, _04708_);
  or (_04713_, _04712_, _04430_);
  and (_04714_, _04713_, _04485_);
  and (_04715_, _04714_, _04705_);
  and (_04716_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_04717_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  or (_04718_, _04717_, _04716_);
  and (_04719_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_04720_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  or (_04721_, _04720_, _04719_);
  or (_04722_, _04721_, _04718_);
  or (_04723_, _04722_, _04430_);
  and (_04724_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_04725_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  or (_04726_, _04725_, _04724_);
  and (_04727_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_04728_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  or (_04729_, _04728_, _04727_);
  or (_04730_, _04729_, _04726_);
  or (_04731_, _04730_, _04445_);
  and (_04732_, _04731_, _04426_);
  and (_04733_, _04732_, _04723_);
  or (_04734_, _04733_, _04715_);
  and (_04735_, _04734_, _04476_);
  and (_04736_, _04735_, _04697_);
  nor (_04737_, _04735_, _04697_);
  and (_04738_, _02500_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01920_);
  nor (_04740_, _04739_, _04738_);
  not (_04741_, _04740_);
  and (_04742_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_04743_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  or (_04744_, _04743_, _04742_);
  and (_04745_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_04746_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  or (_04747_, _04746_, _04745_);
  or (_04748_, _04747_, _04744_);
  or (_04749_, _04748_, _04430_);
  and (_04750_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_04751_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  or (_04752_, _04751_, _04750_);
  and (_04753_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_04754_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  or (_04755_, _04754_, _04753_);
  or (_04756_, _04755_, _04752_);
  or (_04757_, _04756_, _04445_);
  and (_04758_, _04757_, _04749_);
  or (_04759_, _04758_, _04485_);
  and (_04760_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_04761_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  or (_04762_, _04761_, _04760_);
  and (_04763_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_04764_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  or (_04765_, _04764_, _04763_);
  or (_04766_, _04765_, _04762_);
  or (_04767_, _04766_, _04430_);
  and (_04768_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_04769_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  or (_04770_, _04769_, _04768_);
  and (_04771_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_04772_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  or (_04773_, _04772_, _04771_);
  or (_04774_, _04773_, _04770_);
  or (_04775_, _04774_, _04445_);
  and (_04776_, _04775_, _04767_);
  or (_04777_, _04776_, _04426_);
  and (_04778_, _04777_, _04759_);
  and (_04779_, _04778_, _04476_);
  and (_04780_, _04779_, _04741_);
  and (_04781_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_04782_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  or (_04783_, _04782_, _04781_);
  and (_04784_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_04785_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  or (_04786_, _04785_, _04784_);
  or (_04787_, _04786_, _04783_);
  or (_04788_, _04787_, _04445_);
  and (_04789_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_04790_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or (_04791_, _04790_, _04789_);
  and (_04792_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_04793_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  or (_04794_, _04793_, _04792_);
  or (_04795_, _04794_, _04791_);
  or (_04796_, _04795_, _04430_);
  and (_04797_, _04796_, _04485_);
  and (_04798_, _04797_, _04788_);
  and (_04799_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_04800_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  or (_04801_, _04800_, _04799_);
  and (_04802_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_04803_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  or (_04804_, _04803_, _04802_);
  or (_04805_, _04804_, _04801_);
  or (_04806_, _04805_, _04430_);
  and (_04807_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_04808_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  or (_04809_, _04808_, _04807_);
  and (_04810_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_04811_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  or (_04812_, _04811_, _04810_);
  or (_04813_, _04812_, _04809_);
  or (_04814_, _04813_, _04445_);
  and (_04815_, _04814_, _04426_);
  and (_04816_, _04815_, _04806_);
  or (_04817_, _04816_, _04798_);
  and (_04818_, _04817_, _04476_);
  and (_04819_, _04818_, _02500_);
  and (_04820_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04821_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or (_04822_, _04821_, _04820_);
  and (_04823_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_04824_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  or (_04825_, _04824_, _04823_);
  or (_04826_, _04825_, _04822_);
  or (_04827_, _04826_, _04430_);
  and (_04828_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_04829_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or (_04830_, _04829_, _04828_);
  and (_04831_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04832_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  or (_04833_, _04832_, _04831_);
  or (_04834_, _04833_, _04830_);
  or (_04835_, _04834_, _04445_);
  and (_04836_, _04835_, _04827_);
  or (_04837_, _04836_, _04485_);
  and (_04838_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_04839_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  or (_04840_, _04839_, _04838_);
  and (_04841_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_04842_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or (_04843_, _04842_, _04841_);
  or (_04844_, _04843_, _04840_);
  or (_04845_, _04844_, _04445_);
  and (_04846_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_04847_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or (_04848_, _04847_, _04846_);
  and (_04849_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_04850_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  or (_04851_, _04850_, _04849_);
  or (_04852_, _04851_, _04848_);
  or (_04853_, _04852_, _04430_);
  and (_04854_, _04853_, _04845_);
  or (_04855_, _04854_, _04426_);
  and (_04856_, _04855_, _04837_);
  and (_04857_, _04856_, _04476_);
  and (_04858_, _04857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04859_, _04818_, _02500_);
  nor (_04860_, _04859_, _04819_);
  and (_04861_, _04860_, _04858_);
  nor (_04862_, _04861_, _04819_);
  nor (_04863_, _04779_, _04741_);
  nor (_04864_, _04863_, _04780_);
  not (_04865_, _04864_);
  nor (_04866_, _04865_, _04862_);
  nor (_04867_, _04866_, _04780_);
  nor (_04868_, _04867_, _04737_);
  nor (_04869_, _04868_, _04736_);
  nor (_04870_, _04694_, _04656_);
  nor (_04871_, _04870_, _04695_);
  not (_04872_, _04871_);
  nor (_04873_, _04872_, _04869_);
  nor (_04874_, _04873_, _04695_);
  nor (_04875_, _04874_, _04654_);
  nor (_04876_, _04875_, _04651_);
  nor (_04877_, _04876_, _04610_);
  nor (_04878_, _04877_, _04607_);
  nor (_04879_, _04878_, _04565_);
  or (_04880_, _04879_, _04564_);
  nor (_04881_, _04558_, _04516_);
  nor (_04882_, _04881_, _04559_);
  and (_04883_, _04882_, _04880_);
  and (_04884_, _04883_, _04561_);
  or (_04885_, _04884_, _04559_);
  nor (_04886_, _04885_, _04556_);
  nor (_04887_, _04886_, _04553_);
  and (_04888_, _04887_, _04550_);
  or (_04889_, _04888_, _04548_);
  nor (_04890_, _04889_, _04545_);
  nor (_04891_, _04534_, _04516_);
  nor (_04892_, _04891_, _04535_);
  not (_04893_, _04892_);
  nor (_04894_, _04893_, _04890_);
  and (_04895_, _04894_, _04541_);
  or (_04896_, _04895_, _04539_);
  nor (_04897_, _04896_, _04536_);
  nor (_04898_, _04531_, _04516_);
  nor (_04899_, _04898_, _04532_);
  not (_04900_, _04899_);
  nor (_04901_, _04900_, _04897_);
  nor (_04902_, _04901_, _04532_);
  nor (_04903_, _04529_, _04418_);
  and (_04904_, _04529_, _04418_);
  or (_04905_, _04904_, _04903_);
  and (_04906_, _04905_, _04516_);
  nor (_04907_, _04905_, _04516_);
  nor (_04908_, _04907_, _04906_);
  nor (_04909_, _04908_, _04902_);
  and (_04910_, _04908_, _04902_);
  or (_04911_, _04910_, _04909_);
  nor (_04912_, _04911_, _04421_);
  nor (_04913_, _04905_, cy_reg);
  nor (_04914_, _04913_, _04912_);
  nor (_04915_, _04914_, _02697_);
  and (_04916_, _04914_, _02697_);
  or (_04917_, _04916_, _04915_);
  nor (_04918_, _04894_, _04535_);
  and (_04919_, _04918_, _04541_);
  nor (_04920_, _04918_, _04541_);
  nor (_04921_, _04920_, _04919_);
  nor (_04922_, _04921_, _04421_);
  and (_04923_, _04538_, _04421_);
  nor (_04924_, _04923_, _04922_);
  nor (_04925_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_04926_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_04927_, _04547_, cy_reg);
  nor (_04928_, _04887_, _04544_);
  nor (_04929_, _04928_, _04550_);
  and (_04930_, _04928_, _04550_);
  or (_04931_, _04930_, _04929_);
  nor (_04932_, _04931_, _04421_);
  nor (_04933_, _04932_, _04927_);
  and (_04934_, _04933_, _01924_);
  nor (_04935_, _04933_, _01924_);
  and (_04936_, _04555_, _04421_);
  nor (_04937_, _04883_, _04559_);
  and (_04938_, _04937_, _04561_);
  nor (_04939_, _04937_, _04561_);
  nor (_04940_, _04939_, _04938_);
  nor (_04941_, _04940_, _04421_);
  nor (_04942_, _04941_, _04936_);
  nor (_04943_, _04942_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_04944_, _04942_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_04945_, _04563_, cy_reg);
  nor (_04946_, _04564_, _04565_);
  and (_04947_, _04946_, _04878_);
  nor (_04948_, _04946_, _04878_);
  or (_04949_, _04948_, _04947_);
  nor (_04950_, _04949_, _04421_);
  nor (_04951_, _04950_, _04945_);
  nor (_04952_, _04951_, _02415_);
  and (_04953_, _04951_, _02415_);
  and (_04954_, _04567_, _04421_);
  and (_04955_, _04876_, _04610_);
  nor (_04956_, _04955_, _04877_);
  and (_04957_, _04956_, cy_reg);
  nor (_04958_, _04957_, _04954_);
  and (_04959_, _04958_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_04960_, _04958_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_04961_, _04650_, _04421_);
  and (_04962_, _04874_, _04654_);
  nor (_04963_, _04962_, _04875_);
  and (_04964_, _04963_, cy_reg);
  nor (_04965_, _04964_, _04961_);
  and (_04966_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_04967_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_04968_, _04656_, _04421_);
  and (_04969_, _04872_, _04869_);
  nor (_04970_, _04969_, _04873_);
  and (_04971_, _04970_, cy_reg);
  nor (_04972_, _04971_, _04968_);
  and (_04973_, _04972_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_04974_, _04697_, cy_reg);
  nor (_04975_, _04737_, _04736_);
  nor (_04976_, _04975_, _04867_);
  and (_04977_, _04975_, _04867_);
  or (_04978_, _04977_, _04976_);
  nor (_04979_, _04978_, _04421_);
  nor (_04980_, _04979_, _04974_);
  nor (_04981_, _04980_, _02406_);
  and (_04982_, _04980_, _02406_);
  nor (_04983_, _04740_, cy_reg);
  and (_04984_, _04865_, _04862_);
  nor (_04985_, _04984_, _04866_);
  and (_04986_, _04985_, cy_reg);
  nor (_04987_, _04986_, _04983_);
  and (_04988_, _04987_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04989_, _04857_, cy_reg);
  not (_04990_, _04989_);
  nor (_04991_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04992_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04993_, _04992_, _04991_);
  nor (_04994_, _04993_, _04990_);
  and (_04995_, _04993_, _04990_);
  or (_04996_, _04995_, _04994_);
  nor (_04997_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_04998_, _04860_, _04858_);
  nor (_04999_, _04998_, _04861_);
  and (_05000_, _04999_, cy_reg);
  nor (_05001_, _05000_, _04997_);
  nor (_05002_, _05001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05003_, _05001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_05004_, _05003_, _05002_);
  or (_05005_, _05004_, _04996_);
  nor (_05006_, _04987_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05007_, _05006_, _05005_);
  or (_05008_, _05007_, _04988_);
  or (_05009_, _05008_, _04982_);
  or (_05010_, _05009_, _04981_);
  nor (_05011_, _04972_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_05012_, _05011_, _05010_);
  or (_05013_, _05012_, _04973_);
  or (_05014_, _05013_, _04967_);
  or (_05015_, _05014_, _04966_);
  or (_05016_, _05015_, _04960_);
  or (_05017_, _05016_, _04959_);
  or (_05018_, _05017_, _04953_);
  or (_05019_, _05018_, _04952_);
  and (_05020_, _04558_, _04421_);
  nor (_05021_, _04882_, _04880_);
  nor (_05022_, _05021_, _04883_);
  and (_05023_, _05022_, cy_reg);
  nor (_05024_, _05023_, _05020_);
  nor (_05025_, _05024_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_05026_, _05024_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_05027_, _05026_, _05025_);
  or (_05028_, _05027_, _05019_);
  or (_05029_, _05028_, _04944_);
  or (_05030_, _05029_, _04943_);
  and (_05031_, _04543_, _04421_);
  and (_05032_, _04886_, _04553_);
  nor (_05033_, _05032_, _04887_);
  and (_05034_, _05033_, cy_reg);
  nor (_05035_, _05034_, _05031_);
  and (_05036_, _05035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_05037_, _05035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_05038_, _05037_, _05036_);
  or (_05039_, _05038_, _05030_);
  or (_05040_, _05039_, _04935_);
  or (_05041_, _05040_, _04934_);
  and (_05042_, _04534_, _04421_);
  and (_05043_, _04893_, _04890_);
  nor (_05044_, _05043_, _04894_);
  and (_05045_, _05044_, cy_reg);
  nor (_05046_, _05045_, _05042_);
  and (_05047_, _05046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_05048_, _05046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_05049_, _05048_, _05047_);
  or (_05050_, _05049_, _05041_);
  or (_05051_, _05050_, _04926_);
  or (_05052_, _05051_, _04925_);
  and (_05053_, _04531_, _04421_);
  and (_05054_, _04900_, _04897_);
  nor (_05055_, _05054_, _04901_);
  and (_05056_, _05055_, cy_reg);
  nor (_05057_, _05056_, _05053_);
  and (_05058_, _05057_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_05059_, _05057_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_05060_, _05059_, _05058_);
  or (_05061_, _05060_, _05052_);
  or (_05062_, _05061_, _04917_);
  nor (_05063_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_05064_, _05063_, _02410_);
  nor (_05065_, _05064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05066_, _05064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05067_, _05066_, _05065_);
  or (_05068_, _01960_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05069_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05070_, _05069_, _05068_);
  or (_05071_, _05070_, _05067_);
  and (_05072_, _05063_, _02410_);
  nor (_05073_, _05072_, _05064_);
  not (_05074_, _05073_);
  or (_05075_, _01960_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_05077_, _05076_, _05075_);
  nand (_05078_, _05077_, _05067_);
  and (_05079_, _05078_, _05074_);
  and (_05080_, _05079_, _05071_);
  and (_05081_, _05067_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05082_, _02406_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_05083_, _05082_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_05084_, _05083_, _05081_);
  and (_05085_, _05067_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05086_, _02406_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05087_, _05086_, _01960_);
  or (_05088_, _05087_, _05085_);
  and (_05089_, _05088_, _05073_);
  and (_05090_, _05089_, _05084_);
  or (_05091_, _05090_, _05080_);
  and (_05092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05093_, _05092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_05094_, _05092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_05095_, _05094_, _05093_);
  not (_05096_, _05095_);
  nor (_05097_, _05093_, _02406_);
  and (_05098_, _05093_, _02406_);
  nor (_05099_, _05098_, _05097_);
  or (_05100_, _05099_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_05101_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_05102_, _05101_, _05100_);
  or (_05103_, _05102_, _05096_);
  nand (_05104_, _05099_, _08424_);
  or (_05105_, _05099_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05106_, _05105_, _05104_);
  or (_05107_, _05106_, _05095_);
  and (_05108_, _05107_, _05103_);
  or (_05109_, _05108_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_05110_, _05099_, _08796_);
  and (_05111_, _05099_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05112_, _05111_, _05110_);
  and (_05113_, _05112_, _05096_);
  or (_05114_, _05099_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05115_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05116_, _05115_, _05095_);
  and (_05117_, _05116_, _05114_);
  or (_05118_, _05117_, _01960_);
  or (_05119_, _05118_, _05113_);
  and (_05120_, _02406_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05121_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [15]);
  or (_05122_, _05121_, _05120_);
  and (_05123_, _05122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05124_, _02406_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05125_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05126_, _05125_, _02410_);
  and (_05127_, _05126_, _05124_);
  or (_05128_, _05127_, _05123_);
  and (_05129_, _05128_, _05092_);
  and (_05130_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _01960_);
  or (_05131_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05132_, _02406_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_05133_, _05132_, _05131_);
  or (_05134_, _05133_, _02410_);
  or (_05135_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05136_, _02406_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05137_, _05136_, _05135_);
  or (_05138_, _05137_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05139_, _05138_, _05134_);
  and (_05140_, _05139_, _05130_);
  or (_05141_, _05140_, _05129_);
  and (_05143_, _05128_, _01960_);
  or (_05144_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05145_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05146_, _02406_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05147_, _05146_, _05145_);
  and (_05148_, _05147_, _05144_);
  and (_05149_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _02410_);
  and (_05150_, _05149_, _05133_);
  or (_05151_, _05150_, _05148_);
  or (_05152_, _05151_, _05143_);
  and (_05153_, _05152_, _05141_);
  and (_05154_, _05153_, _05119_);
  and (_05155_, _05154_, _05109_);
  and (_05156_, _05155_, _05091_);
  and (_05157_, _05067_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or (_05158_, _05120_, _05074_);
  or (_05159_, _05158_, _05157_);
  and (_05160_, _05159_, _01960_);
  nor (_05161_, _05067_, _08262_);
  and (_05162_, _05067_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05163_, _05162_, _05161_);
  or (_05164_, _05163_, _05073_);
  and (_05165_, _05164_, _05160_);
  or (_05166_, _05165_, _05151_);
  and (_05167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05168_, _02406_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05169_, _05168_, _05167_);
  and (_05170_, _05169_, _02410_);
  and (_05171_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05172_, _05171_, _05082_);
  and (_05173_, _05172_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05174_, _05173_, _05170_);
  and (_05175_, _05174_, _01960_);
  or (_05176_, _05099_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_05177_, _05131_, _05095_);
  and (_05178_, _05177_, _05176_);
  or (_05179_, _05099_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand (_05180_, _05099_, _08276_);
  and (_05181_, _05180_, _05096_);
  and (_05182_, _05181_, _05179_);
  or (_05183_, _05182_, _05178_);
  and (_05184_, _05183_, _05175_);
  or (_05185_, _05099_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand (_05186_, _05099_, _08262_);
  and (_05187_, _05186_, _05096_);
  and (_05188_, _05187_, _05185_);
  or (_05189_, _05099_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or (_05190_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05191_, _05190_, _05095_);
  and (_05192_, _05191_, _05189_);
  or (_05193_, _05192_, _05188_);
  and (_05194_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_05195_, _05086_, _02410_);
  or (_05196_, _05195_, _05194_);
  or (_05197_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05198_, _02406_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05199_, _05198_, _05197_);
  or (_05200_, _05199_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05201_, _05200_, _05196_);
  and (_05202_, _05201_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05203_, _05172_, _05149_);
  or (_05204_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05205_, _02406_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05206_, _05205_, _05145_);
  and (_05207_, _05206_, _05204_);
  or (_05208_, _05207_, _05203_);
  and (_05209_, _05208_, _05202_);
  and (_05210_, _05209_, _05193_);
  or (_05211_, _05210_, _05184_);
  or (_05212_, _05208_, _05201_);
  and (_05213_, _05212_, _02402_);
  and (_05214_, _05213_, _05211_);
  and (_05215_, _05214_, _05166_);
  or (_05216_, _05215_, _05156_);
  nor (_05217_, _04453_, _01920_);
  nor (_05218_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_05219_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05220_, _05219_, _05218_);
  nand (_05221_, _05220_, _08298_);
  nor (_05222_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05223_, _05222_, _02505_);
  nor (_05224_, _05223_, _05217_);
  and (_05225_, _05224_, _04442_);
  and (_05226_, _05225_, _05221_);
  not (_05227_, _05224_);
  and (_05228_, _05220_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05229_, _05220_, _08424_);
  or (_05230_, _05229_, _05228_);
  and (_05231_, _05230_, _05227_);
  or (_05232_, _05231_, _05226_);
  and (_05233_, _05232_, _04422_);
  nand (_05234_, _05220_, _08967_);
  or (_05235_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05236_, _05235_, _05224_);
  and (_05237_, _05236_, _05234_);
  and (_05238_, _05220_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05239_, _05220_, _08276_);
  or (_05240_, _05239_, _05238_);
  and (_05241_, _05240_, _05227_);
  or (_05242_, _05241_, _05237_);
  and (_05243_, _05242_, _04464_);
  or (_05244_, _05243_, _05233_);
  nand (_05245_, _05220_, _08270_);
  or (_05246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05247_, _05246_, _05224_);
  and (_05248_, _05247_, _05245_);
  and (_05249_, _05220_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05250_, _05220_, _08262_);
  or (_05251_, _05250_, _05249_);
  and (_05252_, _05251_, _05227_);
  or (_05253_, _05252_, _05248_);
  and (_05254_, _05253_, _04453_);
  nand (_05255_, _05220_, _08302_);
  and (_05256_, _05224_, _04431_);
  and (_05257_, _05256_, _05255_);
  and (_05258_, _05220_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05259_, _05220_, _08293_);
  or (_05260_, _05259_, _05258_);
  and (_05261_, _05260_, _05227_);
  or (_05262_, _05261_, _05257_);
  and (_05263_, _05262_, _04440_);
  or (_05264_, _05263_, _05254_);
  or (_05265_, _05264_, _05244_);
  not (_05266_, _04422_);
  nor (_05267_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_05268_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_05269_, _05268_, _05267_);
  or (_05270_, _05269_, _05266_);
  nor (_05271_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_05272_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand (_05273_, _05272_, _05271_);
  nand (_05274_, _05273_, _04440_);
  and (_05275_, _05274_, _05270_);
  nor (_05276_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_05277_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand (_05278_, _05277_, _05276_);
  nand (_05279_, _05278_, _04464_);
  not (_05280_, _04453_);
  nor (_05281_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_05282_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_05283_, _05282_, _05281_);
  or (_05284_, _05283_, _05280_);
  and (_05285_, _05284_, _05279_);
  and (_05286_, _05285_, _05275_);
  and (_05287_, _04422_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_05288_, _04464_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or (_05289_, _05288_, _05287_);
  and (_05290_, _04453_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_05291_, _04440_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or (_05292_, _05291_, _05290_);
  or (_05293_, _05292_, _05289_);
  nand (_05294_, _04464_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_05295_, _04440_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_05296_, _05295_, _05294_);
  nand (_05297_, _04422_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_05298_, _04453_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05299_, _05298_, _05297_);
  and (_05300_, _05299_, _05296_);
  or (_05301_, \oc8051_symbolic_cxrom1.regarray[9] [5], \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nand (_05302_, _05301_, _04440_);
  or (_05303_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nand (_05304_, _05303_, _04464_);
  and (_05305_, _05304_, _05302_);
  or (_05306_, \oc8051_symbolic_cxrom1.regarray[11] [5], \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nand (_05307_, _05306_, _04422_);
  or (_05308_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nand (_05309_, _05308_, _04453_);
  and (_05310_, _05309_, _05307_);
  and (_05311_, _05310_, _05305_);
  and (_05312_, _05311_, _05300_);
  and (_05313_, _05312_, _05293_);
  and (_05314_, _05313_, _05286_);
  or (_05315_, _05314_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_05316_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_05317_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_05318_, _05317_, _05316_);
  or (_05319_, _05318_, _05280_);
  nor (_05320_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_05321_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_05322_, _05321_, _05320_);
  or (_05323_, _05322_, _05266_);
  and (_05324_, _05323_, _05319_);
  nor (_05325_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_05326_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_05327_, _05326_, _05325_);
  nand (_05328_, _05327_, _04464_);
  nor (_05329_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_05330_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand (_05331_, _05330_, _05329_);
  nand (_05332_, _05331_, _04440_);
  and (_05333_, _05332_, _05328_);
  and (_05334_, _05333_, _05324_);
  and (_05335_, _04422_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_05336_, _04464_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or (_05337_, _05336_, _05335_);
  and (_05338_, _04440_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_05339_, _04453_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or (_05340_, _05339_, _05338_);
  or (_05341_, _05340_, _05337_);
  nand (_05342_, _04464_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  or (_05343_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nand (_05344_, _05343_, _04464_);
  and (_05345_, _05344_, _05342_);
  nand (_05346_, _04422_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_05347_, _04453_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_05348_, _05347_, _05346_);
  and (_05349_, _05348_, _05345_);
  nand (_05350_, _04440_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  or (_05351_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand (_05352_, _05351_, _04453_);
  and (_05353_, _05352_, _05350_);
  or (_05354_, \oc8051_symbolic_cxrom1.regarray[15] [5], \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand (_05355_, _05354_, _04422_);
  or (_05356_, \oc8051_symbolic_cxrom1.regarray[13] [5], \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nand (_05357_, _05356_, _04440_);
  and (_05358_, _05357_, _05355_);
  and (_05359_, _05358_, _05353_);
  and (_05360_, _05359_, _05349_);
  and (_05361_, _05360_, _05341_);
  and (_05362_, _05361_, _05334_);
  or (_05363_, _05362_, _01920_);
  and (_05364_, _05363_, _05315_);
  or (_05365_, _05364_, _02512_);
  or (_05366_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand (_05367_, _05366_, _04464_);
  and (_05368_, _05367_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_05369_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand (_05370_, _05369_, _04422_);
  or (_05371_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_05372_, _05371_, _04440_);
  and (_05373_, _05372_, _05370_);
  or (_05374_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand (_05375_, _05374_, _04453_);
  or (_05376_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nand (_05377_, _05376_, _04453_);
  and (_05378_, _05377_, _05375_);
  and (_05379_, _05378_, _05373_);
  and (_05380_, _05379_, _05368_);
  nand (_05381_, _04440_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or (_05382_, \oc8051_symbolic_cxrom1.regarray[5] [5], \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nand (_05383_, _05382_, _04440_);
  and (_05384_, _05383_, _05381_);
  or (_05385_, \oc8051_symbolic_cxrom1.regarray[7] [5], \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand (_05386_, _05385_, _04422_);
  or (_05387_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nand (_05388_, _05387_, _04464_);
  and (_05389_, _05388_, _05386_);
  and (_05390_, _05389_, _05384_);
  nand (_05391_, _04464_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  or (_05392_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand (_05393_, _05392_, _04453_);
  and (_05394_, _05393_, _05391_);
  nand (_05395_, _04422_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_05396_, _04453_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_05397_, _05396_, _05395_);
  and (_05398_, _05397_, _05394_);
  and (_05399_, _05398_, _05390_);
  and (_05400_, _04440_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_05401_, _04453_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or (_05402_, _05401_, _05400_);
  and (_05403_, _04422_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_05404_, _04464_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or (_05405_, _05404_, _05403_);
  or (_05406_, _05405_, _05402_);
  or (_05407_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand (_05408_, _05407_, _04464_);
  or (_05409_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand (_05410_, _05409_, _04422_);
  or (_05411_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand (_05412_, _05411_, _04440_);
  and (_05413_, _05412_, _05410_);
  and (_05414_, _05413_, _05408_);
  and (_05415_, _05414_, _05406_);
  and (_05416_, _05415_, _05399_);
  and (_05417_, _05416_, _05380_);
  nand (_05418_, _04440_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_05419_, _05418_, _01920_);
  or (_05420_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nand (_05421_, _05420_, _04453_);
  or (_05422_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand (_05423_, _05422_, _04453_);
  and (_05424_, _05423_, _05421_);
  or (_05425_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand (_05426_, _05425_, _04464_);
  or (_05427_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_05428_, _05427_, _04440_);
  and (_05429_, _05428_, _05426_);
  and (_05430_, _05429_, _05424_);
  and (_05431_, _05430_, _05419_);
  nand (_05432_, _04453_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  or (_05433_, \oc8051_symbolic_cxrom1.regarray[1] [5], \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand (_05434_, _05433_, _04440_);
  and (_05435_, _05434_, _05432_);
  or (_05436_, \oc8051_symbolic_cxrom1.regarray[3] [5], \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand (_05437_, _05436_, _04422_);
  or (_05438_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nand (_05439_, _05438_, _04464_);
  and (_05440_, _05439_, _05437_);
  and (_05441_, _05440_, _05435_);
  nand (_05442_, _04464_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_05443_, _04422_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_05444_, _05443_, _05442_);
  or (_05445_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand (_05446_, _05445_, _04422_);
  or (_05447_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand (_05448_, _05447_, _04453_);
  and (_05449_, _05448_, _05446_);
  and (_05450_, _05449_, _05444_);
  and (_05451_, _05450_, _05441_);
  and (_05452_, _04453_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_05453_, _04440_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or (_05454_, _05453_, _05452_);
  and (_05455_, _04464_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_05456_, _04422_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  or (_05457_, _05456_, _05455_);
  or (_05458_, _05457_, _05454_);
  or (_05459_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand (_05460_, _05459_, _04464_);
  or (_05461_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand (_05462_, _05461_, _04422_);
  or (_05463_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand (_05464_, _05463_, _04440_);
  and (_05465_, _05464_, _05462_);
  and (_05466_, _05465_, _05460_);
  and (_05467_, _05466_, _05458_);
  and (_05468_, _05467_, _05451_);
  and (_05469_, _05468_, _05431_);
  or (_05470_, _05469_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05471_, _05470_, _05417_);
  and (_05472_, _05246_, _04466_);
  or (_05473_, _05472_, _01920_);
  or (_05474_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05475_, _02512_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05476_, _05475_, _05474_);
  or (_05477_, _05476_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05478_, _05477_, _05473_);
  and (_05479_, _05478_, _04440_);
  and (_05480_, _04464_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_05481_, _02512_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05482_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05483_, _05482_, _05481_);
  and (_05484_, _05483_, _05480_);
  or (_05485_, _02512_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05486_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05487_, _05486_, _05485_);
  and (_05488_, _05487_, _04423_);
  or (_05489_, _05488_, _05484_);
  or (_05490_, _05489_, _05479_);
  or (_05491_, _02512_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05492_, _05491_, _04431_);
  or (_05493_, _05492_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05494_, _05235_, _04455_);
  or (_05495_, _05494_, _02505_);
  and (_05496_, _05495_, _04739_);
  and (_05497_, _05496_, _05493_);
  or (_05498_, _02512_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05499_, _04442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05500_, _05499_, _05498_);
  or (_05501_, _02512_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05502_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_05503_, _05502_, _01920_);
  and (_05504_, _05503_, _05501_);
  or (_05505_, _05504_, _05500_);
  and (_05506_, _05505_, _04453_);
  or (_05507_, _05506_, _05497_);
  or (_05508_, _05507_, _05490_);
  and (_05509_, _05505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05510_, _05492_, _04738_);
  or (_05511_, _02512_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05513_, _05512_, _05222_);
  and (_05514_, _05513_, _05511_);
  or (_05515_, _05514_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_05516_, _05515_, _05510_);
  or (_05517_, _05516_, _05509_);
  and (_05518_, _05478_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05519_, _05494_, _04738_);
  and (_05520_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05521_, _02512_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05522_, _05521_, _05520_);
  and (_05523_, _05522_, _05222_);
  or (_05524_, _05523_, _02505_);
  or (_05525_, _05524_, _05519_);
  or (_05526_, _05525_, _05518_);
  nor (_05527_, _01956_, first_instr);
  and (_05528_, _05527_, _05526_);
  and (_05529_, _05528_, _05517_);
  and (_05530_, _05529_, _05508_);
  and (_05531_, _05530_, _05471_);
  and (_05532_, _05531_, _05365_);
  and (_05533_, _05532_, _04476_);
  and (_05534_, _05533_, _05265_);
  and (_05535_, _05534_, _05216_);
  and (property_invalid_jc, _05535_, _05062_);
  or (_05536_, pc_log_change_r, _04421_);
  nand (_05537_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_00000_, _05537_, _05536_);
  and (_05538_, _01956_, first_instr);
  or (_00001_, _05538_, rst);
  dff (cy_reg, _00000_);
  dff (pc_log_change_r, pc_log_change);
  dff (first_instr, _00001_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _13870_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _13871_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _13872_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _13873_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _13874_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _13875_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _13876_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _13877_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _09923_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _09925_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _09926_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _09929_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _09932_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _09935_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _09939_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _09941_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _13869_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _09832_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _09836_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _09840_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _09842_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _09845_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _09847_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _09850_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _09751_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _09755_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _09758_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _09760_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _09762_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _09765_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _09769_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _09772_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _13861_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _13862_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _13863_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _13864_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _13865_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _13866_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _13867_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _13868_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _13853_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _13854_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _13855_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _13856_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _13857_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _13858_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _13859_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _13860_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _13898_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _13899_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _13900_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _13901_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _13902_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _13903_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _13904_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _13905_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _09403_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _09408_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _13892_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _13893_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _13894_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _13895_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _13896_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _13897_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _13884_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _13885_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _13886_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _13887_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _13888_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _13889_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _13890_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _13891_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _09217_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _09220_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _09224_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _09229_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _09233_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _09235_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _09238_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _09242_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _09110_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _09115_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _09120_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _09125_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _09129_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _09134_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _09138_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _09141_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _08705_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _08709_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _08712_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _08715_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _08717_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _08719_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _08721_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _08724_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _08586_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _08591_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _08597_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _08600_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _08606_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _08612_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _08617_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _08619_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _13879_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _08899_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _08902_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _08907_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _08912_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _08916_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _08919_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _08922_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _08801_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _08805_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _08810_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _08814_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _08817_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _13878_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _08822_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _08825_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _09011_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _09016_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _13880_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _13881_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _13882_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _13883_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _09034_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _09037_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _07256_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _07287_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _07324_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _07361_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _07415_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _07480_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _07541_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _07615_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _07673_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _07739_);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _07829_);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _07927_);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _08032_);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _08119_);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _08231_);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _07207_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _04128_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _04074_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _04054_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _04050_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _12807_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _03846_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03614_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _10695_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _13506_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _13470_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _00331_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _00235_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _00205_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _00153_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _00085_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _03883_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11685_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _10840_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _06005_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _06036_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _06017_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _06013_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _06007_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11741_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _12386_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _06548_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _00475_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _00910_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _01737_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _03645_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04571_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _03742_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _06907_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _06909_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _06912_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _06914_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _06917_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _06920_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _06923_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06780_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _12033_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _01125_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12598_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _04080_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _01436_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _07502_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _04142_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _02378_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _04144_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _07409_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _07268_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _03600_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _03347_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _07341_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _02850_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _02838_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _04168_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _04091_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03548_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04062_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03824_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _04176_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _04490_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _10247_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _04179_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _10693_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _10282_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04181_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03671_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _04184_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _11293_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _11295_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03558_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _04186_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _11720_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _04188_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _04221_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _00251_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _00328_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _02609_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _02612_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _01932_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _02330_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _02545_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _02503_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _03324_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _04166_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _02536_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _03720_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _05581_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _01631_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _11191_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _02190_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _03332_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _02413_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _06961_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _03673_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _11681_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _10816_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _05578_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12281_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _03446_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03914_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _13761_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _00219_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _02471_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _00060_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _10361_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _02165_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _00076_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _11882_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _06623_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _02353_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _03769_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _13682_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _04052_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03636_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _03850_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _06610_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _11755_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _12772_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _11298_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _11748_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _11302_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _13157_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _03888_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _00025_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _11229_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _02818_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _11880_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _02286_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _11869_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01895_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _00247_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _08551_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _08614_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _03270_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _02012_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _02010_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _08845_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _03566_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _00122_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _02597_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _11963_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _11184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _13222_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _11375_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _01437_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _00999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _01447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _01444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _00996_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01077_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _01453_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _01449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _00992_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _01493_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _01459_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _00962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _01135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _01150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _02604_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _01569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _00941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01584_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01571_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _00938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _01065_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _01593_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _01587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _00933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _01596_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _01594_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _00925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _01062_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _01130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _04429_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _03454_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04082_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _04044_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _03936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _03902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _03873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _11974_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _11165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _11355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _11551_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _00549_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _04015_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _04352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _04284_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _04275_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _04017_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _11984_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _00395_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _07338_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03784_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _01666_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _05764_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _11981_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _11162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _12011_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _01193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _08287_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _11992_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _02450_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _00159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _11259_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _03750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _12003_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _11156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03441_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _03439_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _03436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _03433_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _05672_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _06468_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _01918_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _00894_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _12370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _12361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _12346_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _12343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _12286_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _12275_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _12065_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _12440_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _12523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _12520_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _12058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _11110_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _11826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _11798_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _10889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _11168_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _11146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _11013_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _12087_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _11588_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _11369_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _11554_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _11438_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11417_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _12078_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _11096_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _10302_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _10263_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _10298_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _08560_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _11498_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _01864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _11504_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _00606_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _07307_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _01713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _02537_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12105_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _07083_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _06264_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _01884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _06607_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _12102_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _01887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _11143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _11350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _11047_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _11319_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _11517_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _02376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _02382_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _01899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _02089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _12110_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _11044_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _03705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _03467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _06484_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11034_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11314_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _03660_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _03771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _03712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _03679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _12135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _06592_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _06691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _08435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _02706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _02519_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _02238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _10089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _10928_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _10269_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _10033_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11104_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _10640_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _12070_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _10637_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _00071_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _12079_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _10634_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _10813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _10916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _10985_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _00206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _00201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _10631_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _00771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _00291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _10628_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _10810_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _01797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _01352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _10625_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _02571_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _01817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _10623_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _10807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _10903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _02708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _03415_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _02253_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _01664_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _01761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _03814_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _03775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _10604_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _10731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _02255_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _04133_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _12084_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _12115_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _12113_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04039_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _04154_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _04147_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _11841_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _11897_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _11894_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _11888_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _11885_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03665_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03526_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _11659_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _07973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _02456_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _11049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _02458_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _01630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _07968_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _05610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _03603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _00815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _00807_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _03593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _00533_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _00530_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _03638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03895_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _07109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _02168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _05866_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _03398_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _05929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07080_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _05899_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _02153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _04295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _05932_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12026_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _10951_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _02677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _13282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _13271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _13279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _13276_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _02867_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _13296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _02498_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _02636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _04077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _03681_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _13262_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _13250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _03329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _02668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _13150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _12455_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _13142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _13175_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _00274_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _00269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08444_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _10257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _13109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _13106_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _02889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _10254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _13569_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _13564_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _13558_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _02805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _13590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _13587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _13580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _00336_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _13543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _02815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _02654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _13493_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _13490_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _13483_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _02821_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _04414_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _03138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _03305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _03136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _03172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _03623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _03283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _03132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _03162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _05142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _03311_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _03160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _02004_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _03126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _03317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03287_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _03286_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _03158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _06900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _06894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _06964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _07223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _07139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _04069_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _00271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _13680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _03675_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _13726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _13709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _13720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _13717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _13714_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _03651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01080_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _01083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _13154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _13163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _13167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _13135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _13132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _13129_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _13139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _01094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _13197_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _13191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _13194_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _13212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _13203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _13209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _13206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _01088_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _01092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _01090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _13219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _13215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13301_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _01042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13370_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13364_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13340_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13351_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _01046_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _01044_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13376_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13378_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13396_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13393_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _01057_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _03495_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _02435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _02074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _01549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _01547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _01545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _01542_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _01539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _01490_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _01480_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _09910_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _01421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _01403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _01363_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _01395_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _01391_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _01387_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _01366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01794_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _03966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _01265_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _01216_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _01201_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _01211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _01207_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _01182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _01169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _03493_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _01143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _01103_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _01097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _01086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _01037_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _01034_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _01028_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _03078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _00793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _00990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _00970_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _00966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _00930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _00928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _00922_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _00917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _00514_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _05541_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _05540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _05539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _02328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01099_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _02117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01904_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _11021_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _03276_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _00342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _00604_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _02834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _11823_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _01686_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _10954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _02779_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _03346_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _01680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _03881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _07822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _11357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _06338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _07180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _07858_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _02540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _06460_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _10900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _02468_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _02465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _02474_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _11758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _09164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _02831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _02739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _02836_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _02736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _00684_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _00682_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _12067_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _12055_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _03048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _03014_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _12049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _12191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _12326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _12358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _03153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _03075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _02853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _03714_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _03522_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _12042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _12158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _12323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _03844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _03718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _02851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _03974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _12023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _12151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _12294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _12356_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _12383_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _04020_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02726_);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
